
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_regfile ( suppress_key_tlvs, kme_interrupt, .rbus_ring_o( {
	\rbus_ring_o.addr [15], \rbus_ring_o.addr [14], 
	\rbus_ring_o.addr [13], \rbus_ring_o.addr [12], 
	\rbus_ring_o.addr [11], \rbus_ring_o.addr [10], 
	\rbus_ring_o.addr [9], \rbus_ring_o.addr [8], \rbus_ring_o.addr [7], 
	\rbus_ring_o.addr [6], \rbus_ring_o.addr [5], \rbus_ring_o.addr [4], 
	\rbus_ring_o.addr [3], \rbus_ring_o.addr [2], \rbus_ring_o.addr [1], 
	\rbus_ring_o.addr [0], \rbus_ring_o.wr_strb , 
	\rbus_ring_o.wr_data [31], \rbus_ring_o.wr_data [30], 
	\rbus_ring_o.wr_data [29], \rbus_ring_o.wr_data [28], 
	\rbus_ring_o.wr_data [27], \rbus_ring_o.wr_data [26], 
	\rbus_ring_o.wr_data [25], \rbus_ring_o.wr_data [24], 
	\rbus_ring_o.wr_data [23], \rbus_ring_o.wr_data [22], 
	\rbus_ring_o.wr_data [21], \rbus_ring_o.wr_data [20], 
	\rbus_ring_o.wr_data [19], \rbus_ring_o.wr_data [18], 
	\rbus_ring_o.wr_data [17], \rbus_ring_o.wr_data [16], 
	\rbus_ring_o.wr_data [15], \rbus_ring_o.wr_data [14], 
	\rbus_ring_o.wr_data [13], \rbus_ring_o.wr_data [12], 
	\rbus_ring_o.wr_data [11], \rbus_ring_o.wr_data [10], 
	\rbus_ring_o.wr_data [9], \rbus_ring_o.wr_data [8], 
	\rbus_ring_o.wr_data [7], \rbus_ring_o.wr_data [6], 
	\rbus_ring_o.wr_data [5], \rbus_ring_o.wr_data [4], 
	\rbus_ring_o.wr_data [3], \rbus_ring_o.wr_data [2], 
	\rbus_ring_o.wr_data [1], \rbus_ring_o.wr_data [0], 
	\rbus_ring_o.rd_strb , \rbus_ring_o.rd_data [31], 
	\rbus_ring_o.rd_data [30], \rbus_ring_o.rd_data [29], 
	\rbus_ring_o.rd_data [28], \rbus_ring_o.rd_data [27], 
	\rbus_ring_o.rd_data [26], \rbus_ring_o.rd_data [25], 
	\rbus_ring_o.rd_data [24], \rbus_ring_o.rd_data [23], 
	\rbus_ring_o.rd_data [22], \rbus_ring_o.rd_data [21], 
	\rbus_ring_o.rd_data [20], \rbus_ring_o.rd_data [19], 
	\rbus_ring_o.rd_data [18], \rbus_ring_o.rd_data [17], 
	\rbus_ring_o.rd_data [16], \rbus_ring_o.rd_data [15], 
	\rbus_ring_o.rd_data [14], \rbus_ring_o.rd_data [13], 
	\rbus_ring_o.rd_data [12], \rbus_ring_o.rd_data [11], 
	\rbus_ring_o.rd_data [10], \rbus_ring_o.rd_data [9], 
	\rbus_ring_o.rd_data [8], \rbus_ring_o.rd_data [7], 
	\rbus_ring_o.rd_data [6], \rbus_ring_o.rd_data [5], 
	\rbus_ring_o.rd_data [4], \rbus_ring_o.rd_data [3], 
	\rbus_ring_o.rd_data [2], \rbus_ring_o.rd_data [1], 
	\rbus_ring_o.rd_data [0], \rbus_ring_o.ack , \rbus_ring_o.err_ack } ), 
	.kme_cceip0_ob_out( {\kme_cceip0_ob_out.tvalid , 
	\kme_cceip0_ob_out.tlast , \kme_cceip0_ob_out.tid [0], 
	\kme_cceip0_ob_out.tstrb [7], \kme_cceip0_ob_out.tstrb [6], 
	\kme_cceip0_ob_out.tstrb [5], \kme_cceip0_ob_out.tstrb [4], 
	\kme_cceip0_ob_out.tstrb [3], \kme_cceip0_ob_out.tstrb [2], 
	\kme_cceip0_ob_out.tstrb [1], \kme_cceip0_ob_out.tstrb [0], 
	\kme_cceip0_ob_out.tuser [7], \kme_cceip0_ob_out.tuser [6], 
	\kme_cceip0_ob_out.tuser [5], \kme_cceip0_ob_out.tuser [4], 
	\kme_cceip0_ob_out.tuser [3], \kme_cceip0_ob_out.tuser [2], 
	\kme_cceip0_ob_out.tuser [1], \kme_cceip0_ob_out.tuser [0], 
	\kme_cceip0_ob_out.tdata [63], \kme_cceip0_ob_out.tdata [62], 
	\kme_cceip0_ob_out.tdata [61], \kme_cceip0_ob_out.tdata [60], 
	\kme_cceip0_ob_out.tdata [59], \kme_cceip0_ob_out.tdata [58], 
	\kme_cceip0_ob_out.tdata [57], \kme_cceip0_ob_out.tdata [56], 
	\kme_cceip0_ob_out.tdata [55], \kme_cceip0_ob_out.tdata [54], 
	\kme_cceip0_ob_out.tdata [53], \kme_cceip0_ob_out.tdata [52], 
	\kme_cceip0_ob_out.tdata [51], \kme_cceip0_ob_out.tdata [50], 
	\kme_cceip0_ob_out.tdata [49], \kme_cceip0_ob_out.tdata [48], 
	\kme_cceip0_ob_out.tdata [47], \kme_cceip0_ob_out.tdata [46], 
	\kme_cceip0_ob_out.tdata [45], \kme_cceip0_ob_out.tdata [44], 
	\kme_cceip0_ob_out.tdata [43], \kme_cceip0_ob_out.tdata [42], 
	\kme_cceip0_ob_out.tdata [41], \kme_cceip0_ob_out.tdata [40], 
	\kme_cceip0_ob_out.tdata [39], \kme_cceip0_ob_out.tdata [38], 
	\kme_cceip0_ob_out.tdata [37], \kme_cceip0_ob_out.tdata [36], 
	\kme_cceip0_ob_out.tdata [35], \kme_cceip0_ob_out.tdata [34], 
	\kme_cceip0_ob_out.tdata [33], \kme_cceip0_ob_out.tdata [32], 
	\kme_cceip0_ob_out.tdata [31], \kme_cceip0_ob_out.tdata [30], 
	\kme_cceip0_ob_out.tdata [29], \kme_cceip0_ob_out.tdata [28], 
	\kme_cceip0_ob_out.tdata [27], \kme_cceip0_ob_out.tdata [26], 
	\kme_cceip0_ob_out.tdata [25], \kme_cceip0_ob_out.tdata [24], 
	\kme_cceip0_ob_out.tdata [23], \kme_cceip0_ob_out.tdata [22], 
	\kme_cceip0_ob_out.tdata [21], \kme_cceip0_ob_out.tdata [20], 
	\kme_cceip0_ob_out.tdata [19], \kme_cceip0_ob_out.tdata [18], 
	\kme_cceip0_ob_out.tdata [17], \kme_cceip0_ob_out.tdata [16], 
	\kme_cceip0_ob_out.tdata [15], \kme_cceip0_ob_out.tdata [14], 
	\kme_cceip0_ob_out.tdata [13], \kme_cceip0_ob_out.tdata [12], 
	\kme_cceip0_ob_out.tdata [11], \kme_cceip0_ob_out.tdata [10], 
	\kme_cceip0_ob_out.tdata [9], \kme_cceip0_ob_out.tdata [8], 
	\kme_cceip0_ob_out.tdata [7], \kme_cceip0_ob_out.tdata [6], 
	\kme_cceip0_ob_out.tdata [5], \kme_cceip0_ob_out.tdata [4], 
	\kme_cceip0_ob_out.tdata [3], \kme_cceip0_ob_out.tdata [2], 
	\kme_cceip0_ob_out.tdata [1], \kme_cceip0_ob_out.tdata [0]} ), 
	.kme_cceip0_ob_in_mod( {\kme_cceip0_ob_in_mod.tready } ), 
	.kme_cceip1_ob_out( {\kme_cceip1_ob_out.tvalid , 
	\kme_cceip1_ob_out.tlast , \kme_cceip1_ob_out.tid [0], 
	\kme_cceip1_ob_out.tstrb [7], \kme_cceip1_ob_out.tstrb [6], 
	\kme_cceip1_ob_out.tstrb [5], \kme_cceip1_ob_out.tstrb [4], 
	\kme_cceip1_ob_out.tstrb [3], \kme_cceip1_ob_out.tstrb [2], 
	\kme_cceip1_ob_out.tstrb [1], \kme_cceip1_ob_out.tstrb [0], 
	\kme_cceip1_ob_out.tuser [7], \kme_cceip1_ob_out.tuser [6], 
	\kme_cceip1_ob_out.tuser [5], \kme_cceip1_ob_out.tuser [4], 
	\kme_cceip1_ob_out.tuser [3], \kme_cceip1_ob_out.tuser [2], 
	\kme_cceip1_ob_out.tuser [1], \kme_cceip1_ob_out.tuser [0], 
	\kme_cceip1_ob_out.tdata [63], \kme_cceip1_ob_out.tdata [62], 
	\kme_cceip1_ob_out.tdata [61], \kme_cceip1_ob_out.tdata [60], 
	\kme_cceip1_ob_out.tdata [59], \kme_cceip1_ob_out.tdata [58], 
	\kme_cceip1_ob_out.tdata [57], \kme_cceip1_ob_out.tdata [56], 
	\kme_cceip1_ob_out.tdata [55], \kme_cceip1_ob_out.tdata [54], 
	\kme_cceip1_ob_out.tdata [53], \kme_cceip1_ob_out.tdata [52], 
	\kme_cceip1_ob_out.tdata [51], \kme_cceip1_ob_out.tdata [50], 
	\kme_cceip1_ob_out.tdata [49], \kme_cceip1_ob_out.tdata [48], 
	\kme_cceip1_ob_out.tdata [47], \kme_cceip1_ob_out.tdata [46], 
	\kme_cceip1_ob_out.tdata [45], \kme_cceip1_ob_out.tdata [44], 
	\kme_cceip1_ob_out.tdata [43], \kme_cceip1_ob_out.tdata [42], 
	\kme_cceip1_ob_out.tdata [41], \kme_cceip1_ob_out.tdata [40], 
	\kme_cceip1_ob_out.tdata [39], \kme_cceip1_ob_out.tdata [38], 
	\kme_cceip1_ob_out.tdata [37], \kme_cceip1_ob_out.tdata [36], 
	\kme_cceip1_ob_out.tdata [35], \kme_cceip1_ob_out.tdata [34], 
	\kme_cceip1_ob_out.tdata [33], \kme_cceip1_ob_out.tdata [32], 
	\kme_cceip1_ob_out.tdata [31], \kme_cceip1_ob_out.tdata [30], 
	\kme_cceip1_ob_out.tdata [29], \kme_cceip1_ob_out.tdata [28], 
	\kme_cceip1_ob_out.tdata [27], \kme_cceip1_ob_out.tdata [26], 
	\kme_cceip1_ob_out.tdata [25], \kme_cceip1_ob_out.tdata [24], 
	\kme_cceip1_ob_out.tdata [23], \kme_cceip1_ob_out.tdata [22], 
	\kme_cceip1_ob_out.tdata [21], \kme_cceip1_ob_out.tdata [20], 
	\kme_cceip1_ob_out.tdata [19], \kme_cceip1_ob_out.tdata [18], 
	\kme_cceip1_ob_out.tdata [17], \kme_cceip1_ob_out.tdata [16], 
	\kme_cceip1_ob_out.tdata [15], \kme_cceip1_ob_out.tdata [14], 
	\kme_cceip1_ob_out.tdata [13], \kme_cceip1_ob_out.tdata [12], 
	\kme_cceip1_ob_out.tdata [11], \kme_cceip1_ob_out.tdata [10], 
	\kme_cceip1_ob_out.tdata [9], \kme_cceip1_ob_out.tdata [8], 
	\kme_cceip1_ob_out.tdata [7], \kme_cceip1_ob_out.tdata [6], 
	\kme_cceip1_ob_out.tdata [5], \kme_cceip1_ob_out.tdata [4], 
	\kme_cceip1_ob_out.tdata [3], \kme_cceip1_ob_out.tdata [2], 
	\kme_cceip1_ob_out.tdata [1], \kme_cceip1_ob_out.tdata [0]} ), 
	.kme_cceip1_ob_in_mod( {\kme_cceip1_ob_in_mod.tready } ), 
	.kme_cceip2_ob_out( {\kme_cceip2_ob_out.tvalid , 
	\kme_cceip2_ob_out.tlast , \kme_cceip2_ob_out.tid [0], 
	\kme_cceip2_ob_out.tstrb [7], \kme_cceip2_ob_out.tstrb [6], 
	\kme_cceip2_ob_out.tstrb [5], \kme_cceip2_ob_out.tstrb [4], 
	\kme_cceip2_ob_out.tstrb [3], \kme_cceip2_ob_out.tstrb [2], 
	\kme_cceip2_ob_out.tstrb [1], \kme_cceip2_ob_out.tstrb [0], 
	\kme_cceip2_ob_out.tuser [7], \kme_cceip2_ob_out.tuser [6], 
	\kme_cceip2_ob_out.tuser [5], \kme_cceip2_ob_out.tuser [4], 
	\kme_cceip2_ob_out.tuser [3], \kme_cceip2_ob_out.tuser [2], 
	\kme_cceip2_ob_out.tuser [1], \kme_cceip2_ob_out.tuser [0], 
	\kme_cceip2_ob_out.tdata [63], \kme_cceip2_ob_out.tdata [62], 
	\kme_cceip2_ob_out.tdata [61], \kme_cceip2_ob_out.tdata [60], 
	\kme_cceip2_ob_out.tdata [59], \kme_cceip2_ob_out.tdata [58], 
	\kme_cceip2_ob_out.tdata [57], \kme_cceip2_ob_out.tdata [56], 
	\kme_cceip2_ob_out.tdata [55], \kme_cceip2_ob_out.tdata [54], 
	\kme_cceip2_ob_out.tdata [53], \kme_cceip2_ob_out.tdata [52], 
	\kme_cceip2_ob_out.tdata [51], \kme_cceip2_ob_out.tdata [50], 
	\kme_cceip2_ob_out.tdata [49], \kme_cceip2_ob_out.tdata [48], 
	\kme_cceip2_ob_out.tdata [47], \kme_cceip2_ob_out.tdata [46], 
	\kme_cceip2_ob_out.tdata [45], \kme_cceip2_ob_out.tdata [44], 
	\kme_cceip2_ob_out.tdata [43], \kme_cceip2_ob_out.tdata [42], 
	\kme_cceip2_ob_out.tdata [41], \kme_cceip2_ob_out.tdata [40], 
	\kme_cceip2_ob_out.tdata [39], \kme_cceip2_ob_out.tdata [38], 
	\kme_cceip2_ob_out.tdata [37], \kme_cceip2_ob_out.tdata [36], 
	\kme_cceip2_ob_out.tdata [35], \kme_cceip2_ob_out.tdata [34], 
	\kme_cceip2_ob_out.tdata [33], \kme_cceip2_ob_out.tdata [32], 
	\kme_cceip2_ob_out.tdata [31], \kme_cceip2_ob_out.tdata [30], 
	\kme_cceip2_ob_out.tdata [29], \kme_cceip2_ob_out.tdata [28], 
	\kme_cceip2_ob_out.tdata [27], \kme_cceip2_ob_out.tdata [26], 
	\kme_cceip2_ob_out.tdata [25], \kme_cceip2_ob_out.tdata [24], 
	\kme_cceip2_ob_out.tdata [23], \kme_cceip2_ob_out.tdata [22], 
	\kme_cceip2_ob_out.tdata [21], \kme_cceip2_ob_out.tdata [20], 
	\kme_cceip2_ob_out.tdata [19], \kme_cceip2_ob_out.tdata [18], 
	\kme_cceip2_ob_out.tdata [17], \kme_cceip2_ob_out.tdata [16], 
	\kme_cceip2_ob_out.tdata [15], \kme_cceip2_ob_out.tdata [14], 
	\kme_cceip2_ob_out.tdata [13], \kme_cceip2_ob_out.tdata [12], 
	\kme_cceip2_ob_out.tdata [11], \kme_cceip2_ob_out.tdata [10], 
	\kme_cceip2_ob_out.tdata [9], \kme_cceip2_ob_out.tdata [8], 
	\kme_cceip2_ob_out.tdata [7], \kme_cceip2_ob_out.tdata [6], 
	\kme_cceip2_ob_out.tdata [5], \kme_cceip2_ob_out.tdata [4], 
	\kme_cceip2_ob_out.tdata [3], \kme_cceip2_ob_out.tdata [2], 
	\kme_cceip2_ob_out.tdata [1], \kme_cceip2_ob_out.tdata [0]} ), 
	.kme_cceip2_ob_in_mod( {\kme_cceip2_ob_in_mod.tready } ), 
	.kme_cceip3_ob_out( {\kme_cceip3_ob_out.tvalid , 
	\kme_cceip3_ob_out.tlast , \kme_cceip3_ob_out.tid [0], 
	\kme_cceip3_ob_out.tstrb [7], \kme_cceip3_ob_out.tstrb [6], 
	\kme_cceip3_ob_out.tstrb [5], \kme_cceip3_ob_out.tstrb [4], 
	\kme_cceip3_ob_out.tstrb [3], \kme_cceip3_ob_out.tstrb [2], 
	\kme_cceip3_ob_out.tstrb [1], \kme_cceip3_ob_out.tstrb [0], 
	\kme_cceip3_ob_out.tuser [7], \kme_cceip3_ob_out.tuser [6], 
	\kme_cceip3_ob_out.tuser [5], \kme_cceip3_ob_out.tuser [4], 
	\kme_cceip3_ob_out.tuser [3], \kme_cceip3_ob_out.tuser [2], 
	\kme_cceip3_ob_out.tuser [1], \kme_cceip3_ob_out.tuser [0], 
	\kme_cceip3_ob_out.tdata [63], \kme_cceip3_ob_out.tdata [62], 
	\kme_cceip3_ob_out.tdata [61], \kme_cceip3_ob_out.tdata [60], 
	\kme_cceip3_ob_out.tdata [59], \kme_cceip3_ob_out.tdata [58], 
	\kme_cceip3_ob_out.tdata [57], \kme_cceip3_ob_out.tdata [56], 
	\kme_cceip3_ob_out.tdata [55], \kme_cceip3_ob_out.tdata [54], 
	\kme_cceip3_ob_out.tdata [53], \kme_cceip3_ob_out.tdata [52], 
	\kme_cceip3_ob_out.tdata [51], \kme_cceip3_ob_out.tdata [50], 
	\kme_cceip3_ob_out.tdata [49], \kme_cceip3_ob_out.tdata [48], 
	\kme_cceip3_ob_out.tdata [47], \kme_cceip3_ob_out.tdata [46], 
	\kme_cceip3_ob_out.tdata [45], \kme_cceip3_ob_out.tdata [44], 
	\kme_cceip3_ob_out.tdata [43], \kme_cceip3_ob_out.tdata [42], 
	\kme_cceip3_ob_out.tdata [41], \kme_cceip3_ob_out.tdata [40], 
	\kme_cceip3_ob_out.tdata [39], \kme_cceip3_ob_out.tdata [38], 
	\kme_cceip3_ob_out.tdata [37], \kme_cceip3_ob_out.tdata [36], 
	\kme_cceip3_ob_out.tdata [35], \kme_cceip3_ob_out.tdata [34], 
	\kme_cceip3_ob_out.tdata [33], \kme_cceip3_ob_out.tdata [32], 
	\kme_cceip3_ob_out.tdata [31], \kme_cceip3_ob_out.tdata [30], 
	\kme_cceip3_ob_out.tdata [29], \kme_cceip3_ob_out.tdata [28], 
	\kme_cceip3_ob_out.tdata [27], \kme_cceip3_ob_out.tdata [26], 
	\kme_cceip3_ob_out.tdata [25], \kme_cceip3_ob_out.tdata [24], 
	\kme_cceip3_ob_out.tdata [23], \kme_cceip3_ob_out.tdata [22], 
	\kme_cceip3_ob_out.tdata [21], \kme_cceip3_ob_out.tdata [20], 
	\kme_cceip3_ob_out.tdata [19], \kme_cceip3_ob_out.tdata [18], 
	\kme_cceip3_ob_out.tdata [17], \kme_cceip3_ob_out.tdata [16], 
	\kme_cceip3_ob_out.tdata [15], \kme_cceip3_ob_out.tdata [14], 
	\kme_cceip3_ob_out.tdata [13], \kme_cceip3_ob_out.tdata [12], 
	\kme_cceip3_ob_out.tdata [11], \kme_cceip3_ob_out.tdata [10], 
	\kme_cceip3_ob_out.tdata [9], \kme_cceip3_ob_out.tdata [8], 
	\kme_cceip3_ob_out.tdata [7], \kme_cceip3_ob_out.tdata [6], 
	\kme_cceip3_ob_out.tdata [5], \kme_cceip3_ob_out.tdata [4], 
	\kme_cceip3_ob_out.tdata [3], \kme_cceip3_ob_out.tdata [2], 
	\kme_cceip3_ob_out.tdata [1], \kme_cceip3_ob_out.tdata [0]} ), 
	.kme_cceip3_ob_in_mod( {\kme_cceip3_ob_in_mod.tready } ), 
	.kme_cddip0_ob_out( {\kme_cddip0_ob_out.tvalid , 
	\kme_cddip0_ob_out.tlast , \kme_cddip0_ob_out.tid [0], 
	\kme_cddip0_ob_out.tstrb [7], \kme_cddip0_ob_out.tstrb [6], 
	\kme_cddip0_ob_out.tstrb [5], \kme_cddip0_ob_out.tstrb [4], 
	\kme_cddip0_ob_out.tstrb [3], \kme_cddip0_ob_out.tstrb [2], 
	\kme_cddip0_ob_out.tstrb [1], \kme_cddip0_ob_out.tstrb [0], 
	\kme_cddip0_ob_out.tuser [7], \kme_cddip0_ob_out.tuser [6], 
	\kme_cddip0_ob_out.tuser [5], \kme_cddip0_ob_out.tuser [4], 
	\kme_cddip0_ob_out.tuser [3], \kme_cddip0_ob_out.tuser [2], 
	\kme_cddip0_ob_out.tuser [1], \kme_cddip0_ob_out.tuser [0], 
	\kme_cddip0_ob_out.tdata [63], \kme_cddip0_ob_out.tdata [62], 
	\kme_cddip0_ob_out.tdata [61], \kme_cddip0_ob_out.tdata [60], 
	\kme_cddip0_ob_out.tdata [59], \kme_cddip0_ob_out.tdata [58], 
	\kme_cddip0_ob_out.tdata [57], \kme_cddip0_ob_out.tdata [56], 
	\kme_cddip0_ob_out.tdata [55], \kme_cddip0_ob_out.tdata [54], 
	\kme_cddip0_ob_out.tdata [53], \kme_cddip0_ob_out.tdata [52], 
	\kme_cddip0_ob_out.tdata [51], \kme_cddip0_ob_out.tdata [50], 
	\kme_cddip0_ob_out.tdata [49], \kme_cddip0_ob_out.tdata [48], 
	\kme_cddip0_ob_out.tdata [47], \kme_cddip0_ob_out.tdata [46], 
	\kme_cddip0_ob_out.tdata [45], \kme_cddip0_ob_out.tdata [44], 
	\kme_cddip0_ob_out.tdata [43], \kme_cddip0_ob_out.tdata [42], 
	\kme_cddip0_ob_out.tdata [41], \kme_cddip0_ob_out.tdata [40], 
	\kme_cddip0_ob_out.tdata [39], \kme_cddip0_ob_out.tdata [38], 
	\kme_cddip0_ob_out.tdata [37], \kme_cddip0_ob_out.tdata [36], 
	\kme_cddip0_ob_out.tdata [35], \kme_cddip0_ob_out.tdata [34], 
	\kme_cddip0_ob_out.tdata [33], \kme_cddip0_ob_out.tdata [32], 
	\kme_cddip0_ob_out.tdata [31], \kme_cddip0_ob_out.tdata [30], 
	\kme_cddip0_ob_out.tdata [29], \kme_cddip0_ob_out.tdata [28], 
	\kme_cddip0_ob_out.tdata [27], \kme_cddip0_ob_out.tdata [26], 
	\kme_cddip0_ob_out.tdata [25], \kme_cddip0_ob_out.tdata [24], 
	\kme_cddip0_ob_out.tdata [23], \kme_cddip0_ob_out.tdata [22], 
	\kme_cddip0_ob_out.tdata [21], \kme_cddip0_ob_out.tdata [20], 
	\kme_cddip0_ob_out.tdata [19], \kme_cddip0_ob_out.tdata [18], 
	\kme_cddip0_ob_out.tdata [17], \kme_cddip0_ob_out.tdata [16], 
	\kme_cddip0_ob_out.tdata [15], \kme_cddip0_ob_out.tdata [14], 
	\kme_cddip0_ob_out.tdata [13], \kme_cddip0_ob_out.tdata [12], 
	\kme_cddip0_ob_out.tdata [11], \kme_cddip0_ob_out.tdata [10], 
	\kme_cddip0_ob_out.tdata [9], \kme_cddip0_ob_out.tdata [8], 
	\kme_cddip0_ob_out.tdata [7], \kme_cddip0_ob_out.tdata [6], 
	\kme_cddip0_ob_out.tdata [5], \kme_cddip0_ob_out.tdata [4], 
	\kme_cddip0_ob_out.tdata [3], \kme_cddip0_ob_out.tdata [2], 
	\kme_cddip0_ob_out.tdata [1], \kme_cddip0_ob_out.tdata [0]} ), 
	.kme_cddip0_ob_in_mod( {\kme_cddip0_ob_in_mod.tready } ), 
	.kme_cddip1_ob_out( {\kme_cddip1_ob_out.tvalid , 
	\kme_cddip1_ob_out.tlast , \kme_cddip1_ob_out.tid [0], 
	\kme_cddip1_ob_out.tstrb [7], \kme_cddip1_ob_out.tstrb [6], 
	\kme_cddip1_ob_out.tstrb [5], \kme_cddip1_ob_out.tstrb [4], 
	\kme_cddip1_ob_out.tstrb [3], \kme_cddip1_ob_out.tstrb [2], 
	\kme_cddip1_ob_out.tstrb [1], \kme_cddip1_ob_out.tstrb [0], 
	\kme_cddip1_ob_out.tuser [7], \kme_cddip1_ob_out.tuser [6], 
	\kme_cddip1_ob_out.tuser [5], \kme_cddip1_ob_out.tuser [4], 
	\kme_cddip1_ob_out.tuser [3], \kme_cddip1_ob_out.tuser [2], 
	\kme_cddip1_ob_out.tuser [1], \kme_cddip1_ob_out.tuser [0], 
	\kme_cddip1_ob_out.tdata [63], \kme_cddip1_ob_out.tdata [62], 
	\kme_cddip1_ob_out.tdata [61], \kme_cddip1_ob_out.tdata [60], 
	\kme_cddip1_ob_out.tdata [59], \kme_cddip1_ob_out.tdata [58], 
	\kme_cddip1_ob_out.tdata [57], \kme_cddip1_ob_out.tdata [56], 
	\kme_cddip1_ob_out.tdata [55], \kme_cddip1_ob_out.tdata [54], 
	\kme_cddip1_ob_out.tdata [53], \kme_cddip1_ob_out.tdata [52], 
	\kme_cddip1_ob_out.tdata [51], \kme_cddip1_ob_out.tdata [50], 
	\kme_cddip1_ob_out.tdata [49], \kme_cddip1_ob_out.tdata [48], 
	\kme_cddip1_ob_out.tdata [47], \kme_cddip1_ob_out.tdata [46], 
	\kme_cddip1_ob_out.tdata [45], \kme_cddip1_ob_out.tdata [44], 
	\kme_cddip1_ob_out.tdata [43], \kme_cddip1_ob_out.tdata [42], 
	\kme_cddip1_ob_out.tdata [41], \kme_cddip1_ob_out.tdata [40], 
	\kme_cddip1_ob_out.tdata [39], \kme_cddip1_ob_out.tdata [38], 
	\kme_cddip1_ob_out.tdata [37], \kme_cddip1_ob_out.tdata [36], 
	\kme_cddip1_ob_out.tdata [35], \kme_cddip1_ob_out.tdata [34], 
	\kme_cddip1_ob_out.tdata [33], \kme_cddip1_ob_out.tdata [32], 
	\kme_cddip1_ob_out.tdata [31], \kme_cddip1_ob_out.tdata [30], 
	\kme_cddip1_ob_out.tdata [29], \kme_cddip1_ob_out.tdata [28], 
	\kme_cddip1_ob_out.tdata [27], \kme_cddip1_ob_out.tdata [26], 
	\kme_cddip1_ob_out.tdata [25], \kme_cddip1_ob_out.tdata [24], 
	\kme_cddip1_ob_out.tdata [23], \kme_cddip1_ob_out.tdata [22], 
	\kme_cddip1_ob_out.tdata [21], \kme_cddip1_ob_out.tdata [20], 
	\kme_cddip1_ob_out.tdata [19], \kme_cddip1_ob_out.tdata [18], 
	\kme_cddip1_ob_out.tdata [17], \kme_cddip1_ob_out.tdata [16], 
	\kme_cddip1_ob_out.tdata [15], \kme_cddip1_ob_out.tdata [14], 
	\kme_cddip1_ob_out.tdata [13], \kme_cddip1_ob_out.tdata [12], 
	\kme_cddip1_ob_out.tdata [11], \kme_cddip1_ob_out.tdata [10], 
	\kme_cddip1_ob_out.tdata [9], \kme_cddip1_ob_out.tdata [8], 
	\kme_cddip1_ob_out.tdata [7], \kme_cddip1_ob_out.tdata [6], 
	\kme_cddip1_ob_out.tdata [5], \kme_cddip1_ob_out.tdata [4], 
	\kme_cddip1_ob_out.tdata [3], \kme_cddip1_ob_out.tdata [2], 
	\kme_cddip1_ob_out.tdata [1], \kme_cddip1_ob_out.tdata [0]} ), 
	.kme_cddip1_ob_in_mod( {\kme_cddip1_ob_in_mod.tready } ), 
	.kme_cddip2_ob_out( {\kme_cddip2_ob_out.tvalid , 
	\kme_cddip2_ob_out.tlast , \kme_cddip2_ob_out.tid [0], 
	\kme_cddip2_ob_out.tstrb [7], \kme_cddip2_ob_out.tstrb [6], 
	\kme_cddip2_ob_out.tstrb [5], \kme_cddip2_ob_out.tstrb [4], 
	\kme_cddip2_ob_out.tstrb [3], \kme_cddip2_ob_out.tstrb [2], 
	\kme_cddip2_ob_out.tstrb [1], \kme_cddip2_ob_out.tstrb [0], 
	\kme_cddip2_ob_out.tuser [7], \kme_cddip2_ob_out.tuser [6], 
	\kme_cddip2_ob_out.tuser [5], \kme_cddip2_ob_out.tuser [4], 
	\kme_cddip2_ob_out.tuser [3], \kme_cddip2_ob_out.tuser [2], 
	\kme_cddip2_ob_out.tuser [1], \kme_cddip2_ob_out.tuser [0], 
	\kme_cddip2_ob_out.tdata [63], \kme_cddip2_ob_out.tdata [62], 
	\kme_cddip2_ob_out.tdata [61], \kme_cddip2_ob_out.tdata [60], 
	\kme_cddip2_ob_out.tdata [59], \kme_cddip2_ob_out.tdata [58], 
	\kme_cddip2_ob_out.tdata [57], \kme_cddip2_ob_out.tdata [56], 
	\kme_cddip2_ob_out.tdata [55], \kme_cddip2_ob_out.tdata [54], 
	\kme_cddip2_ob_out.tdata [53], \kme_cddip2_ob_out.tdata [52], 
	\kme_cddip2_ob_out.tdata [51], \kme_cddip2_ob_out.tdata [50], 
	\kme_cddip2_ob_out.tdata [49], \kme_cddip2_ob_out.tdata [48], 
	\kme_cddip2_ob_out.tdata [47], \kme_cddip2_ob_out.tdata [46], 
	\kme_cddip2_ob_out.tdata [45], \kme_cddip2_ob_out.tdata [44], 
	\kme_cddip2_ob_out.tdata [43], \kme_cddip2_ob_out.tdata [42], 
	\kme_cddip2_ob_out.tdata [41], \kme_cddip2_ob_out.tdata [40], 
	\kme_cddip2_ob_out.tdata [39], \kme_cddip2_ob_out.tdata [38], 
	\kme_cddip2_ob_out.tdata [37], \kme_cddip2_ob_out.tdata [36], 
	\kme_cddip2_ob_out.tdata [35], \kme_cddip2_ob_out.tdata [34], 
	\kme_cddip2_ob_out.tdata [33], \kme_cddip2_ob_out.tdata [32], 
	\kme_cddip2_ob_out.tdata [31], \kme_cddip2_ob_out.tdata [30], 
	\kme_cddip2_ob_out.tdata [29], \kme_cddip2_ob_out.tdata [28], 
	\kme_cddip2_ob_out.tdata [27], \kme_cddip2_ob_out.tdata [26], 
	\kme_cddip2_ob_out.tdata [25], \kme_cddip2_ob_out.tdata [24], 
	\kme_cddip2_ob_out.tdata [23], \kme_cddip2_ob_out.tdata [22], 
	\kme_cddip2_ob_out.tdata [21], \kme_cddip2_ob_out.tdata [20], 
	\kme_cddip2_ob_out.tdata [19], \kme_cddip2_ob_out.tdata [18], 
	\kme_cddip2_ob_out.tdata [17], \kme_cddip2_ob_out.tdata [16], 
	\kme_cddip2_ob_out.tdata [15], \kme_cddip2_ob_out.tdata [14], 
	\kme_cddip2_ob_out.tdata [13], \kme_cddip2_ob_out.tdata [12], 
	\kme_cddip2_ob_out.tdata [11], \kme_cddip2_ob_out.tdata [10], 
	\kme_cddip2_ob_out.tdata [9], \kme_cddip2_ob_out.tdata [8], 
	\kme_cddip2_ob_out.tdata [7], \kme_cddip2_ob_out.tdata [6], 
	\kme_cddip2_ob_out.tdata [5], \kme_cddip2_ob_out.tdata [4], 
	\kme_cddip2_ob_out.tdata [3], \kme_cddip2_ob_out.tdata [2], 
	\kme_cddip2_ob_out.tdata [1], \kme_cddip2_ob_out.tdata [0]} ), 
	.kme_cddip2_ob_in_mod( {\kme_cddip2_ob_in_mod.tready } ), 
	.kme_cddip3_ob_out( {\kme_cddip3_ob_out.tvalid , 
	\kme_cddip3_ob_out.tlast , \kme_cddip3_ob_out.tid [0], 
	\kme_cddip3_ob_out.tstrb [7], \kme_cddip3_ob_out.tstrb [6], 
	\kme_cddip3_ob_out.tstrb [5], \kme_cddip3_ob_out.tstrb [4], 
	\kme_cddip3_ob_out.tstrb [3], \kme_cddip3_ob_out.tstrb [2], 
	\kme_cddip3_ob_out.tstrb [1], \kme_cddip3_ob_out.tstrb [0], 
	\kme_cddip3_ob_out.tuser [7], \kme_cddip3_ob_out.tuser [6], 
	\kme_cddip3_ob_out.tuser [5], \kme_cddip3_ob_out.tuser [4], 
	\kme_cddip3_ob_out.tuser [3], \kme_cddip3_ob_out.tuser [2], 
	\kme_cddip3_ob_out.tuser [1], \kme_cddip3_ob_out.tuser [0], 
	\kme_cddip3_ob_out.tdata [63], \kme_cddip3_ob_out.tdata [62], 
	\kme_cddip3_ob_out.tdata [61], \kme_cddip3_ob_out.tdata [60], 
	\kme_cddip3_ob_out.tdata [59], \kme_cddip3_ob_out.tdata [58], 
	\kme_cddip3_ob_out.tdata [57], \kme_cddip3_ob_out.tdata [56], 
	\kme_cddip3_ob_out.tdata [55], \kme_cddip3_ob_out.tdata [54], 
	\kme_cddip3_ob_out.tdata [53], \kme_cddip3_ob_out.tdata [52], 
	\kme_cddip3_ob_out.tdata [51], \kme_cddip3_ob_out.tdata [50], 
	\kme_cddip3_ob_out.tdata [49], \kme_cddip3_ob_out.tdata [48], 
	\kme_cddip3_ob_out.tdata [47], \kme_cddip3_ob_out.tdata [46], 
	\kme_cddip3_ob_out.tdata [45], \kme_cddip3_ob_out.tdata [44], 
	\kme_cddip3_ob_out.tdata [43], \kme_cddip3_ob_out.tdata [42], 
	\kme_cddip3_ob_out.tdata [41], \kme_cddip3_ob_out.tdata [40], 
	\kme_cddip3_ob_out.tdata [39], \kme_cddip3_ob_out.tdata [38], 
	\kme_cddip3_ob_out.tdata [37], \kme_cddip3_ob_out.tdata [36], 
	\kme_cddip3_ob_out.tdata [35], \kme_cddip3_ob_out.tdata [34], 
	\kme_cddip3_ob_out.tdata [33], \kme_cddip3_ob_out.tdata [32], 
	\kme_cddip3_ob_out.tdata [31], \kme_cddip3_ob_out.tdata [30], 
	\kme_cddip3_ob_out.tdata [29], \kme_cddip3_ob_out.tdata [28], 
	\kme_cddip3_ob_out.tdata [27], \kme_cddip3_ob_out.tdata [26], 
	\kme_cddip3_ob_out.tdata [25], \kme_cddip3_ob_out.tdata [24], 
	\kme_cddip3_ob_out.tdata [23], \kme_cddip3_ob_out.tdata [22], 
	\kme_cddip3_ob_out.tdata [21], \kme_cddip3_ob_out.tdata [20], 
	\kme_cddip3_ob_out.tdata [19], \kme_cddip3_ob_out.tdata [18], 
	\kme_cddip3_ob_out.tdata [17], \kme_cddip3_ob_out.tdata [16], 
	\kme_cddip3_ob_out.tdata [15], \kme_cddip3_ob_out.tdata [14], 
	\kme_cddip3_ob_out.tdata [13], \kme_cddip3_ob_out.tdata [12], 
	\kme_cddip3_ob_out.tdata [11], \kme_cddip3_ob_out.tdata [10], 
	\kme_cddip3_ob_out.tdata [9], \kme_cddip3_ob_out.tdata [8], 
	\kme_cddip3_ob_out.tdata [7], \kme_cddip3_ob_out.tdata [6], 
	\kme_cddip3_ob_out.tdata [5], \kme_cddip3_ob_out.tdata [4], 
	\kme_cddip3_ob_out.tdata [3], \kme_cddip3_ob_out.tdata [2], 
	\kme_cddip3_ob_out.tdata [1], \kme_cddip3_ob_out.tdata [0]} ), 
	.kme_cddip3_ob_in_mod( {\kme_cddip3_ob_in_mod.tready } ), ckv_dout, 
	ckv_mbe, .kim_dout( {\kim_dout.valid [0], \kim_dout.label_index [2], 
	\kim_dout.label_index [1], \kim_dout.label_index [0], 
	\kim_dout.ckv_length [1], \kim_dout.ckv_length [0], 
	\kim_dout.ckv_pointer [14], \kim_dout.ckv_pointer [13], 
	\kim_dout.ckv_pointer [12], \kim_dout.ckv_pointer [11], 
	\kim_dout.ckv_pointer [10], \kim_dout.ckv_pointer [9], 
	\kim_dout.ckv_pointer [8], \kim_dout.ckv_pointer [7], 
	\kim_dout.ckv_pointer [6], \kim_dout.ckv_pointer [5], 
	\kim_dout.ckv_pointer [4], \kim_dout.ckv_pointer [3], 
	\kim_dout.ckv_pointer [2], \kim_dout.ckv_pointer [1], 
	\kim_dout.ckv_pointer [0], \kim_dout.pf_num [3], 
	\kim_dout.pf_num [2], \kim_dout.pf_num [1], \kim_dout.pf_num [0], 
	\kim_dout.vf_num [11], \kim_dout.vf_num [10], \kim_dout.vf_num [9], 
	\kim_dout.vf_num [8], \kim_dout.vf_num [7], \kim_dout.vf_num [6], 
	\kim_dout.vf_num [5], \kim_dout.vf_num [4], \kim_dout.vf_num [3], 
	\kim_dout.vf_num [2], \kim_dout.vf_num [1], \kim_dout.vf_num [0], 
	\kim_dout.vf_valid [0]} ), kim_mbe, bimc_rst_n, 
	cceip_encrypt_bimc_isync, cceip_encrypt_bimc_idat, 
	cceip_validate_bimc_isync, cceip_validate_bimc_idat, 
	cddip_decrypt_bimc_isync, cddip_decrypt_bimc_idat, axi_bimc_isync, 
	axi_bimc_idat, .labels( {\labels[7].guid_size[0] , 
	\labels[7].label_size[5] , \labels[7].label_size[4] , 
	\labels[7].label_size[3] , \labels[7].label_size[2] , 
	\labels[7].label_size[1] , \labels[7].label_size[0] , 
	\labels[7].label[255] , \labels[7].label[254] , 
	\labels[7].label[253] , \labels[7].label[252] , 
	\labels[7].label[251] , \labels[7].label[250] , 
	\labels[7].label[249] , \labels[7].label[248] , 
	\labels[7].label[247] , \labels[7].label[246] , 
	\labels[7].label[245] , \labels[7].label[244] , 
	\labels[7].label[243] , \labels[7].label[242] , 
	\labels[7].label[241] , \labels[7].label[240] , 
	\labels[7].label[239] , \labels[7].label[238] , 
	\labels[7].label[237] , \labels[7].label[236] , 
	\labels[7].label[235] , \labels[7].label[234] , 
	\labels[7].label[233] , \labels[7].label[232] , 
	\labels[7].label[231] , \labels[7].label[230] , 
	\labels[7].label[229] , \labels[7].label[228] , 
	\labels[7].label[227] , \labels[7].label[226] , 
	\labels[7].label[225] , \labels[7].label[224] , 
	\labels[7].label[223] , \labels[7].label[222] , 
	\labels[7].label[221] , \labels[7].label[220] , 
	\labels[7].label[219] , \labels[7].label[218] , 
	\labels[7].label[217] , \labels[7].label[216] , 
	\labels[7].label[215] , \labels[7].label[214] , 
	\labels[7].label[213] , \labels[7].label[212] , 
	\labels[7].label[211] , \labels[7].label[210] , 
	\labels[7].label[209] , \labels[7].label[208] , 
	\labels[7].label[207] , \labels[7].label[206] , 
	\labels[7].label[205] , \labels[7].label[204] , 
	\labels[7].label[203] , \labels[7].label[202] , 
	\labels[7].label[201] , \labels[7].label[200] , 
	\labels[7].label[199] , \labels[7].label[198] , 
	\labels[7].label[197] , \labels[7].label[196] , 
	\labels[7].label[195] , \labels[7].label[194] , 
	\labels[7].label[193] , \labels[7].label[192] , 
	\labels[7].label[191] , \labels[7].label[190] , 
	\labels[7].label[189] , \labels[7].label[188] , 
	\labels[7].label[187] , \labels[7].label[186] , 
	\labels[7].label[185] , \labels[7].label[184] , 
	\labels[7].label[183] , \labels[7].label[182] , 
	\labels[7].label[181] , \labels[7].label[180] , 
	\labels[7].label[179] , \labels[7].label[178] , 
	\labels[7].label[177] , \labels[7].label[176] , 
	\labels[7].label[175] , \labels[7].label[174] , 
	\labels[7].label[173] , \labels[7].label[172] , 
	\labels[7].label[171] , \labels[7].label[170] , 
	\labels[7].label[169] , \labels[7].label[168] , 
	\labels[7].label[167] , \labels[7].label[166] , 
	\labels[7].label[165] , \labels[7].label[164] , 
	\labels[7].label[163] , \labels[7].label[162] , 
	\labels[7].label[161] , \labels[7].label[160] , 
	\labels[7].label[159] , \labels[7].label[158] , 
	\labels[7].label[157] , \labels[7].label[156] , 
	\labels[7].label[155] , \labels[7].label[154] , 
	\labels[7].label[153] , \labels[7].label[152] , 
	\labels[7].label[151] , \labels[7].label[150] , 
	\labels[7].label[149] , \labels[7].label[148] , 
	\labels[7].label[147] , \labels[7].label[146] , 
	\labels[7].label[145] , \labels[7].label[144] , 
	\labels[7].label[143] , \labels[7].label[142] , 
	\labels[7].label[141] , \labels[7].label[140] , 
	\labels[7].label[139] , \labels[7].label[138] , 
	\labels[7].label[137] , \labels[7].label[136] , 
	\labels[7].label[135] , \labels[7].label[134] , 
	\labels[7].label[133] , \labels[7].label[132] , 
	\labels[7].label[131] , \labels[7].label[130] , 
	\labels[7].label[129] , \labels[7].label[128] , 
	\labels[7].label[127] , \labels[7].label[126] , 
	\labels[7].label[125] , \labels[7].label[124] , 
	\labels[7].label[123] , \labels[7].label[122] , 
	\labels[7].label[121] , \labels[7].label[120] , 
	\labels[7].label[119] , \labels[7].label[118] , 
	\labels[7].label[117] , \labels[7].label[116] , 
	\labels[7].label[115] , \labels[7].label[114] , 
	\labels[7].label[113] , \labels[7].label[112] , 
	\labels[7].label[111] , \labels[7].label[110] , 
	\labels[7].label[109] , \labels[7].label[108] , 
	\labels[7].label[107] , \labels[7].label[106] , 
	\labels[7].label[105] , \labels[7].label[104] , 
	\labels[7].label[103] , \labels[7].label[102] , 
	\labels[7].label[101] , \labels[7].label[100] , 
	\labels[7].label[99] , \labels[7].label[98] , \labels[7].label[97] , 
	\labels[7].label[96] , \labels[7].label[95] , \labels[7].label[94] , 
	\labels[7].label[93] , \labels[7].label[92] , \labels[7].label[91] , 
	\labels[7].label[90] , \labels[7].label[89] , \labels[7].label[88] , 
	\labels[7].label[87] , \labels[7].label[86] , \labels[7].label[85] , 
	\labels[7].label[84] , \labels[7].label[83] , \labels[7].label[82] , 
	\labels[7].label[81] , \labels[7].label[80] , \labels[7].label[79] , 
	\labels[7].label[78] , \labels[7].label[77] , \labels[7].label[76] , 
	\labels[7].label[75] , \labels[7].label[74] , \labels[7].label[73] , 
	\labels[7].label[72] , \labels[7].label[71] , \labels[7].label[70] , 
	\labels[7].label[69] , \labels[7].label[68] , \labels[7].label[67] , 
	\labels[7].label[66] , \labels[7].label[65] , \labels[7].label[64] , 
	\labels[7].label[63] , \labels[7].label[62] , \labels[7].label[61] , 
	\labels[7].label[60] , \labels[7].label[59] , \labels[7].label[58] , 
	\labels[7].label[57] , \labels[7].label[56] , \labels[7].label[55] , 
	\labels[7].label[54] , \labels[7].label[53] , \labels[7].label[52] , 
	\labels[7].label[51] , \labels[7].label[50] , \labels[7].label[49] , 
	\labels[7].label[48] , \labels[7].label[47] , \labels[7].label[46] , 
	\labels[7].label[45] , \labels[7].label[44] , \labels[7].label[43] , 
	\labels[7].label[42] , \labels[7].label[41] , \labels[7].label[40] , 
	\labels[7].label[39] , \labels[7].label[38] , \labels[7].label[37] , 
	\labels[7].label[36] , \labels[7].label[35] , \labels[7].label[34] , 
	\labels[7].label[33] , \labels[7].label[32] , \labels[7].label[31] , 
	\labels[7].label[30] , \labels[7].label[29] , \labels[7].label[28] , 
	\labels[7].label[27] , \labels[7].label[26] , \labels[7].label[25] , 
	\labels[7].label[24] , \labels[7].label[23] , \labels[7].label[22] , 
	\labels[7].label[21] , \labels[7].label[20] , \labels[7].label[19] , 
	\labels[7].label[18] , \labels[7].label[17] , \labels[7].label[16] , 
	\labels[7].label[15] , \labels[7].label[14] , \labels[7].label[13] , 
	\labels[7].label[12] , \labels[7].label[11] , \labels[7].label[10] , 
	\labels[7].label[9] , \labels[7].label[8] , \labels[7].label[7] , 
	\labels[7].label[6] , \labels[7].label[5] , \labels[7].label[4] , 
	\labels[7].label[3] , \labels[7].label[2] , \labels[7].label[1] , 
	\labels[7].label[0] , \labels[7].delimiter_valid[0] , 
	\labels[7].delimiter[7] , \labels[7].delimiter[6] , 
	\labels[7].delimiter[5] , \labels[7].delimiter[4] , 
	\labels[7].delimiter[3] , \labels[7].delimiter[2] , 
	\labels[7].delimiter[1] , \labels[7].delimiter[0] , 
	\labels[6].guid_size[0] , \labels[6].label_size[5] , 
	\labels[6].label_size[4] , \labels[6].label_size[3] , 
	\labels[6].label_size[2] , \labels[6].label_size[1] , 
	\labels[6].label_size[0] , \labels[6].label[255] , 
	\labels[6].label[254] , \labels[6].label[253] , 
	\labels[6].label[252] , \labels[6].label[251] , 
	\labels[6].label[250] , \labels[6].label[249] , 
	\labels[6].label[248] , \labels[6].label[247] , 
	\labels[6].label[246] , \labels[6].label[245] , 
	\labels[6].label[244] , \labels[6].label[243] , 
	\labels[6].label[242] , \labels[6].label[241] , 
	\labels[6].label[240] , \labels[6].label[239] , 
	\labels[6].label[238] , \labels[6].label[237] , 
	\labels[6].label[236] , \labels[6].label[235] , 
	\labels[6].label[234] , \labels[6].label[233] , 
	\labels[6].label[232] , \labels[6].label[231] , 
	\labels[6].label[230] , \labels[6].label[229] , 
	\labels[6].label[228] , \labels[6].label[227] , 
	\labels[6].label[226] , \labels[6].label[225] , 
	\labels[6].label[224] , \labels[6].label[223] , 
	\labels[6].label[222] , \labels[6].label[221] , 
	\labels[6].label[220] , \labels[6].label[219] , 
	\labels[6].label[218] , \labels[6].label[217] , 
	\labels[6].label[216] , \labels[6].label[215] , 
	\labels[6].label[214] , \labels[6].label[213] , 
	\labels[6].label[212] , \labels[6].label[211] , 
	\labels[6].label[210] , \labels[6].label[209] , 
	\labels[6].label[208] , \labels[6].label[207] , 
	\labels[6].label[206] , \labels[6].label[205] , 
	\labels[6].label[204] , \labels[6].label[203] , 
	\labels[6].label[202] , \labels[6].label[201] , 
	\labels[6].label[200] , \labels[6].label[199] , 
	\labels[6].label[198] , \labels[6].label[197] , 
	\labels[6].label[196] , \labels[6].label[195] , 
	\labels[6].label[194] , \labels[6].label[193] , 
	\labels[6].label[192] , \labels[6].label[191] , 
	\labels[6].label[190] , \labels[6].label[189] , 
	\labels[6].label[188] , \labels[6].label[187] , 
	\labels[6].label[186] , \labels[6].label[185] , 
	\labels[6].label[184] , \labels[6].label[183] , 
	\labels[6].label[182] , \labels[6].label[181] , 
	\labels[6].label[180] , \labels[6].label[179] , 
	\labels[6].label[178] , \labels[6].label[177] , 
	\labels[6].label[176] , \labels[6].label[175] , 
	\labels[6].label[174] , \labels[6].label[173] , 
	\labels[6].label[172] , \labels[6].label[171] , 
	\labels[6].label[170] , \labels[6].label[169] , 
	\labels[6].label[168] , \labels[6].label[167] , 
	\labels[6].label[166] , \labels[6].label[165] , 
	\labels[6].label[164] , \labels[6].label[163] , 
	\labels[6].label[162] , \labels[6].label[161] , 
	\labels[6].label[160] , \labels[6].label[159] , 
	\labels[6].label[158] , \labels[6].label[157] , 
	\labels[6].label[156] , \labels[6].label[155] , 
	\labels[6].label[154] , \labels[6].label[153] , 
	\labels[6].label[152] , \labels[6].label[151] , 
	\labels[6].label[150] , \labels[6].label[149] , 
	\labels[6].label[148] , \labels[6].label[147] , 
	\labels[6].label[146] , \labels[6].label[145] , 
	\labels[6].label[144] , \labels[6].label[143] , 
	\labels[6].label[142] , \labels[6].label[141] , 
	\labels[6].label[140] , \labels[6].label[139] , 
	\labels[6].label[138] , \labels[6].label[137] , 
	\labels[6].label[136] , \labels[6].label[135] , 
	\labels[6].label[134] , \labels[6].label[133] , 
	\labels[6].label[132] , \labels[6].label[131] , 
	\labels[6].label[130] , \labels[6].label[129] , 
	\labels[6].label[128] , \labels[6].label[127] , 
	\labels[6].label[126] , \labels[6].label[125] , 
	\labels[6].label[124] , \labels[6].label[123] , 
	\labels[6].label[122] , \labels[6].label[121] , 
	\labels[6].label[120] , \labels[6].label[119] , 
	\labels[6].label[118] , \labels[6].label[117] , 
	\labels[6].label[116] , \labels[6].label[115] , 
	\labels[6].label[114] , \labels[6].label[113] , 
	\labels[6].label[112] , \labels[6].label[111] , 
	\labels[6].label[110] , \labels[6].label[109] , 
	\labels[6].label[108] , \labels[6].label[107] , 
	\labels[6].label[106] , \labels[6].label[105] , 
	\labels[6].label[104] , \labels[6].label[103] , 
	\labels[6].label[102] , \labels[6].label[101] , 
	\labels[6].label[100] , \labels[6].label[99] , \labels[6].label[98] , 
	\labels[6].label[97] , \labels[6].label[96] , \labels[6].label[95] , 
	\labels[6].label[94] , \labels[6].label[93] , \labels[6].label[92] , 
	\labels[6].label[91] , \labels[6].label[90] , \labels[6].label[89] , 
	\labels[6].label[88] , \labels[6].label[87] , \labels[6].label[86] , 
	\labels[6].label[85] , \labels[6].label[84] , \labels[6].label[83] , 
	\labels[6].label[82] , \labels[6].label[81] , \labels[6].label[80] , 
	\labels[6].label[79] , \labels[6].label[78] , \labels[6].label[77] , 
	\labels[6].label[76] , \labels[6].label[75] , \labels[6].label[74] , 
	\labels[6].label[73] , \labels[6].label[72] , \labels[6].label[71] , 
	\labels[6].label[70] , \labels[6].label[69] , \labels[6].label[68] , 
	\labels[6].label[67] , \labels[6].label[66] , \labels[6].label[65] , 
	\labels[6].label[64] , \labels[6].label[63] , \labels[6].label[62] , 
	\labels[6].label[61] , \labels[6].label[60] , \labels[6].label[59] , 
	\labels[6].label[58] , \labels[6].label[57] , \labels[6].label[56] , 
	\labels[6].label[55] , \labels[6].label[54] , \labels[6].label[53] , 
	\labels[6].label[52] , \labels[6].label[51] , \labels[6].label[50] , 
	\labels[6].label[49] , \labels[6].label[48] , \labels[6].label[47] , 
	\labels[6].label[46] , \labels[6].label[45] , \labels[6].label[44] , 
	\labels[6].label[43] , \labels[6].label[42] , \labels[6].label[41] , 
	\labels[6].label[40] , \labels[6].label[39] , \labels[6].label[38] , 
	\labels[6].label[37] , \labels[6].label[36] , \labels[6].label[35] , 
	\labels[6].label[34] , \labels[6].label[33] , \labels[6].label[32] , 
	\labels[6].label[31] , \labels[6].label[30] , \labels[6].label[29] , 
	\labels[6].label[28] , \labels[6].label[27] , \labels[6].label[26] , 
	\labels[6].label[25] , \labels[6].label[24] , \labels[6].label[23] , 
	\labels[6].label[22] , \labels[6].label[21] , \labels[6].label[20] , 
	\labels[6].label[19] , \labels[6].label[18] , \labels[6].label[17] , 
	\labels[6].label[16] , \labels[6].label[15] , \labels[6].label[14] , 
	\labels[6].label[13] , \labels[6].label[12] , \labels[6].label[11] , 
	\labels[6].label[10] , \labels[6].label[9] , \labels[6].label[8] , 
	\labels[6].label[7] , \labels[6].label[6] , \labels[6].label[5] , 
	\labels[6].label[4] , \labels[6].label[3] , \labels[6].label[2] , 
	\labels[6].label[1] , \labels[6].label[0] , 
	\labels[6].delimiter_valid[0] , \labels[6].delimiter[7] , 
	\labels[6].delimiter[6] , \labels[6].delimiter[5] , 
	\labels[6].delimiter[4] , \labels[6].delimiter[3] , 
	\labels[6].delimiter[2] , \labels[6].delimiter[1] , 
	\labels[6].delimiter[0] , \labels[5].guid_size[0] , 
	\labels[5].label_size[5] , \labels[5].label_size[4] , 
	\labels[5].label_size[3] , \labels[5].label_size[2] , 
	\labels[5].label_size[1] , \labels[5].label_size[0] , 
	\labels[5].label[255] , \labels[5].label[254] , 
	\labels[5].label[253] , \labels[5].label[252] , 
	\labels[5].label[251] , \labels[5].label[250] , 
	\labels[5].label[249] , \labels[5].label[248] , 
	\labels[5].label[247] , \labels[5].label[246] , 
	\labels[5].label[245] , \labels[5].label[244] , 
	\labels[5].label[243] , \labels[5].label[242] , 
	\labels[5].label[241] , \labels[5].label[240] , 
	\labels[5].label[239] , \labels[5].label[238] , 
	\labels[5].label[237] , \labels[5].label[236] , 
	\labels[5].label[235] , \labels[5].label[234] , 
	\labels[5].label[233] , \labels[5].label[232] , 
	\labels[5].label[231] , \labels[5].label[230] , 
	\labels[5].label[229] , \labels[5].label[228] , 
	\labels[5].label[227] , \labels[5].label[226] , 
	\labels[5].label[225] , \labels[5].label[224] , 
	\labels[5].label[223] , \labels[5].label[222] , 
	\labels[5].label[221] , \labels[5].label[220] , 
	\labels[5].label[219] , \labels[5].label[218] , 
	\labels[5].label[217] , \labels[5].label[216] , 
	\labels[5].label[215] , \labels[5].label[214] , 
	\labels[5].label[213] , \labels[5].label[212] , 
	\labels[5].label[211] , \labels[5].label[210] , 
	\labels[5].label[209] , \labels[5].label[208] , 
	\labels[5].label[207] , \labels[5].label[206] , 
	\labels[5].label[205] , \labels[5].label[204] , 
	\labels[5].label[203] , \labels[5].label[202] , 
	\labels[5].label[201] , \labels[5].label[200] , 
	\labels[5].label[199] , \labels[5].label[198] , 
	\labels[5].label[197] , \labels[5].label[196] , 
	\labels[5].label[195] , \labels[5].label[194] , 
	\labels[5].label[193] , \labels[5].label[192] , 
	\labels[5].label[191] , \labels[5].label[190] , 
	\labels[5].label[189] , \labels[5].label[188] , 
	\labels[5].label[187] , \labels[5].label[186] , 
	\labels[5].label[185] , \labels[5].label[184] , 
	\labels[5].label[183] , \labels[5].label[182] , 
	\labels[5].label[181] , \labels[5].label[180] , 
	\labels[5].label[179] , \labels[5].label[178] , 
	\labels[5].label[177] , \labels[5].label[176] , 
	\labels[5].label[175] , \labels[5].label[174] , 
	\labels[5].label[173] , \labels[5].label[172] , 
	\labels[5].label[171] , \labels[5].label[170] , 
	\labels[5].label[169] , \labels[5].label[168] , 
	\labels[5].label[167] , \labels[5].label[166] , 
	\labels[5].label[165] , \labels[5].label[164] , 
	\labels[5].label[163] , \labels[5].label[162] , 
	\labels[5].label[161] , \labels[5].label[160] , 
	\labels[5].label[159] , \labels[5].label[158] , 
	\labels[5].label[157] , \labels[5].label[156] , 
	\labels[5].label[155] , \labels[5].label[154] , 
	\labels[5].label[153] , \labels[5].label[152] , 
	\labels[5].label[151] , \labels[5].label[150] , 
	\labels[5].label[149] , \labels[5].label[148] , 
	\labels[5].label[147] , \labels[5].label[146] , 
	\labels[5].label[145] , \labels[5].label[144] , 
	\labels[5].label[143] , \labels[5].label[142] , 
	\labels[5].label[141] , \labels[5].label[140] , 
	\labels[5].label[139] , \labels[5].label[138] , 
	\labels[5].label[137] , \labels[5].label[136] , 
	\labels[5].label[135] , \labels[5].label[134] , 
	\labels[5].label[133] , \labels[5].label[132] , 
	\labels[5].label[131] , \labels[5].label[130] , 
	\labels[5].label[129] , \labels[5].label[128] , 
	\labels[5].label[127] , \labels[5].label[126] , 
	\labels[5].label[125] , \labels[5].label[124] , 
	\labels[5].label[123] , \labels[5].label[122] , 
	\labels[5].label[121] , \labels[5].label[120] , 
	\labels[5].label[119] , \labels[5].label[118] , 
	\labels[5].label[117] , \labels[5].label[116] , 
	\labels[5].label[115] , \labels[5].label[114] , 
	\labels[5].label[113] , \labels[5].label[112] , 
	\labels[5].label[111] , \labels[5].label[110] , 
	\labels[5].label[109] , \labels[5].label[108] , 
	\labels[5].label[107] , \labels[5].label[106] , 
	\labels[5].label[105] , \labels[5].label[104] , 
	\labels[5].label[103] , \labels[5].label[102] , 
	\labels[5].label[101] , \labels[5].label[100] , 
	\labels[5].label[99] , \labels[5].label[98] , \labels[5].label[97] , 
	\labels[5].label[96] , \labels[5].label[95] , \labels[5].label[94] , 
	\labels[5].label[93] , \labels[5].label[92] , \labels[5].label[91] , 
	\labels[5].label[90] , \labels[5].label[89] , \labels[5].label[88] , 
	\labels[5].label[87] , \labels[5].label[86] , \labels[5].label[85] , 
	\labels[5].label[84] , \labels[5].label[83] , \labels[5].label[82] , 
	\labels[5].label[81] , \labels[5].label[80] , \labels[5].label[79] , 
	\labels[5].label[78] , \labels[5].label[77] , \labels[5].label[76] , 
	\labels[5].label[75] , \labels[5].label[74] , \labels[5].label[73] , 
	\labels[5].label[72] , \labels[5].label[71] , \labels[5].label[70] , 
	\labels[5].label[69] , \labels[5].label[68] , \labels[5].label[67] , 
	\labels[5].label[66] , \labels[5].label[65] , \labels[5].label[64] , 
	\labels[5].label[63] , \labels[5].label[62] , \labels[5].label[61] , 
	\labels[5].label[60] , \labels[5].label[59] , \labels[5].label[58] , 
	\labels[5].label[57] , \labels[5].label[56] , \labels[5].label[55] , 
	\labels[5].label[54] , \labels[5].label[53] , \labels[5].label[52] , 
	\labels[5].label[51] , \labels[5].label[50] , \labels[5].label[49] , 
	\labels[5].label[48] , \labels[5].label[47] , \labels[5].label[46] , 
	\labels[5].label[45] , \labels[5].label[44] , \labels[5].label[43] , 
	\labels[5].label[42] , \labels[5].label[41] , \labels[5].label[40] , 
	\labels[5].label[39] , \labels[5].label[38] , \labels[5].label[37] , 
	\labels[5].label[36] , \labels[5].label[35] , \labels[5].label[34] , 
	\labels[5].label[33] , \labels[5].label[32] , \labels[5].label[31] , 
	\labels[5].label[30] , \labels[5].label[29] , \labels[5].label[28] , 
	\labels[5].label[27] , \labels[5].label[26] , \labels[5].label[25] , 
	\labels[5].label[24] , \labels[5].label[23] , \labels[5].label[22] , 
	\labels[5].label[21] , \labels[5].label[20] , \labels[5].label[19] , 
	\labels[5].label[18] , \labels[5].label[17] , \labels[5].label[16] , 
	\labels[5].label[15] , \labels[5].label[14] , \labels[5].label[13] , 
	\labels[5].label[12] , \labels[5].label[11] , \labels[5].label[10] , 
	\labels[5].label[9] , \labels[5].label[8] , \labels[5].label[7] , 
	\labels[5].label[6] , \labels[5].label[5] , \labels[5].label[4] , 
	\labels[5].label[3] , \labels[5].label[2] , \labels[5].label[1] , 
	\labels[5].label[0] , \labels[5].delimiter_valid[0] , 
	\labels[5].delimiter[7] , \labels[5].delimiter[6] , 
	\labels[5].delimiter[5] , \labels[5].delimiter[4] , 
	\labels[5].delimiter[3] , \labels[5].delimiter[2] , 
	\labels[5].delimiter[1] , \labels[5].delimiter[0] , 
	\labels[4].guid_size[0] , \labels[4].label_size[5] , 
	\labels[4].label_size[4] , \labels[4].label_size[3] , 
	\labels[4].label_size[2] , \labels[4].label_size[1] , 
	\labels[4].label_size[0] , \labels[4].label[255] , 
	\labels[4].label[254] , \labels[4].label[253] , 
	\labels[4].label[252] , \labels[4].label[251] , 
	\labels[4].label[250] , \labels[4].label[249] , 
	\labels[4].label[248] , \labels[4].label[247] , 
	\labels[4].label[246] , \labels[4].label[245] , 
	\labels[4].label[244] , \labels[4].label[243] , 
	\labels[4].label[242] , \labels[4].label[241] , 
	\labels[4].label[240] , \labels[4].label[239] , 
	\labels[4].label[238] , \labels[4].label[237] , 
	\labels[4].label[236] , \labels[4].label[235] , 
	\labels[4].label[234] , \labels[4].label[233] , 
	\labels[4].label[232] , \labels[4].label[231] , 
	\labels[4].label[230] , \labels[4].label[229] , 
	\labels[4].label[228] , \labels[4].label[227] , 
	\labels[4].label[226] , \labels[4].label[225] , 
	\labels[4].label[224] , \labels[4].label[223] , 
	\labels[4].label[222] , \labels[4].label[221] , 
	\labels[4].label[220] , \labels[4].label[219] , 
	\labels[4].label[218] , \labels[4].label[217] , 
	\labels[4].label[216] , \labels[4].label[215] , 
	\labels[4].label[214] , \labels[4].label[213] , 
	\labels[4].label[212] , \labels[4].label[211] , 
	\labels[4].label[210] , \labels[4].label[209] , 
	\labels[4].label[208] , \labels[4].label[207] , 
	\labels[4].label[206] , \labels[4].label[205] , 
	\labels[4].label[204] , \labels[4].label[203] , 
	\labels[4].label[202] , \labels[4].label[201] , 
	\labels[4].label[200] , \labels[4].label[199] , 
	\labels[4].label[198] , \labels[4].label[197] , 
	\labels[4].label[196] , \labels[4].label[195] , 
	\labels[4].label[194] , \labels[4].label[193] , 
	\labels[4].label[192] , \labels[4].label[191] , 
	\labels[4].label[190] , \labels[4].label[189] , 
	\labels[4].label[188] , \labels[4].label[187] , 
	\labels[4].label[186] , \labels[4].label[185] , 
	\labels[4].label[184] , \labels[4].label[183] , 
	\labels[4].label[182] , \labels[4].label[181] , 
	\labels[4].label[180] , \labels[4].label[179] , 
	\labels[4].label[178] , \labels[4].label[177] , 
	\labels[4].label[176] , \labels[4].label[175] , 
	\labels[4].label[174] , \labels[4].label[173] , 
	\labels[4].label[172] , \labels[4].label[171] , 
	\labels[4].label[170] , \labels[4].label[169] , 
	\labels[4].label[168] , \labels[4].label[167] , 
	\labels[4].label[166] , \labels[4].label[165] , 
	\labels[4].label[164] , \labels[4].label[163] , 
	\labels[4].label[162] , \labels[4].label[161] , 
	\labels[4].label[160] , \labels[4].label[159] , 
	\labels[4].label[158] , \labels[4].label[157] , 
	\labels[4].label[156] , \labels[4].label[155] , 
	\labels[4].label[154] , \labels[4].label[153] , 
	\labels[4].label[152] , \labels[4].label[151] , 
	\labels[4].label[150] , \labels[4].label[149] , 
	\labels[4].label[148] , \labels[4].label[147] , 
	\labels[4].label[146] , \labels[4].label[145] , 
	\labels[4].label[144] , \labels[4].label[143] , 
	\labels[4].label[142] , \labels[4].label[141] , 
	\labels[4].label[140] , \labels[4].label[139] , 
	\labels[4].label[138] , \labels[4].label[137] , 
	\labels[4].label[136] , \labels[4].label[135] , 
	\labels[4].label[134] , \labels[4].label[133] , 
	\labels[4].label[132] , \labels[4].label[131] , 
	\labels[4].label[130] , \labels[4].label[129] , 
	\labels[4].label[128] , \labels[4].label[127] , 
	\labels[4].label[126] , \labels[4].label[125] , 
	\labels[4].label[124] , \labels[4].label[123] , 
	\labels[4].label[122] , \labels[4].label[121] , 
	\labels[4].label[120] , \labels[4].label[119] , 
	\labels[4].label[118] , \labels[4].label[117] , 
	\labels[4].label[116] , \labels[4].label[115] , 
	\labels[4].label[114] , \labels[4].label[113] , 
	\labels[4].label[112] , \labels[4].label[111] , 
	\labels[4].label[110] , \labels[4].label[109] , 
	\labels[4].label[108] , \labels[4].label[107] , 
	\labels[4].label[106] , \labels[4].label[105] , 
	\labels[4].label[104] , \labels[4].label[103] , 
	\labels[4].label[102] , \labels[4].label[101] , 
	\labels[4].label[100] , \labels[4].label[99] , \labels[4].label[98] , 
	\labels[4].label[97] , \labels[4].label[96] , \labels[4].label[95] , 
	\labels[4].label[94] , \labels[4].label[93] , \labels[4].label[92] , 
	\labels[4].label[91] , \labels[4].label[90] , \labels[4].label[89] , 
	\labels[4].label[88] , \labels[4].label[87] , \labels[4].label[86] , 
	\labels[4].label[85] , \labels[4].label[84] , \labels[4].label[83] , 
	\labels[4].label[82] , \labels[4].label[81] , \labels[4].label[80] , 
	\labels[4].label[79] , \labels[4].label[78] , \labels[4].label[77] , 
	\labels[4].label[76] , \labels[4].label[75] , \labels[4].label[74] , 
	\labels[4].label[73] , \labels[4].label[72] , \labels[4].label[71] , 
	\labels[4].label[70] , \labels[4].label[69] , \labels[4].label[68] , 
	\labels[4].label[67] , \labels[4].label[66] , \labels[4].label[65] , 
	\labels[4].label[64] , \labels[4].label[63] , \labels[4].label[62] , 
	\labels[4].label[61] , \labels[4].label[60] , \labels[4].label[59] , 
	\labels[4].label[58] , \labels[4].label[57] , \labels[4].label[56] , 
	\labels[4].label[55] , \labels[4].label[54] , \labels[4].label[53] , 
	\labels[4].label[52] , \labels[4].label[51] , \labels[4].label[50] , 
	\labels[4].label[49] , \labels[4].label[48] , \labels[4].label[47] , 
	\labels[4].label[46] , \labels[4].label[45] , \labels[4].label[44] , 
	\labels[4].label[43] , \labels[4].label[42] , \labels[4].label[41] , 
	\labels[4].label[40] , \labels[4].label[39] , \labels[4].label[38] , 
	\labels[4].label[37] , \labels[4].label[36] , \labels[4].label[35] , 
	\labels[4].label[34] , \labels[4].label[33] , \labels[4].label[32] , 
	\labels[4].label[31] , \labels[4].label[30] , \labels[4].label[29] , 
	\labels[4].label[28] , \labels[4].label[27] , \labels[4].label[26] , 
	\labels[4].label[25] , \labels[4].label[24] , \labels[4].label[23] , 
	\labels[4].label[22] , \labels[4].label[21] , \labels[4].label[20] , 
	\labels[4].label[19] , \labels[4].label[18] , \labels[4].label[17] , 
	\labels[4].label[16] , \labels[4].label[15] , \labels[4].label[14] , 
	\labels[4].label[13] , \labels[4].label[12] , \labels[4].label[11] , 
	\labels[4].label[10] , \labels[4].label[9] , \labels[4].label[8] , 
	\labels[4].label[7] , \labels[4].label[6] , \labels[4].label[5] , 
	\labels[4].label[4] , \labels[4].label[3] , \labels[4].label[2] , 
	\labels[4].label[1] , \labels[4].label[0] , 
	\labels[4].delimiter_valid[0] , \labels[4].delimiter[7] , 
	\labels[4].delimiter[6] , \labels[4].delimiter[5] , 
	\labels[4].delimiter[4] , \labels[4].delimiter[3] , 
	\labels[4].delimiter[2] , \labels[4].delimiter[1] , 
	\labels[4].delimiter[0] , \labels[3].guid_size[0] , 
	\labels[3].label_size[5] , \labels[3].label_size[4] , 
	\labels[3].label_size[3] , \labels[3].label_size[2] , 
	\labels[3].label_size[1] , \labels[3].label_size[0] , 
	\labels[3].label[255] , \labels[3].label[254] , 
	\labels[3].label[253] , \labels[3].label[252] , 
	\labels[3].label[251] , \labels[3].label[250] , 
	\labels[3].label[249] , \labels[3].label[248] , 
	\labels[3].label[247] , \labels[3].label[246] , 
	\labels[3].label[245] , \labels[3].label[244] , 
	\labels[3].label[243] , \labels[3].label[242] , 
	\labels[3].label[241] , \labels[3].label[240] , 
	\labels[3].label[239] , \labels[3].label[238] , 
	\labels[3].label[237] , \labels[3].label[236] , 
	\labels[3].label[235] , \labels[3].label[234] , 
	\labels[3].label[233] , \labels[3].label[232] , 
	\labels[3].label[231] , \labels[3].label[230] , 
	\labels[3].label[229] , \labels[3].label[228] , 
	\labels[3].label[227] , \labels[3].label[226] , 
	\labels[3].label[225] , \labels[3].label[224] , 
	\labels[3].label[223] , \labels[3].label[222] , 
	\labels[3].label[221] , \labels[3].label[220] , 
	\labels[3].label[219] , \labels[3].label[218] , 
	\labels[3].label[217] , \labels[3].label[216] , 
	\labels[3].label[215] , \labels[3].label[214] , 
	\labels[3].label[213] , \labels[3].label[212] , 
	\labels[3].label[211] , \labels[3].label[210] , 
	\labels[3].label[209] , \labels[3].label[208] , 
	\labels[3].label[207] , \labels[3].label[206] , 
	\labels[3].label[205] , \labels[3].label[204] , 
	\labels[3].label[203] , \labels[3].label[202] , 
	\labels[3].label[201] , \labels[3].label[200] , 
	\labels[3].label[199] , \labels[3].label[198] , 
	\labels[3].label[197] , \labels[3].label[196] , 
	\labels[3].label[195] , \labels[3].label[194] , 
	\labels[3].label[193] , \labels[3].label[192] , 
	\labels[3].label[191] , \labels[3].label[190] , 
	\labels[3].label[189] , \labels[3].label[188] , 
	\labels[3].label[187] , \labels[3].label[186] , 
	\labels[3].label[185] , \labels[3].label[184] , 
	\labels[3].label[183] , \labels[3].label[182] , 
	\labels[3].label[181] , \labels[3].label[180] , 
	\labels[3].label[179] , \labels[3].label[178] , 
	\labels[3].label[177] , \labels[3].label[176] , 
	\labels[3].label[175] , \labels[3].label[174] , 
	\labels[3].label[173] , \labels[3].label[172] , 
	\labels[3].label[171] , \labels[3].label[170] , 
	\labels[3].label[169] , \labels[3].label[168] , 
	\labels[3].label[167] , \labels[3].label[166] , 
	\labels[3].label[165] , \labels[3].label[164] , 
	\labels[3].label[163] , \labels[3].label[162] , 
	\labels[3].label[161] , \labels[3].label[160] , 
	\labels[3].label[159] , \labels[3].label[158] , 
	\labels[3].label[157] , \labels[3].label[156] , 
	\labels[3].label[155] , \labels[3].label[154] , 
	\labels[3].label[153] , \labels[3].label[152] , 
	\labels[3].label[151] , \labels[3].label[150] , 
	\labels[3].label[149] , \labels[3].label[148] , 
	\labels[3].label[147] , \labels[3].label[146] , 
	\labels[3].label[145] , \labels[3].label[144] , 
	\labels[3].label[143] , \labels[3].label[142] , 
	\labels[3].label[141] , \labels[3].label[140] , 
	\labels[3].label[139] , \labels[3].label[138] , 
	\labels[3].label[137] , \labels[3].label[136] , 
	\labels[3].label[135] , \labels[3].label[134] , 
	\labels[3].label[133] , \labels[3].label[132] , 
	\labels[3].label[131] , \labels[3].label[130] , 
	\labels[3].label[129] , \labels[3].label[128] , 
	\labels[3].label[127] , \labels[3].label[126] , 
	\labels[3].label[125] , \labels[3].label[124] , 
	\labels[3].label[123] , \labels[3].label[122] , 
	\labels[3].label[121] , \labels[3].label[120] , 
	\labels[3].label[119] , \labels[3].label[118] , 
	\labels[3].label[117] , \labels[3].label[116] , 
	\labels[3].label[115] , \labels[3].label[114] , 
	\labels[3].label[113] , \labels[3].label[112] , 
	\labels[3].label[111] , \labels[3].label[110] , 
	\labels[3].label[109] , \labels[3].label[108] , 
	\labels[3].label[107] , \labels[3].label[106] , 
	\labels[3].label[105] , \labels[3].label[104] , 
	\labels[3].label[103] , \labels[3].label[102] , 
	\labels[3].label[101] , \labels[3].label[100] , 
	\labels[3].label[99] , \labels[3].label[98] , \labels[3].label[97] , 
	\labels[3].label[96] , \labels[3].label[95] , \labels[3].label[94] , 
	\labels[3].label[93] , \labels[3].label[92] , \labels[3].label[91] , 
	\labels[3].label[90] , \labels[3].label[89] , \labels[3].label[88] , 
	\labels[3].label[87] , \labels[3].label[86] , \labels[3].label[85] , 
	\labels[3].label[84] , \labels[3].label[83] , \labels[3].label[82] , 
	\labels[3].label[81] , \labels[3].label[80] , \labels[3].label[79] , 
	\labels[3].label[78] , \labels[3].label[77] , \labels[3].label[76] , 
	\labels[3].label[75] , \labels[3].label[74] , \labels[3].label[73] , 
	\labels[3].label[72] , \labels[3].label[71] , \labels[3].label[70] , 
	\labels[3].label[69] , \labels[3].label[68] , \labels[3].label[67] , 
	\labels[3].label[66] , \labels[3].label[65] , \labels[3].label[64] , 
	\labels[3].label[63] , \labels[3].label[62] , \labels[3].label[61] , 
	\labels[3].label[60] , \labels[3].label[59] , \labels[3].label[58] , 
	\labels[3].label[57] , \labels[3].label[56] , \labels[3].label[55] , 
	\labels[3].label[54] , \labels[3].label[53] , \labels[3].label[52] , 
	\labels[3].label[51] , \labels[3].label[50] , \labels[3].label[49] , 
	\labels[3].label[48] , \labels[3].label[47] , \labels[3].label[46] , 
	\labels[3].label[45] , \labels[3].label[44] , \labels[3].label[43] , 
	\labels[3].label[42] , \labels[3].label[41] , \labels[3].label[40] , 
	\labels[3].label[39] , \labels[3].label[38] , \labels[3].label[37] , 
	\labels[3].label[36] , \labels[3].label[35] , \labels[3].label[34] , 
	\labels[3].label[33] , \labels[3].label[32] , \labels[3].label[31] , 
	\labels[3].label[30] , \labels[3].label[29] , \labels[3].label[28] , 
	\labels[3].label[27] , \labels[3].label[26] , \labels[3].label[25] , 
	\labels[3].label[24] , \labels[3].label[23] , \labels[3].label[22] , 
	\labels[3].label[21] , \labels[3].label[20] , \labels[3].label[19] , 
	\labels[3].label[18] , \labels[3].label[17] , \labels[3].label[16] , 
	\labels[3].label[15] , \labels[3].label[14] , \labels[3].label[13] , 
	\labels[3].label[12] , \labels[3].label[11] , \labels[3].label[10] , 
	\labels[3].label[9] , \labels[3].label[8] , \labels[3].label[7] , 
	\labels[3].label[6] , \labels[3].label[5] , \labels[3].label[4] , 
	\labels[3].label[3] , \labels[3].label[2] , \labels[3].label[1] , 
	\labels[3].label[0] , \labels[3].delimiter_valid[0] , 
	\labels[3].delimiter[7] , \labels[3].delimiter[6] , 
	\labels[3].delimiter[5] , \labels[3].delimiter[4] , 
	\labels[3].delimiter[3] , \labels[3].delimiter[2] , 
	\labels[3].delimiter[1] , \labels[3].delimiter[0] , 
	\labels[2].guid_size[0] , \labels[2].label_size[5] , 
	\labels[2].label_size[4] , \labels[2].label_size[3] , 
	\labels[2].label_size[2] , \labels[2].label_size[1] , 
	\labels[2].label_size[0] , \labels[2].label[255] , 
	\labels[2].label[254] , \labels[2].label[253] , 
	\labels[2].label[252] , \labels[2].label[251] , 
	\labels[2].label[250] , \labels[2].label[249] , 
	\labels[2].label[248] , \labels[2].label[247] , 
	\labels[2].label[246] , \labels[2].label[245] , 
	\labels[2].label[244] , \labels[2].label[243] , 
	\labels[2].label[242] , \labels[2].label[241] , 
	\labels[2].label[240] , \labels[2].label[239] , 
	\labels[2].label[238] , \labels[2].label[237] , 
	\labels[2].label[236] , \labels[2].label[235] , 
	\labels[2].label[234] , \labels[2].label[233] , 
	\labels[2].label[232] , \labels[2].label[231] , 
	\labels[2].label[230] , \labels[2].label[229] , 
	\labels[2].label[228] , \labels[2].label[227] , 
	\labels[2].label[226] , \labels[2].label[225] , 
	\labels[2].label[224] , \labels[2].label[223] , 
	\labels[2].label[222] , \labels[2].label[221] , 
	\labels[2].label[220] , \labels[2].label[219] , 
	\labels[2].label[218] , \labels[2].label[217] , 
	\labels[2].label[216] , \labels[2].label[215] , 
	\labels[2].label[214] , \labels[2].label[213] , 
	\labels[2].label[212] , \labels[2].label[211] , 
	\labels[2].label[210] , \labels[2].label[209] , 
	\labels[2].label[208] , \labels[2].label[207] , 
	\labels[2].label[206] , \labels[2].label[205] , 
	\labels[2].label[204] , \labels[2].label[203] , 
	\labels[2].label[202] , \labels[2].label[201] , 
	\labels[2].label[200] , \labels[2].label[199] , 
	\labels[2].label[198] , \labels[2].label[197] , 
	\labels[2].label[196] , \labels[2].label[195] , 
	\labels[2].label[194] , \labels[2].label[193] , 
	\labels[2].label[192] , \labels[2].label[191] , 
	\labels[2].label[190] , \labels[2].label[189] , 
	\labels[2].label[188] , \labels[2].label[187] , 
	\labels[2].label[186] , \labels[2].label[185] , 
	\labels[2].label[184] , \labels[2].label[183] , 
	\labels[2].label[182] , \labels[2].label[181] , 
	\labels[2].label[180] , \labels[2].label[179] , 
	\labels[2].label[178] , \labels[2].label[177] , 
	\labels[2].label[176] , \labels[2].label[175] , 
	\labels[2].label[174] , \labels[2].label[173] , 
	\labels[2].label[172] , \labels[2].label[171] , 
	\labels[2].label[170] , \labels[2].label[169] , 
	\labels[2].label[168] , \labels[2].label[167] , 
	\labels[2].label[166] , \labels[2].label[165] , 
	\labels[2].label[164] , \labels[2].label[163] , 
	\labels[2].label[162] , \labels[2].label[161] , 
	\labels[2].label[160] , \labels[2].label[159] , 
	\labels[2].label[158] , \labels[2].label[157] , 
	\labels[2].label[156] , \labels[2].label[155] , 
	\labels[2].label[154] , \labels[2].label[153] , 
	\labels[2].label[152] , \labels[2].label[151] , 
	\labels[2].label[150] , \labels[2].label[149] , 
	\labels[2].label[148] , \labels[2].label[147] , 
	\labels[2].label[146] , \labels[2].label[145] , 
	\labels[2].label[144] , \labels[2].label[143] , 
	\labels[2].label[142] , \labels[2].label[141] , 
	\labels[2].label[140] , \labels[2].label[139] , 
	\labels[2].label[138] , \labels[2].label[137] , 
	\labels[2].label[136] , \labels[2].label[135] , 
	\labels[2].label[134] , \labels[2].label[133] , 
	\labels[2].label[132] , \labels[2].label[131] , 
	\labels[2].label[130] , \labels[2].label[129] , 
	\labels[2].label[128] , \labels[2].label[127] , 
	\labels[2].label[126] , \labels[2].label[125] , 
	\labels[2].label[124] , \labels[2].label[123] , 
	\labels[2].label[122] , \labels[2].label[121] , 
	\labels[2].label[120] , \labels[2].label[119] , 
	\labels[2].label[118] , \labels[2].label[117] , 
	\labels[2].label[116] , \labels[2].label[115] , 
	\labels[2].label[114] , \labels[2].label[113] , 
	\labels[2].label[112] , \labels[2].label[111] , 
	\labels[2].label[110] , \labels[2].label[109] , 
	\labels[2].label[108] , \labels[2].label[107] , 
	\labels[2].label[106] , \labels[2].label[105] , 
	\labels[2].label[104] , \labels[2].label[103] , 
	\labels[2].label[102] , \labels[2].label[101] , 
	\labels[2].label[100] , \labels[2].label[99] , \labels[2].label[98] , 
	\labels[2].label[97] , \labels[2].label[96] , \labels[2].label[95] , 
	\labels[2].label[94] , \labels[2].label[93] , \labels[2].label[92] , 
	\labels[2].label[91] , \labels[2].label[90] , \labels[2].label[89] , 
	\labels[2].label[88] , \labels[2].label[87] , \labels[2].label[86] , 
	\labels[2].label[85] , \labels[2].label[84] , \labels[2].label[83] , 
	\labels[2].label[82] , \labels[2].label[81] , \labels[2].label[80] , 
	\labels[2].label[79] , \labels[2].label[78] , \labels[2].label[77] , 
	\labels[2].label[76] , \labels[2].label[75] , \labels[2].label[74] , 
	\labels[2].label[73] , \labels[2].label[72] , \labels[2].label[71] , 
	\labels[2].label[70] , \labels[2].label[69] , \labels[2].label[68] , 
	\labels[2].label[67] , \labels[2].label[66] , \labels[2].label[65] , 
	\labels[2].label[64] , \labels[2].label[63] , \labels[2].label[62] , 
	\labels[2].label[61] , \labels[2].label[60] , \labels[2].label[59] , 
	\labels[2].label[58] , \labels[2].label[57] , \labels[2].label[56] , 
	\labels[2].label[55] , \labels[2].label[54] , \labels[2].label[53] , 
	\labels[2].label[52] , \labels[2].label[51] , \labels[2].label[50] , 
	\labels[2].label[49] , \labels[2].label[48] , \labels[2].label[47] , 
	\labels[2].label[46] , \labels[2].label[45] , \labels[2].label[44] , 
	\labels[2].label[43] , \labels[2].label[42] , \labels[2].label[41] , 
	\labels[2].label[40] , \labels[2].label[39] , \labels[2].label[38] , 
	\labels[2].label[37] , \labels[2].label[36] , \labels[2].label[35] , 
	\labels[2].label[34] , \labels[2].label[33] , \labels[2].label[32] , 
	\labels[2].label[31] , \labels[2].label[30] , \labels[2].label[29] , 
	\labels[2].label[28] , \labels[2].label[27] , \labels[2].label[26] , 
	\labels[2].label[25] , \labels[2].label[24] , \labels[2].label[23] , 
	\labels[2].label[22] , \labels[2].label[21] , \labels[2].label[20] , 
	\labels[2].label[19] , \labels[2].label[18] , \labels[2].label[17] , 
	\labels[2].label[16] , \labels[2].label[15] , \labels[2].label[14] , 
	\labels[2].label[13] , \labels[2].label[12] , \labels[2].label[11] , 
	\labels[2].label[10] , \labels[2].label[9] , \labels[2].label[8] , 
	\labels[2].label[7] , \labels[2].label[6] , \labels[2].label[5] , 
	\labels[2].label[4] , \labels[2].label[3] , \labels[2].label[2] , 
	\labels[2].label[1] , \labels[2].label[0] , 
	\labels[2].delimiter_valid[0] , \labels[2].delimiter[7] , 
	\labels[2].delimiter[6] , \labels[2].delimiter[5] , 
	\labels[2].delimiter[4] , \labels[2].delimiter[3] , 
	\labels[2].delimiter[2] , \labels[2].delimiter[1] , 
	\labels[2].delimiter[0] , \labels[1].guid_size[0] , 
	\labels[1].label_size[5] , \labels[1].label_size[4] , 
	\labels[1].label_size[3] , \labels[1].label_size[2] , 
	\labels[1].label_size[1] , \labels[1].label_size[0] , 
	\labels[1].label[255] , \labels[1].label[254] , 
	\labels[1].label[253] , \labels[1].label[252] , 
	\labels[1].label[251] , \labels[1].label[250] , 
	\labels[1].label[249] , \labels[1].label[248] , 
	\labels[1].label[247] , \labels[1].label[246] , 
	\labels[1].label[245] , \labels[1].label[244] , 
	\labels[1].label[243] , \labels[1].label[242] , 
	\labels[1].label[241] , \labels[1].label[240] , 
	\labels[1].label[239] , \labels[1].label[238] , 
	\labels[1].label[237] , \labels[1].label[236] , 
	\labels[1].label[235] , \labels[1].label[234] , 
	\labels[1].label[233] , \labels[1].label[232] , 
	\labels[1].label[231] , \labels[1].label[230] , 
	\labels[1].label[229] , \labels[1].label[228] , 
	\labels[1].label[227] , \labels[1].label[226] , 
	\labels[1].label[225] , \labels[1].label[224] , 
	\labels[1].label[223] , \labels[1].label[222] , 
	\labels[1].label[221] , \labels[1].label[220] , 
	\labels[1].label[219] , \labels[1].label[218] , 
	\labels[1].label[217] , \labels[1].label[216] , 
	\labels[1].label[215] , \labels[1].label[214] , 
	\labels[1].label[213] , \labels[1].label[212] , 
	\labels[1].label[211] , \labels[1].label[210] , 
	\labels[1].label[209] , \labels[1].label[208] , 
	\labels[1].label[207] , \labels[1].label[206] , 
	\labels[1].label[205] , \labels[1].label[204] , 
	\labels[1].label[203] , \labels[1].label[202] , 
	\labels[1].label[201] , \labels[1].label[200] , 
	\labels[1].label[199] , \labels[1].label[198] , 
	\labels[1].label[197] , \labels[1].label[196] , 
	\labels[1].label[195] , \labels[1].label[194] , 
	\labels[1].label[193] , \labels[1].label[192] , 
	\labels[1].label[191] , \labels[1].label[190] , 
	\labels[1].label[189] , \labels[1].label[188] , 
	\labels[1].label[187] , \labels[1].label[186] , 
	\labels[1].label[185] , \labels[1].label[184] , 
	\labels[1].label[183] , \labels[1].label[182] , 
	\labels[1].label[181] , \labels[1].label[180] , 
	\labels[1].label[179] , \labels[1].label[178] , 
	\labels[1].label[177] , \labels[1].label[176] , 
	\labels[1].label[175] , \labels[1].label[174] , 
	\labels[1].label[173] , \labels[1].label[172] , 
	\labels[1].label[171] , \labels[1].label[170] , 
	\labels[1].label[169] , \labels[1].label[168] , 
	\labels[1].label[167] , \labels[1].label[166] , 
	\labels[1].label[165] , \labels[1].label[164] , 
	\labels[1].label[163] , \labels[1].label[162] , 
	\labels[1].label[161] , \labels[1].label[160] , 
	\labels[1].label[159] , \labels[1].label[158] , 
	\labels[1].label[157] , \labels[1].label[156] , 
	\labels[1].label[155] , \labels[1].label[154] , 
	\labels[1].label[153] , \labels[1].label[152] , 
	\labels[1].label[151] , \labels[1].label[150] , 
	\labels[1].label[149] , \labels[1].label[148] , 
	\labels[1].label[147] , \labels[1].label[146] , 
	\labels[1].label[145] , \labels[1].label[144] , 
	\labels[1].label[143] , \labels[1].label[142] , 
	\labels[1].label[141] , \labels[1].label[140] , 
	\labels[1].label[139] , \labels[1].label[138] , 
	\labels[1].label[137] , \labels[1].label[136] , 
	\labels[1].label[135] , \labels[1].label[134] , 
	\labels[1].label[133] , \labels[1].label[132] , 
	\labels[1].label[131] , \labels[1].label[130] , 
	\labels[1].label[129] , \labels[1].label[128] , 
	\labels[1].label[127] , \labels[1].label[126] , 
	\labels[1].label[125] , \labels[1].label[124] , 
	\labels[1].label[123] , \labels[1].label[122] , 
	\labels[1].label[121] , \labels[1].label[120] , 
	\labels[1].label[119] , \labels[1].label[118] , 
	\labels[1].label[117] , \labels[1].label[116] , 
	\labels[1].label[115] , \labels[1].label[114] , 
	\labels[1].label[113] , \labels[1].label[112] , 
	\labels[1].label[111] , \labels[1].label[110] , 
	\labels[1].label[109] , \labels[1].label[108] , 
	\labels[1].label[107] , \labels[1].label[106] , 
	\labels[1].label[105] , \labels[1].label[104] , 
	\labels[1].label[103] , \labels[1].label[102] , 
	\labels[1].label[101] , \labels[1].label[100] , 
	\labels[1].label[99] , \labels[1].label[98] , \labels[1].label[97] , 
	\labels[1].label[96] , \labels[1].label[95] , \labels[1].label[94] , 
	\labels[1].label[93] , \labels[1].label[92] , \labels[1].label[91] , 
	\labels[1].label[90] , \labels[1].label[89] , \labels[1].label[88] , 
	\labels[1].label[87] , \labels[1].label[86] , \labels[1].label[85] , 
	\labels[1].label[84] , \labels[1].label[83] , \labels[1].label[82] , 
	\labels[1].label[81] , \labels[1].label[80] , \labels[1].label[79] , 
	\labels[1].label[78] , \labels[1].label[77] , \labels[1].label[76] , 
	\labels[1].label[75] , \labels[1].label[74] , \labels[1].label[73] , 
	\labels[1].label[72] , \labels[1].label[71] , \labels[1].label[70] , 
	\labels[1].label[69] , \labels[1].label[68] , \labels[1].label[67] , 
	\labels[1].label[66] , \labels[1].label[65] , \labels[1].label[64] , 
	\labels[1].label[63] , \labels[1].label[62] , \labels[1].label[61] , 
	\labels[1].label[60] , \labels[1].label[59] , \labels[1].label[58] , 
	\labels[1].label[57] , \labels[1].label[56] , \labels[1].label[55] , 
	\labels[1].label[54] , \labels[1].label[53] , \labels[1].label[52] , 
	\labels[1].label[51] , \labels[1].label[50] , \labels[1].label[49] , 
	\labels[1].label[48] , \labels[1].label[47] , \labels[1].label[46] , 
	\labels[1].label[45] , \labels[1].label[44] , \labels[1].label[43] , 
	\labels[1].label[42] , \labels[1].label[41] , \labels[1].label[40] , 
	\labels[1].label[39] , \labels[1].label[38] , \labels[1].label[37] , 
	\labels[1].label[36] , \labels[1].label[35] , \labels[1].label[34] , 
	\labels[1].label[33] , \labels[1].label[32] , \labels[1].label[31] , 
	\labels[1].label[30] , \labels[1].label[29] , \labels[1].label[28] , 
	\labels[1].label[27] , \labels[1].label[26] , \labels[1].label[25] , 
	\labels[1].label[24] , \labels[1].label[23] , \labels[1].label[22] , 
	\labels[1].label[21] , \labels[1].label[20] , \labels[1].label[19] , 
	\labels[1].label[18] , \labels[1].label[17] , \labels[1].label[16] , 
	\labels[1].label[15] , \labels[1].label[14] , \labels[1].label[13] , 
	\labels[1].label[12] , \labels[1].label[11] , \labels[1].label[10] , 
	\labels[1].label[9] , \labels[1].label[8] , \labels[1].label[7] , 
	\labels[1].label[6] , \labels[1].label[5] , \labels[1].label[4] , 
	\labels[1].label[3] , \labels[1].label[2] , \labels[1].label[1] , 
	\labels[1].label[0] , \labels[1].delimiter_valid[0] , 
	\labels[1].delimiter[7] , \labels[1].delimiter[6] , 
	\labels[1].delimiter[5] , \labels[1].delimiter[4] , 
	\labels[1].delimiter[3] , \labels[1].delimiter[2] , 
	\labels[1].delimiter[1] , \labels[1].delimiter[0] , 
	\labels[0].guid_size[0] , \labels[0].label_size[5] , 
	\labels[0].label_size[4] , \labels[0].label_size[3] , 
	\labels[0].label_size[2] , \labels[0].label_size[1] , 
	\labels[0].label_size[0] , \labels[0].label[255] , 
	\labels[0].label[254] , \labels[0].label[253] , 
	\labels[0].label[252] , \labels[0].label[251] , 
	\labels[0].label[250] , \labels[0].label[249] , 
	\labels[0].label[248] , \labels[0].label[247] , 
	\labels[0].label[246] , \labels[0].label[245] , 
	\labels[0].label[244] , \labels[0].label[243] , 
	\labels[0].label[242] , \labels[0].label[241] , 
	\labels[0].label[240] , \labels[0].label[239] , 
	\labels[0].label[238] , \labels[0].label[237] , 
	\labels[0].label[236] , \labels[0].label[235] , 
	\labels[0].label[234] , \labels[0].label[233] , 
	\labels[0].label[232] , \labels[0].label[231] , 
	\labels[0].label[230] , \labels[0].label[229] , 
	\labels[0].label[228] , \labels[0].label[227] , 
	\labels[0].label[226] , \labels[0].label[225] , 
	\labels[0].label[224] , \labels[0].label[223] , 
	\labels[0].label[222] , \labels[0].label[221] , 
	\labels[0].label[220] , \labels[0].label[219] , 
	\labels[0].label[218] , \labels[0].label[217] , 
	\labels[0].label[216] , \labels[0].label[215] , 
	\labels[0].label[214] , \labels[0].label[213] , 
	\labels[0].label[212] , \labels[0].label[211] , 
	\labels[0].label[210] , \labels[0].label[209] , 
	\labels[0].label[208] , \labels[0].label[207] , 
	\labels[0].label[206] , \labels[0].label[205] , 
	\labels[0].label[204] , \labels[0].label[203] , 
	\labels[0].label[202] , \labels[0].label[201] , 
	\labels[0].label[200] , \labels[0].label[199] , 
	\labels[0].label[198] , \labels[0].label[197] , 
	\labels[0].label[196] , \labels[0].label[195] , 
	\labels[0].label[194] , \labels[0].label[193] , 
	\labels[0].label[192] , \labels[0].label[191] , 
	\labels[0].label[190] , \labels[0].label[189] , 
	\labels[0].label[188] , \labels[0].label[187] , 
	\labels[0].label[186] , \labels[0].label[185] , 
	\labels[0].label[184] , \labels[0].label[183] , 
	\labels[0].label[182] , \labels[0].label[181] , 
	\labels[0].label[180] , \labels[0].label[179] , 
	\labels[0].label[178] , \labels[0].label[177] , 
	\labels[0].label[176] , \labels[0].label[175] , 
	\labels[0].label[174] , \labels[0].label[173] , 
	\labels[0].label[172] , \labels[0].label[171] , 
	\labels[0].label[170] , \labels[0].label[169] , 
	\labels[0].label[168] , \labels[0].label[167] , 
	\labels[0].label[166] , \labels[0].label[165] , 
	\labels[0].label[164] , \labels[0].label[163] , 
	\labels[0].label[162] , \labels[0].label[161] , 
	\labels[0].label[160] , \labels[0].label[159] , 
	\labels[0].label[158] , \labels[0].label[157] , 
	\labels[0].label[156] , \labels[0].label[155] , 
	\labels[0].label[154] , \labels[0].label[153] , 
	\labels[0].label[152] , \labels[0].label[151] , 
	\labels[0].label[150] , \labels[0].label[149] , 
	\labels[0].label[148] , \labels[0].label[147] , 
	\labels[0].label[146] , \labels[0].label[145] , 
	\labels[0].label[144] , \labels[0].label[143] , 
	\labels[0].label[142] , \labels[0].label[141] , 
	\labels[0].label[140] , \labels[0].label[139] , 
	\labels[0].label[138] , \labels[0].label[137] , 
	\labels[0].label[136] , \labels[0].label[135] , 
	\labels[0].label[134] , \labels[0].label[133] , 
	\labels[0].label[132] , \labels[0].label[131] , 
	\labels[0].label[130] , \labels[0].label[129] , 
	\labels[0].label[128] , \labels[0].label[127] , 
	\labels[0].label[126] , \labels[0].label[125] , 
	\labels[0].label[124] , \labels[0].label[123] , 
	\labels[0].label[122] , \labels[0].label[121] , 
	\labels[0].label[120] , \labels[0].label[119] , 
	\labels[0].label[118] , \labels[0].label[117] , 
	\labels[0].label[116] , \labels[0].label[115] , 
	\labels[0].label[114] , \labels[0].label[113] , 
	\labels[0].label[112] , \labels[0].label[111] , 
	\labels[0].label[110] , \labels[0].label[109] , 
	\labels[0].label[108] , \labels[0].label[107] , 
	\labels[0].label[106] , \labels[0].label[105] , 
	\labels[0].label[104] , \labels[0].label[103] , 
	\labels[0].label[102] , \labels[0].label[101] , 
	\labels[0].label[100] , \labels[0].label[99] , \labels[0].label[98] , 
	\labels[0].label[97] , \labels[0].label[96] , \labels[0].label[95] , 
	\labels[0].label[94] , \labels[0].label[93] , \labels[0].label[92] , 
	\labels[0].label[91] , \labels[0].label[90] , \labels[0].label[89] , 
	\labels[0].label[88] , \labels[0].label[87] , \labels[0].label[86] , 
	\labels[0].label[85] , \labels[0].label[84] , \labels[0].label[83] , 
	\labels[0].label[82] , \labels[0].label[81] , \labels[0].label[80] , 
	\labels[0].label[79] , \labels[0].label[78] , \labels[0].label[77] , 
	\labels[0].label[76] , \labels[0].label[75] , \labels[0].label[74] , 
	\labels[0].label[73] , \labels[0].label[72] , \labels[0].label[71] , 
	\labels[0].label[70] , \labels[0].label[69] , \labels[0].label[68] , 
	\labels[0].label[67] , \labels[0].label[66] , \labels[0].label[65] , 
	\labels[0].label[64] , \labels[0].label[63] , \labels[0].label[62] , 
	\labels[0].label[61] , \labels[0].label[60] , \labels[0].label[59] , 
	\labels[0].label[58] , \labels[0].label[57] , \labels[0].label[56] , 
	\labels[0].label[55] , \labels[0].label[54] , \labels[0].label[53] , 
	\labels[0].label[52] , \labels[0].label[51] , \labels[0].label[50] , 
	\labels[0].label[49] , \labels[0].label[48] , \labels[0].label[47] , 
	\labels[0].label[46] , \labels[0].label[45] , \labels[0].label[44] , 
	\labels[0].label[43] , \labels[0].label[42] , \labels[0].label[41] , 
	\labels[0].label[40] , \labels[0].label[39] , \labels[0].label[38] , 
	\labels[0].label[37] , \labels[0].label[36] , \labels[0].label[35] , 
	\labels[0].label[34] , \labels[0].label[33] , \labels[0].label[32] , 
	\labels[0].label[31] , \labels[0].label[30] , \labels[0].label[29] , 
	\labels[0].label[28] , \labels[0].label[27] , \labels[0].label[26] , 
	\labels[0].label[25] , \labels[0].label[24] , \labels[0].label[23] , 
	\labels[0].label[22] , \labels[0].label[21] , \labels[0].label[20] , 
	\labels[0].label[19] , \labels[0].label[18] , \labels[0].label[17] , 
	\labels[0].label[16] , \labels[0].label[15] , \labels[0].label[14] , 
	\labels[0].label[13] , \labels[0].label[12] , \labels[0].label[11] , 
	\labels[0].label[10] , \labels[0].label[9] , \labels[0].label[8] , 
	\labels[0].label[7] , \labels[0].label[6] , \labels[0].label[5] , 
	\labels[0].label[4] , \labels[0].label[3] , \labels[0].label[2] , 
	\labels[0].label[1] , \labels[0].label[0] , 
	\labels[0].delimiter_valid[0] , \labels[0].delimiter[7] , 
	\labels[0].delimiter[6] , \labels[0].delimiter[5] , 
	\labels[0].delimiter[4] , \labels[0].delimiter[3] , 
	\labels[0].delimiter[2] , \labels[0].delimiter[1] , 
	\labels[0].delimiter[0] } ), seed0_valid, seed0_internal_state_key, 
	seed0_internal_state_value, seed0_reseed_interval, seed1_valid, 
	seed1_internal_state_key, seed1_internal_state_value, 
	seed1_reseed_interval, .tready_override( {
	\tready_override.r.part0 [8], \tready_override.r.part0 [7], 
	\tready_override.r.part0 [6], \tready_override.r.part0 [5], 
	\tready_override.r.part0 [4], \tready_override.r.part0 [3], 
	\tready_override.r.part0 [2], \tready_override.r.part0 [1], 
	\tready_override.r.part0 [0]} ), .cceip_encrypt_kop_fifo_override( {
	\cceip_encrypt_kop_fifo_override.r.part0 [6], 
	\cceip_encrypt_kop_fifo_override.r.part0 [5], 
	\cceip_encrypt_kop_fifo_override.r.part0 [4], 
	\cceip_encrypt_kop_fifo_override.r.part0 [3], 
	\cceip_encrypt_kop_fifo_override.r.part0 [2], 
	\cceip_encrypt_kop_fifo_override.r.part0 [1], 
	\cceip_encrypt_kop_fifo_override.r.part0 [0]} ), 
	.cceip_validate_kop_fifo_override( {
	\cceip_validate_kop_fifo_override.r.part0 [6], 
	\cceip_validate_kop_fifo_override.r.part0 [5], 
	\cceip_validate_kop_fifo_override.r.part0 [4], 
	\cceip_validate_kop_fifo_override.r.part0 [3], 
	\cceip_validate_kop_fifo_override.r.part0 [2], 
	\cceip_validate_kop_fifo_override.r.part0 [1], 
	\cceip_validate_kop_fifo_override.r.part0 [0]} ), 
	.cddip_decrypt_kop_fifo_override( {
	\cddip_decrypt_kop_fifo_override.r.part0 [6], 
	\cddip_decrypt_kop_fifo_override.r.part0 [5], 
	\cddip_decrypt_kop_fifo_override.r.part0 [4], 
	\cddip_decrypt_kop_fifo_override.r.part0 [3], 
	\cddip_decrypt_kop_fifo_override.r.part0 [2], 
	\cddip_decrypt_kop_fifo_override.r.part0 [1], 
	\cddip_decrypt_kop_fifo_override.r.part0 [0]} ), manual_txc, 
	always_validate_kim_ref, kdf_test_mode_en, kdf_test_key_size, 
	.sa_global_ctrl( {\sa_global_ctrl.r.part0 [31], 
	\sa_global_ctrl.r.part0 [30], \sa_global_ctrl.r.part0 [29], 
	\sa_global_ctrl.r.part0 [28], \sa_global_ctrl.r.part0 [27], 
	\sa_global_ctrl.r.part0 [26], \sa_global_ctrl.r.part0 [25], 
	\sa_global_ctrl.r.part0 [24], \sa_global_ctrl.r.part0 [23], 
	\sa_global_ctrl.r.part0 [22], \sa_global_ctrl.r.part0 [21], 
	\sa_global_ctrl.r.part0 [20], \sa_global_ctrl.r.part0 [19], 
	\sa_global_ctrl.r.part0 [18], \sa_global_ctrl.r.part0 [17], 
	\sa_global_ctrl.r.part0 [16], \sa_global_ctrl.r.part0 [15], 
	\sa_global_ctrl.r.part0 [14], \sa_global_ctrl.r.part0 [13], 
	\sa_global_ctrl.r.part0 [12], \sa_global_ctrl.r.part0 [11], 
	\sa_global_ctrl.r.part0 [10], \sa_global_ctrl.r.part0 [9], 
	\sa_global_ctrl.r.part0 [8], \sa_global_ctrl.r.part0 [7], 
	\sa_global_ctrl.r.part0 [6], \sa_global_ctrl.r.part0 [5], 
	\sa_global_ctrl.r.part0 [4], \sa_global_ctrl.r.part0 [3], 
	\sa_global_ctrl.r.part0 [2], \sa_global_ctrl.r.part0 [1], 
	\sa_global_ctrl.r.part0 [0]} ), .sa_ctrl( {
	\sa_ctrl[31].r.part0[31] , \sa_ctrl[31].r.part0[30] , 
	\sa_ctrl[31].r.part0[29] , \sa_ctrl[31].r.part0[28] , 
	\sa_ctrl[31].r.part0[27] , \sa_ctrl[31].r.part0[26] , 
	\sa_ctrl[31].r.part0[25] , \sa_ctrl[31].r.part0[24] , 
	\sa_ctrl[31].r.part0[23] , \sa_ctrl[31].r.part0[22] , 
	\sa_ctrl[31].r.part0[21] , \sa_ctrl[31].r.part0[20] , 
	\sa_ctrl[31].r.part0[19] , \sa_ctrl[31].r.part0[18] , 
	\sa_ctrl[31].r.part0[17] , \sa_ctrl[31].r.part0[16] , 
	\sa_ctrl[31].r.part0[15] , \sa_ctrl[31].r.part0[14] , 
	\sa_ctrl[31].r.part0[13] , \sa_ctrl[31].r.part0[12] , 
	\sa_ctrl[31].r.part0[11] , \sa_ctrl[31].r.part0[10] , 
	\sa_ctrl[31].r.part0[9] , \sa_ctrl[31].r.part0[8] , 
	\sa_ctrl[31].r.part0[7] , \sa_ctrl[31].r.part0[6] , 
	\sa_ctrl[31].r.part0[5] , \sa_ctrl[31].r.part0[4] , 
	\sa_ctrl[31].r.part0[3] , \sa_ctrl[31].r.part0[2] , 
	\sa_ctrl[31].r.part0[1] , \sa_ctrl[31].r.part0[0] , 
	\sa_ctrl[30].r.part0[31] , \sa_ctrl[30].r.part0[30] , 
	\sa_ctrl[30].r.part0[29] , \sa_ctrl[30].r.part0[28] , 
	\sa_ctrl[30].r.part0[27] , \sa_ctrl[30].r.part0[26] , 
	\sa_ctrl[30].r.part0[25] , \sa_ctrl[30].r.part0[24] , 
	\sa_ctrl[30].r.part0[23] , \sa_ctrl[30].r.part0[22] , 
	\sa_ctrl[30].r.part0[21] , \sa_ctrl[30].r.part0[20] , 
	\sa_ctrl[30].r.part0[19] , \sa_ctrl[30].r.part0[18] , 
	\sa_ctrl[30].r.part0[17] , \sa_ctrl[30].r.part0[16] , 
	\sa_ctrl[30].r.part0[15] , \sa_ctrl[30].r.part0[14] , 
	\sa_ctrl[30].r.part0[13] , \sa_ctrl[30].r.part0[12] , 
	\sa_ctrl[30].r.part0[11] , \sa_ctrl[30].r.part0[10] , 
	\sa_ctrl[30].r.part0[9] , \sa_ctrl[30].r.part0[8] , 
	\sa_ctrl[30].r.part0[7] , \sa_ctrl[30].r.part0[6] , 
	\sa_ctrl[30].r.part0[5] , \sa_ctrl[30].r.part0[4] , 
	\sa_ctrl[30].r.part0[3] , \sa_ctrl[30].r.part0[2] , 
	\sa_ctrl[30].r.part0[1] , \sa_ctrl[30].r.part0[0] , 
	\sa_ctrl[29].r.part0[31] , \sa_ctrl[29].r.part0[30] , 
	\sa_ctrl[29].r.part0[29] , \sa_ctrl[29].r.part0[28] , 
	\sa_ctrl[29].r.part0[27] , \sa_ctrl[29].r.part0[26] , 
	\sa_ctrl[29].r.part0[25] , \sa_ctrl[29].r.part0[24] , 
	\sa_ctrl[29].r.part0[23] , \sa_ctrl[29].r.part0[22] , 
	\sa_ctrl[29].r.part0[21] , \sa_ctrl[29].r.part0[20] , 
	\sa_ctrl[29].r.part0[19] , \sa_ctrl[29].r.part0[18] , 
	\sa_ctrl[29].r.part0[17] , \sa_ctrl[29].r.part0[16] , 
	\sa_ctrl[29].r.part0[15] , \sa_ctrl[29].r.part0[14] , 
	\sa_ctrl[29].r.part0[13] , \sa_ctrl[29].r.part0[12] , 
	\sa_ctrl[29].r.part0[11] , \sa_ctrl[29].r.part0[10] , 
	\sa_ctrl[29].r.part0[9] , \sa_ctrl[29].r.part0[8] , 
	\sa_ctrl[29].r.part0[7] , \sa_ctrl[29].r.part0[6] , 
	\sa_ctrl[29].r.part0[5] , \sa_ctrl[29].r.part0[4] , 
	\sa_ctrl[29].r.part0[3] , \sa_ctrl[29].r.part0[2] , 
	\sa_ctrl[29].r.part0[1] , \sa_ctrl[29].r.part0[0] , 
	\sa_ctrl[28].r.part0[31] , \sa_ctrl[28].r.part0[30] , 
	\sa_ctrl[28].r.part0[29] , \sa_ctrl[28].r.part0[28] , 
	\sa_ctrl[28].r.part0[27] , \sa_ctrl[28].r.part0[26] , 
	\sa_ctrl[28].r.part0[25] , \sa_ctrl[28].r.part0[24] , 
	\sa_ctrl[28].r.part0[23] , \sa_ctrl[28].r.part0[22] , 
	\sa_ctrl[28].r.part0[21] , \sa_ctrl[28].r.part0[20] , 
	\sa_ctrl[28].r.part0[19] , \sa_ctrl[28].r.part0[18] , 
	\sa_ctrl[28].r.part0[17] , \sa_ctrl[28].r.part0[16] , 
	\sa_ctrl[28].r.part0[15] , \sa_ctrl[28].r.part0[14] , 
	\sa_ctrl[28].r.part0[13] , \sa_ctrl[28].r.part0[12] , 
	\sa_ctrl[28].r.part0[11] , \sa_ctrl[28].r.part0[10] , 
	\sa_ctrl[28].r.part0[9] , \sa_ctrl[28].r.part0[8] , 
	\sa_ctrl[28].r.part0[7] , \sa_ctrl[28].r.part0[6] , 
	\sa_ctrl[28].r.part0[5] , \sa_ctrl[28].r.part0[4] , 
	\sa_ctrl[28].r.part0[3] , \sa_ctrl[28].r.part0[2] , 
	\sa_ctrl[28].r.part0[1] , \sa_ctrl[28].r.part0[0] , 
	\sa_ctrl[27].r.part0[31] , \sa_ctrl[27].r.part0[30] , 
	\sa_ctrl[27].r.part0[29] , \sa_ctrl[27].r.part0[28] , 
	\sa_ctrl[27].r.part0[27] , \sa_ctrl[27].r.part0[26] , 
	\sa_ctrl[27].r.part0[25] , \sa_ctrl[27].r.part0[24] , 
	\sa_ctrl[27].r.part0[23] , \sa_ctrl[27].r.part0[22] , 
	\sa_ctrl[27].r.part0[21] , \sa_ctrl[27].r.part0[20] , 
	\sa_ctrl[27].r.part0[19] , \sa_ctrl[27].r.part0[18] , 
	\sa_ctrl[27].r.part0[17] , \sa_ctrl[27].r.part0[16] , 
	\sa_ctrl[27].r.part0[15] , \sa_ctrl[27].r.part0[14] , 
	\sa_ctrl[27].r.part0[13] , \sa_ctrl[27].r.part0[12] , 
	\sa_ctrl[27].r.part0[11] , \sa_ctrl[27].r.part0[10] , 
	\sa_ctrl[27].r.part0[9] , \sa_ctrl[27].r.part0[8] , 
	\sa_ctrl[27].r.part0[7] , \sa_ctrl[27].r.part0[6] , 
	\sa_ctrl[27].r.part0[5] , \sa_ctrl[27].r.part0[4] , 
	\sa_ctrl[27].r.part0[3] , \sa_ctrl[27].r.part0[2] , 
	\sa_ctrl[27].r.part0[1] , \sa_ctrl[27].r.part0[0] , 
	\sa_ctrl[26].r.part0[31] , \sa_ctrl[26].r.part0[30] , 
	\sa_ctrl[26].r.part0[29] , \sa_ctrl[26].r.part0[28] , 
	\sa_ctrl[26].r.part0[27] , \sa_ctrl[26].r.part0[26] , 
	\sa_ctrl[26].r.part0[25] , \sa_ctrl[26].r.part0[24] , 
	\sa_ctrl[26].r.part0[23] , \sa_ctrl[26].r.part0[22] , 
	\sa_ctrl[26].r.part0[21] , \sa_ctrl[26].r.part0[20] , 
	\sa_ctrl[26].r.part0[19] , \sa_ctrl[26].r.part0[18] , 
	\sa_ctrl[26].r.part0[17] , \sa_ctrl[26].r.part0[16] , 
	\sa_ctrl[26].r.part0[15] , \sa_ctrl[26].r.part0[14] , 
	\sa_ctrl[26].r.part0[13] , \sa_ctrl[26].r.part0[12] , 
	\sa_ctrl[26].r.part0[11] , \sa_ctrl[26].r.part0[10] , 
	\sa_ctrl[26].r.part0[9] , \sa_ctrl[26].r.part0[8] , 
	\sa_ctrl[26].r.part0[7] , \sa_ctrl[26].r.part0[6] , 
	\sa_ctrl[26].r.part0[5] , \sa_ctrl[26].r.part0[4] , 
	\sa_ctrl[26].r.part0[3] , \sa_ctrl[26].r.part0[2] , 
	\sa_ctrl[26].r.part0[1] , \sa_ctrl[26].r.part0[0] , 
	\sa_ctrl[25].r.part0[31] , \sa_ctrl[25].r.part0[30] , 
	\sa_ctrl[25].r.part0[29] , \sa_ctrl[25].r.part0[28] , 
	\sa_ctrl[25].r.part0[27] , \sa_ctrl[25].r.part0[26] , 
	\sa_ctrl[25].r.part0[25] , \sa_ctrl[25].r.part0[24] , 
	\sa_ctrl[25].r.part0[23] , \sa_ctrl[25].r.part0[22] , 
	\sa_ctrl[25].r.part0[21] , \sa_ctrl[25].r.part0[20] , 
	\sa_ctrl[25].r.part0[19] , \sa_ctrl[25].r.part0[18] , 
	\sa_ctrl[25].r.part0[17] , \sa_ctrl[25].r.part0[16] , 
	\sa_ctrl[25].r.part0[15] , \sa_ctrl[25].r.part0[14] , 
	\sa_ctrl[25].r.part0[13] , \sa_ctrl[25].r.part0[12] , 
	\sa_ctrl[25].r.part0[11] , \sa_ctrl[25].r.part0[10] , 
	\sa_ctrl[25].r.part0[9] , \sa_ctrl[25].r.part0[8] , 
	\sa_ctrl[25].r.part0[7] , \sa_ctrl[25].r.part0[6] , 
	\sa_ctrl[25].r.part0[5] , \sa_ctrl[25].r.part0[4] , 
	\sa_ctrl[25].r.part0[3] , \sa_ctrl[25].r.part0[2] , 
	\sa_ctrl[25].r.part0[1] , \sa_ctrl[25].r.part0[0] , 
	\sa_ctrl[24].r.part0[31] , \sa_ctrl[24].r.part0[30] , 
	\sa_ctrl[24].r.part0[29] , \sa_ctrl[24].r.part0[28] , 
	\sa_ctrl[24].r.part0[27] , \sa_ctrl[24].r.part0[26] , 
	\sa_ctrl[24].r.part0[25] , \sa_ctrl[24].r.part0[24] , 
	\sa_ctrl[24].r.part0[23] , \sa_ctrl[24].r.part0[22] , 
	\sa_ctrl[24].r.part0[21] , \sa_ctrl[24].r.part0[20] , 
	\sa_ctrl[24].r.part0[19] , \sa_ctrl[24].r.part0[18] , 
	\sa_ctrl[24].r.part0[17] , \sa_ctrl[24].r.part0[16] , 
	\sa_ctrl[24].r.part0[15] , \sa_ctrl[24].r.part0[14] , 
	\sa_ctrl[24].r.part0[13] , \sa_ctrl[24].r.part0[12] , 
	\sa_ctrl[24].r.part0[11] , \sa_ctrl[24].r.part0[10] , 
	\sa_ctrl[24].r.part0[9] , \sa_ctrl[24].r.part0[8] , 
	\sa_ctrl[24].r.part0[7] , \sa_ctrl[24].r.part0[6] , 
	\sa_ctrl[24].r.part0[5] , \sa_ctrl[24].r.part0[4] , 
	\sa_ctrl[24].r.part0[3] , \sa_ctrl[24].r.part0[2] , 
	\sa_ctrl[24].r.part0[1] , \sa_ctrl[24].r.part0[0] , 
	\sa_ctrl[23].r.part0[31] , \sa_ctrl[23].r.part0[30] , 
	\sa_ctrl[23].r.part0[29] , \sa_ctrl[23].r.part0[28] , 
	\sa_ctrl[23].r.part0[27] , \sa_ctrl[23].r.part0[26] , 
	\sa_ctrl[23].r.part0[25] , \sa_ctrl[23].r.part0[24] , 
	\sa_ctrl[23].r.part0[23] , \sa_ctrl[23].r.part0[22] , 
	\sa_ctrl[23].r.part0[21] , \sa_ctrl[23].r.part0[20] , 
	\sa_ctrl[23].r.part0[19] , \sa_ctrl[23].r.part0[18] , 
	\sa_ctrl[23].r.part0[17] , \sa_ctrl[23].r.part0[16] , 
	\sa_ctrl[23].r.part0[15] , \sa_ctrl[23].r.part0[14] , 
	\sa_ctrl[23].r.part0[13] , \sa_ctrl[23].r.part0[12] , 
	\sa_ctrl[23].r.part0[11] , \sa_ctrl[23].r.part0[10] , 
	\sa_ctrl[23].r.part0[9] , \sa_ctrl[23].r.part0[8] , 
	\sa_ctrl[23].r.part0[7] , \sa_ctrl[23].r.part0[6] , 
	\sa_ctrl[23].r.part0[5] , \sa_ctrl[23].r.part0[4] , 
	\sa_ctrl[23].r.part0[3] , \sa_ctrl[23].r.part0[2] , 
	\sa_ctrl[23].r.part0[1] , \sa_ctrl[23].r.part0[0] , 
	\sa_ctrl[22].r.part0[31] , \sa_ctrl[22].r.part0[30] , 
	\sa_ctrl[22].r.part0[29] , \sa_ctrl[22].r.part0[28] , 
	\sa_ctrl[22].r.part0[27] , \sa_ctrl[22].r.part0[26] , 
	\sa_ctrl[22].r.part0[25] , \sa_ctrl[22].r.part0[24] , 
	\sa_ctrl[22].r.part0[23] , \sa_ctrl[22].r.part0[22] , 
	\sa_ctrl[22].r.part0[21] , \sa_ctrl[22].r.part0[20] , 
	\sa_ctrl[22].r.part0[19] , \sa_ctrl[22].r.part0[18] , 
	\sa_ctrl[22].r.part0[17] , \sa_ctrl[22].r.part0[16] , 
	\sa_ctrl[22].r.part0[15] , \sa_ctrl[22].r.part0[14] , 
	\sa_ctrl[22].r.part0[13] , \sa_ctrl[22].r.part0[12] , 
	\sa_ctrl[22].r.part0[11] , \sa_ctrl[22].r.part0[10] , 
	\sa_ctrl[22].r.part0[9] , \sa_ctrl[22].r.part0[8] , 
	\sa_ctrl[22].r.part0[7] , \sa_ctrl[22].r.part0[6] , 
	\sa_ctrl[22].r.part0[5] , \sa_ctrl[22].r.part0[4] , 
	\sa_ctrl[22].r.part0[3] , \sa_ctrl[22].r.part0[2] , 
	\sa_ctrl[22].r.part0[1] , \sa_ctrl[22].r.part0[0] , 
	\sa_ctrl[21].r.part0[31] , \sa_ctrl[21].r.part0[30] , 
	\sa_ctrl[21].r.part0[29] , \sa_ctrl[21].r.part0[28] , 
	\sa_ctrl[21].r.part0[27] , \sa_ctrl[21].r.part0[26] , 
	\sa_ctrl[21].r.part0[25] , \sa_ctrl[21].r.part0[24] , 
	\sa_ctrl[21].r.part0[23] , \sa_ctrl[21].r.part0[22] , 
	\sa_ctrl[21].r.part0[21] , \sa_ctrl[21].r.part0[20] , 
	\sa_ctrl[21].r.part0[19] , \sa_ctrl[21].r.part0[18] , 
	\sa_ctrl[21].r.part0[17] , \sa_ctrl[21].r.part0[16] , 
	\sa_ctrl[21].r.part0[15] , \sa_ctrl[21].r.part0[14] , 
	\sa_ctrl[21].r.part0[13] , \sa_ctrl[21].r.part0[12] , 
	\sa_ctrl[21].r.part0[11] , \sa_ctrl[21].r.part0[10] , 
	\sa_ctrl[21].r.part0[9] , \sa_ctrl[21].r.part0[8] , 
	\sa_ctrl[21].r.part0[7] , \sa_ctrl[21].r.part0[6] , 
	\sa_ctrl[21].r.part0[5] , \sa_ctrl[21].r.part0[4] , 
	\sa_ctrl[21].r.part0[3] , \sa_ctrl[21].r.part0[2] , 
	\sa_ctrl[21].r.part0[1] , \sa_ctrl[21].r.part0[0] , 
	\sa_ctrl[20].r.part0[31] , \sa_ctrl[20].r.part0[30] , 
	\sa_ctrl[20].r.part0[29] , \sa_ctrl[20].r.part0[28] , 
	\sa_ctrl[20].r.part0[27] , \sa_ctrl[20].r.part0[26] , 
	\sa_ctrl[20].r.part0[25] , \sa_ctrl[20].r.part0[24] , 
	\sa_ctrl[20].r.part0[23] , \sa_ctrl[20].r.part0[22] , 
	\sa_ctrl[20].r.part0[21] , \sa_ctrl[20].r.part0[20] , 
	\sa_ctrl[20].r.part0[19] , \sa_ctrl[20].r.part0[18] , 
	\sa_ctrl[20].r.part0[17] , \sa_ctrl[20].r.part0[16] , 
	\sa_ctrl[20].r.part0[15] , \sa_ctrl[20].r.part0[14] , 
	\sa_ctrl[20].r.part0[13] , \sa_ctrl[20].r.part0[12] , 
	\sa_ctrl[20].r.part0[11] , \sa_ctrl[20].r.part0[10] , 
	\sa_ctrl[20].r.part0[9] , \sa_ctrl[20].r.part0[8] , 
	\sa_ctrl[20].r.part0[7] , \sa_ctrl[20].r.part0[6] , 
	\sa_ctrl[20].r.part0[5] , \sa_ctrl[20].r.part0[4] , 
	\sa_ctrl[20].r.part0[3] , \sa_ctrl[20].r.part0[2] , 
	\sa_ctrl[20].r.part0[1] , \sa_ctrl[20].r.part0[0] , 
	\sa_ctrl[19].r.part0[31] , \sa_ctrl[19].r.part0[30] , 
	\sa_ctrl[19].r.part0[29] , \sa_ctrl[19].r.part0[28] , 
	\sa_ctrl[19].r.part0[27] , \sa_ctrl[19].r.part0[26] , 
	\sa_ctrl[19].r.part0[25] , \sa_ctrl[19].r.part0[24] , 
	\sa_ctrl[19].r.part0[23] , \sa_ctrl[19].r.part0[22] , 
	\sa_ctrl[19].r.part0[21] , \sa_ctrl[19].r.part0[20] , 
	\sa_ctrl[19].r.part0[19] , \sa_ctrl[19].r.part0[18] , 
	\sa_ctrl[19].r.part0[17] , \sa_ctrl[19].r.part0[16] , 
	\sa_ctrl[19].r.part0[15] , \sa_ctrl[19].r.part0[14] , 
	\sa_ctrl[19].r.part0[13] , \sa_ctrl[19].r.part0[12] , 
	\sa_ctrl[19].r.part0[11] , \sa_ctrl[19].r.part0[10] , 
	\sa_ctrl[19].r.part0[9] , \sa_ctrl[19].r.part0[8] , 
	\sa_ctrl[19].r.part0[7] , \sa_ctrl[19].r.part0[6] , 
	\sa_ctrl[19].r.part0[5] , \sa_ctrl[19].r.part0[4] , 
	\sa_ctrl[19].r.part0[3] , \sa_ctrl[19].r.part0[2] , 
	\sa_ctrl[19].r.part0[1] , \sa_ctrl[19].r.part0[0] , 
	\sa_ctrl[18].r.part0[31] , \sa_ctrl[18].r.part0[30] , 
	\sa_ctrl[18].r.part0[29] , \sa_ctrl[18].r.part0[28] , 
	\sa_ctrl[18].r.part0[27] , \sa_ctrl[18].r.part0[26] , 
	\sa_ctrl[18].r.part0[25] , \sa_ctrl[18].r.part0[24] , 
	\sa_ctrl[18].r.part0[23] , \sa_ctrl[18].r.part0[22] , 
	\sa_ctrl[18].r.part0[21] , \sa_ctrl[18].r.part0[20] , 
	\sa_ctrl[18].r.part0[19] , \sa_ctrl[18].r.part0[18] , 
	\sa_ctrl[18].r.part0[17] , \sa_ctrl[18].r.part0[16] , 
	\sa_ctrl[18].r.part0[15] , \sa_ctrl[18].r.part0[14] , 
	\sa_ctrl[18].r.part0[13] , \sa_ctrl[18].r.part0[12] , 
	\sa_ctrl[18].r.part0[11] , \sa_ctrl[18].r.part0[10] , 
	\sa_ctrl[18].r.part0[9] , \sa_ctrl[18].r.part0[8] , 
	\sa_ctrl[18].r.part0[7] , \sa_ctrl[18].r.part0[6] , 
	\sa_ctrl[18].r.part0[5] , \sa_ctrl[18].r.part0[4] , 
	\sa_ctrl[18].r.part0[3] , \sa_ctrl[18].r.part0[2] , 
	\sa_ctrl[18].r.part0[1] , \sa_ctrl[18].r.part0[0] , 
	\sa_ctrl[17].r.part0[31] , \sa_ctrl[17].r.part0[30] , 
	\sa_ctrl[17].r.part0[29] , \sa_ctrl[17].r.part0[28] , 
	\sa_ctrl[17].r.part0[27] , \sa_ctrl[17].r.part0[26] , 
	\sa_ctrl[17].r.part0[25] , \sa_ctrl[17].r.part0[24] , 
	\sa_ctrl[17].r.part0[23] , \sa_ctrl[17].r.part0[22] , 
	\sa_ctrl[17].r.part0[21] , \sa_ctrl[17].r.part0[20] , 
	\sa_ctrl[17].r.part0[19] , \sa_ctrl[17].r.part0[18] , 
	\sa_ctrl[17].r.part0[17] , \sa_ctrl[17].r.part0[16] , 
	\sa_ctrl[17].r.part0[15] , \sa_ctrl[17].r.part0[14] , 
	\sa_ctrl[17].r.part0[13] , \sa_ctrl[17].r.part0[12] , 
	\sa_ctrl[17].r.part0[11] , \sa_ctrl[17].r.part0[10] , 
	\sa_ctrl[17].r.part0[9] , \sa_ctrl[17].r.part0[8] , 
	\sa_ctrl[17].r.part0[7] , \sa_ctrl[17].r.part0[6] , 
	\sa_ctrl[17].r.part0[5] , \sa_ctrl[17].r.part0[4] , 
	\sa_ctrl[17].r.part0[3] , \sa_ctrl[17].r.part0[2] , 
	\sa_ctrl[17].r.part0[1] , \sa_ctrl[17].r.part0[0] , 
	\sa_ctrl[16].r.part0[31] , \sa_ctrl[16].r.part0[30] , 
	\sa_ctrl[16].r.part0[29] , \sa_ctrl[16].r.part0[28] , 
	\sa_ctrl[16].r.part0[27] , \sa_ctrl[16].r.part0[26] , 
	\sa_ctrl[16].r.part0[25] , \sa_ctrl[16].r.part0[24] , 
	\sa_ctrl[16].r.part0[23] , \sa_ctrl[16].r.part0[22] , 
	\sa_ctrl[16].r.part0[21] , \sa_ctrl[16].r.part0[20] , 
	\sa_ctrl[16].r.part0[19] , \sa_ctrl[16].r.part0[18] , 
	\sa_ctrl[16].r.part0[17] , \sa_ctrl[16].r.part0[16] , 
	\sa_ctrl[16].r.part0[15] , \sa_ctrl[16].r.part0[14] , 
	\sa_ctrl[16].r.part0[13] , \sa_ctrl[16].r.part0[12] , 
	\sa_ctrl[16].r.part0[11] , \sa_ctrl[16].r.part0[10] , 
	\sa_ctrl[16].r.part0[9] , \sa_ctrl[16].r.part0[8] , 
	\sa_ctrl[16].r.part0[7] , \sa_ctrl[16].r.part0[6] , 
	\sa_ctrl[16].r.part0[5] , \sa_ctrl[16].r.part0[4] , 
	\sa_ctrl[16].r.part0[3] , \sa_ctrl[16].r.part0[2] , 
	\sa_ctrl[16].r.part0[1] , \sa_ctrl[16].r.part0[0] , 
	\sa_ctrl[15].r.part0[31] , \sa_ctrl[15].r.part0[30] , 
	\sa_ctrl[15].r.part0[29] , \sa_ctrl[15].r.part0[28] , 
	\sa_ctrl[15].r.part0[27] , \sa_ctrl[15].r.part0[26] , 
	\sa_ctrl[15].r.part0[25] , \sa_ctrl[15].r.part0[24] , 
	\sa_ctrl[15].r.part0[23] , \sa_ctrl[15].r.part0[22] , 
	\sa_ctrl[15].r.part0[21] , \sa_ctrl[15].r.part0[20] , 
	\sa_ctrl[15].r.part0[19] , \sa_ctrl[15].r.part0[18] , 
	\sa_ctrl[15].r.part0[17] , \sa_ctrl[15].r.part0[16] , 
	\sa_ctrl[15].r.part0[15] , \sa_ctrl[15].r.part0[14] , 
	\sa_ctrl[15].r.part0[13] , \sa_ctrl[15].r.part0[12] , 
	\sa_ctrl[15].r.part0[11] , \sa_ctrl[15].r.part0[10] , 
	\sa_ctrl[15].r.part0[9] , \sa_ctrl[15].r.part0[8] , 
	\sa_ctrl[15].r.part0[7] , \sa_ctrl[15].r.part0[6] , 
	\sa_ctrl[15].r.part0[5] , \sa_ctrl[15].r.part0[4] , 
	\sa_ctrl[15].r.part0[3] , \sa_ctrl[15].r.part0[2] , 
	\sa_ctrl[15].r.part0[1] , \sa_ctrl[15].r.part0[0] , 
	\sa_ctrl[14].r.part0[31] , \sa_ctrl[14].r.part0[30] , 
	\sa_ctrl[14].r.part0[29] , \sa_ctrl[14].r.part0[28] , 
	\sa_ctrl[14].r.part0[27] , \sa_ctrl[14].r.part0[26] , 
	\sa_ctrl[14].r.part0[25] , \sa_ctrl[14].r.part0[24] , 
	\sa_ctrl[14].r.part0[23] , \sa_ctrl[14].r.part0[22] , 
	\sa_ctrl[14].r.part0[21] , \sa_ctrl[14].r.part0[20] , 
	\sa_ctrl[14].r.part0[19] , \sa_ctrl[14].r.part0[18] , 
	\sa_ctrl[14].r.part0[17] , \sa_ctrl[14].r.part0[16] , 
	\sa_ctrl[14].r.part0[15] , \sa_ctrl[14].r.part0[14] , 
	\sa_ctrl[14].r.part0[13] , \sa_ctrl[14].r.part0[12] , 
	\sa_ctrl[14].r.part0[11] , \sa_ctrl[14].r.part0[10] , 
	\sa_ctrl[14].r.part0[9] , \sa_ctrl[14].r.part0[8] , 
	\sa_ctrl[14].r.part0[7] , \sa_ctrl[14].r.part0[6] , 
	\sa_ctrl[14].r.part0[5] , \sa_ctrl[14].r.part0[4] , 
	\sa_ctrl[14].r.part0[3] , \sa_ctrl[14].r.part0[2] , 
	\sa_ctrl[14].r.part0[1] , \sa_ctrl[14].r.part0[0] , 
	\sa_ctrl[13].r.part0[31] , \sa_ctrl[13].r.part0[30] , 
	\sa_ctrl[13].r.part0[29] , \sa_ctrl[13].r.part0[28] , 
	\sa_ctrl[13].r.part0[27] , \sa_ctrl[13].r.part0[26] , 
	\sa_ctrl[13].r.part0[25] , \sa_ctrl[13].r.part0[24] , 
	\sa_ctrl[13].r.part0[23] , \sa_ctrl[13].r.part0[22] , 
	\sa_ctrl[13].r.part0[21] , \sa_ctrl[13].r.part0[20] , 
	\sa_ctrl[13].r.part0[19] , \sa_ctrl[13].r.part0[18] , 
	\sa_ctrl[13].r.part0[17] , \sa_ctrl[13].r.part0[16] , 
	\sa_ctrl[13].r.part0[15] , \sa_ctrl[13].r.part0[14] , 
	\sa_ctrl[13].r.part0[13] , \sa_ctrl[13].r.part0[12] , 
	\sa_ctrl[13].r.part0[11] , \sa_ctrl[13].r.part0[10] , 
	\sa_ctrl[13].r.part0[9] , \sa_ctrl[13].r.part0[8] , 
	\sa_ctrl[13].r.part0[7] , \sa_ctrl[13].r.part0[6] , 
	\sa_ctrl[13].r.part0[5] , \sa_ctrl[13].r.part0[4] , 
	\sa_ctrl[13].r.part0[3] , \sa_ctrl[13].r.part0[2] , 
	\sa_ctrl[13].r.part0[1] , \sa_ctrl[13].r.part0[0] , 
	\sa_ctrl[12].r.part0[31] , \sa_ctrl[12].r.part0[30] , 
	\sa_ctrl[12].r.part0[29] , \sa_ctrl[12].r.part0[28] , 
	\sa_ctrl[12].r.part0[27] , \sa_ctrl[12].r.part0[26] , 
	\sa_ctrl[12].r.part0[25] , \sa_ctrl[12].r.part0[24] , 
	\sa_ctrl[12].r.part0[23] , \sa_ctrl[12].r.part0[22] , 
	\sa_ctrl[12].r.part0[21] , \sa_ctrl[12].r.part0[20] , 
	\sa_ctrl[12].r.part0[19] , \sa_ctrl[12].r.part0[18] , 
	\sa_ctrl[12].r.part0[17] , \sa_ctrl[12].r.part0[16] , 
	\sa_ctrl[12].r.part0[15] , \sa_ctrl[12].r.part0[14] , 
	\sa_ctrl[12].r.part0[13] , \sa_ctrl[12].r.part0[12] , 
	\sa_ctrl[12].r.part0[11] , \sa_ctrl[12].r.part0[10] , 
	\sa_ctrl[12].r.part0[9] , \sa_ctrl[12].r.part0[8] , 
	\sa_ctrl[12].r.part0[7] , \sa_ctrl[12].r.part0[6] , 
	\sa_ctrl[12].r.part0[5] , \sa_ctrl[12].r.part0[4] , 
	\sa_ctrl[12].r.part0[3] , \sa_ctrl[12].r.part0[2] , 
	\sa_ctrl[12].r.part0[1] , \sa_ctrl[12].r.part0[0] , 
	\sa_ctrl[11].r.part0[31] , \sa_ctrl[11].r.part0[30] , 
	\sa_ctrl[11].r.part0[29] , \sa_ctrl[11].r.part0[28] , 
	\sa_ctrl[11].r.part0[27] , \sa_ctrl[11].r.part0[26] , 
	\sa_ctrl[11].r.part0[25] , \sa_ctrl[11].r.part0[24] , 
	\sa_ctrl[11].r.part0[23] , \sa_ctrl[11].r.part0[22] , 
	\sa_ctrl[11].r.part0[21] , \sa_ctrl[11].r.part0[20] , 
	\sa_ctrl[11].r.part0[19] , \sa_ctrl[11].r.part0[18] , 
	\sa_ctrl[11].r.part0[17] , \sa_ctrl[11].r.part0[16] , 
	\sa_ctrl[11].r.part0[15] , \sa_ctrl[11].r.part0[14] , 
	\sa_ctrl[11].r.part0[13] , \sa_ctrl[11].r.part0[12] , 
	\sa_ctrl[11].r.part0[11] , \sa_ctrl[11].r.part0[10] , 
	\sa_ctrl[11].r.part0[9] , \sa_ctrl[11].r.part0[8] , 
	\sa_ctrl[11].r.part0[7] , \sa_ctrl[11].r.part0[6] , 
	\sa_ctrl[11].r.part0[5] , \sa_ctrl[11].r.part0[4] , 
	\sa_ctrl[11].r.part0[3] , \sa_ctrl[11].r.part0[2] , 
	\sa_ctrl[11].r.part0[1] , \sa_ctrl[11].r.part0[0] , 
	\sa_ctrl[10].r.part0[31] , \sa_ctrl[10].r.part0[30] , 
	\sa_ctrl[10].r.part0[29] , \sa_ctrl[10].r.part0[28] , 
	\sa_ctrl[10].r.part0[27] , \sa_ctrl[10].r.part0[26] , 
	\sa_ctrl[10].r.part0[25] , \sa_ctrl[10].r.part0[24] , 
	\sa_ctrl[10].r.part0[23] , \sa_ctrl[10].r.part0[22] , 
	\sa_ctrl[10].r.part0[21] , \sa_ctrl[10].r.part0[20] , 
	\sa_ctrl[10].r.part0[19] , \sa_ctrl[10].r.part0[18] , 
	\sa_ctrl[10].r.part0[17] , \sa_ctrl[10].r.part0[16] , 
	\sa_ctrl[10].r.part0[15] , \sa_ctrl[10].r.part0[14] , 
	\sa_ctrl[10].r.part0[13] , \sa_ctrl[10].r.part0[12] , 
	\sa_ctrl[10].r.part0[11] , \sa_ctrl[10].r.part0[10] , 
	\sa_ctrl[10].r.part0[9] , \sa_ctrl[10].r.part0[8] , 
	\sa_ctrl[10].r.part0[7] , \sa_ctrl[10].r.part0[6] , 
	\sa_ctrl[10].r.part0[5] , \sa_ctrl[10].r.part0[4] , 
	\sa_ctrl[10].r.part0[3] , \sa_ctrl[10].r.part0[2] , 
	\sa_ctrl[10].r.part0[1] , \sa_ctrl[10].r.part0[0] , 
	\sa_ctrl[9].r.part0[31] , \sa_ctrl[9].r.part0[30] , 
	\sa_ctrl[9].r.part0[29] , \sa_ctrl[9].r.part0[28] , 
	\sa_ctrl[9].r.part0[27] , \sa_ctrl[9].r.part0[26] , 
	\sa_ctrl[9].r.part0[25] , \sa_ctrl[9].r.part0[24] , 
	\sa_ctrl[9].r.part0[23] , \sa_ctrl[9].r.part0[22] , 
	\sa_ctrl[9].r.part0[21] , \sa_ctrl[9].r.part0[20] , 
	\sa_ctrl[9].r.part0[19] , \sa_ctrl[9].r.part0[18] , 
	\sa_ctrl[9].r.part0[17] , \sa_ctrl[9].r.part0[16] , 
	\sa_ctrl[9].r.part0[15] , \sa_ctrl[9].r.part0[14] , 
	\sa_ctrl[9].r.part0[13] , \sa_ctrl[9].r.part0[12] , 
	\sa_ctrl[9].r.part0[11] , \sa_ctrl[9].r.part0[10] , 
	\sa_ctrl[9].r.part0[9] , \sa_ctrl[9].r.part0[8] , 
	\sa_ctrl[9].r.part0[7] , \sa_ctrl[9].r.part0[6] , 
	\sa_ctrl[9].r.part0[5] , \sa_ctrl[9].r.part0[4] , 
	\sa_ctrl[9].r.part0[3] , \sa_ctrl[9].r.part0[2] , 
	\sa_ctrl[9].r.part0[1] , \sa_ctrl[9].r.part0[0] , 
	\sa_ctrl[8].r.part0[31] , \sa_ctrl[8].r.part0[30] , 
	\sa_ctrl[8].r.part0[29] , \sa_ctrl[8].r.part0[28] , 
	\sa_ctrl[8].r.part0[27] , \sa_ctrl[8].r.part0[26] , 
	\sa_ctrl[8].r.part0[25] , \sa_ctrl[8].r.part0[24] , 
	\sa_ctrl[8].r.part0[23] , \sa_ctrl[8].r.part0[22] , 
	\sa_ctrl[8].r.part0[21] , \sa_ctrl[8].r.part0[20] , 
	\sa_ctrl[8].r.part0[19] , \sa_ctrl[8].r.part0[18] , 
	\sa_ctrl[8].r.part0[17] , \sa_ctrl[8].r.part0[16] , 
	\sa_ctrl[8].r.part0[15] , \sa_ctrl[8].r.part0[14] , 
	\sa_ctrl[8].r.part0[13] , \sa_ctrl[8].r.part0[12] , 
	\sa_ctrl[8].r.part0[11] , \sa_ctrl[8].r.part0[10] , 
	\sa_ctrl[8].r.part0[9] , \sa_ctrl[8].r.part0[8] , 
	\sa_ctrl[8].r.part0[7] , \sa_ctrl[8].r.part0[6] , 
	\sa_ctrl[8].r.part0[5] , \sa_ctrl[8].r.part0[4] , 
	\sa_ctrl[8].r.part0[3] , \sa_ctrl[8].r.part0[2] , 
	\sa_ctrl[8].r.part0[1] , \sa_ctrl[8].r.part0[0] , 
	\sa_ctrl[7].r.part0[31] , \sa_ctrl[7].r.part0[30] , 
	\sa_ctrl[7].r.part0[29] , \sa_ctrl[7].r.part0[28] , 
	\sa_ctrl[7].r.part0[27] , \sa_ctrl[7].r.part0[26] , 
	\sa_ctrl[7].r.part0[25] , \sa_ctrl[7].r.part0[24] , 
	\sa_ctrl[7].r.part0[23] , \sa_ctrl[7].r.part0[22] , 
	\sa_ctrl[7].r.part0[21] , \sa_ctrl[7].r.part0[20] , 
	\sa_ctrl[7].r.part0[19] , \sa_ctrl[7].r.part0[18] , 
	\sa_ctrl[7].r.part0[17] , \sa_ctrl[7].r.part0[16] , 
	\sa_ctrl[7].r.part0[15] , \sa_ctrl[7].r.part0[14] , 
	\sa_ctrl[7].r.part0[13] , \sa_ctrl[7].r.part0[12] , 
	\sa_ctrl[7].r.part0[11] , \sa_ctrl[7].r.part0[10] , 
	\sa_ctrl[7].r.part0[9] , \sa_ctrl[7].r.part0[8] , 
	\sa_ctrl[7].r.part0[7] , \sa_ctrl[7].r.part0[6] , 
	\sa_ctrl[7].r.part0[5] , \sa_ctrl[7].r.part0[4] , 
	\sa_ctrl[7].r.part0[3] , \sa_ctrl[7].r.part0[2] , 
	\sa_ctrl[7].r.part0[1] , \sa_ctrl[7].r.part0[0] , 
	\sa_ctrl[6].r.part0[31] , \sa_ctrl[6].r.part0[30] , 
	\sa_ctrl[6].r.part0[29] , \sa_ctrl[6].r.part0[28] , 
	\sa_ctrl[6].r.part0[27] , \sa_ctrl[6].r.part0[26] , 
	\sa_ctrl[6].r.part0[25] , \sa_ctrl[6].r.part0[24] , 
	\sa_ctrl[6].r.part0[23] , \sa_ctrl[6].r.part0[22] , 
	\sa_ctrl[6].r.part0[21] , \sa_ctrl[6].r.part0[20] , 
	\sa_ctrl[6].r.part0[19] , \sa_ctrl[6].r.part0[18] , 
	\sa_ctrl[6].r.part0[17] , \sa_ctrl[6].r.part0[16] , 
	\sa_ctrl[6].r.part0[15] , \sa_ctrl[6].r.part0[14] , 
	\sa_ctrl[6].r.part0[13] , \sa_ctrl[6].r.part0[12] , 
	\sa_ctrl[6].r.part0[11] , \sa_ctrl[6].r.part0[10] , 
	\sa_ctrl[6].r.part0[9] , \sa_ctrl[6].r.part0[8] , 
	\sa_ctrl[6].r.part0[7] , \sa_ctrl[6].r.part0[6] , 
	\sa_ctrl[6].r.part0[5] , \sa_ctrl[6].r.part0[4] , 
	\sa_ctrl[6].r.part0[3] , \sa_ctrl[6].r.part0[2] , 
	\sa_ctrl[6].r.part0[1] , \sa_ctrl[6].r.part0[0] , 
	\sa_ctrl[5].r.part0[31] , \sa_ctrl[5].r.part0[30] , 
	\sa_ctrl[5].r.part0[29] , \sa_ctrl[5].r.part0[28] , 
	\sa_ctrl[5].r.part0[27] , \sa_ctrl[5].r.part0[26] , 
	\sa_ctrl[5].r.part0[25] , \sa_ctrl[5].r.part0[24] , 
	\sa_ctrl[5].r.part0[23] , \sa_ctrl[5].r.part0[22] , 
	\sa_ctrl[5].r.part0[21] , \sa_ctrl[5].r.part0[20] , 
	\sa_ctrl[5].r.part0[19] , \sa_ctrl[5].r.part0[18] , 
	\sa_ctrl[5].r.part0[17] , \sa_ctrl[5].r.part0[16] , 
	\sa_ctrl[5].r.part0[15] , \sa_ctrl[5].r.part0[14] , 
	\sa_ctrl[5].r.part0[13] , \sa_ctrl[5].r.part0[12] , 
	\sa_ctrl[5].r.part0[11] , \sa_ctrl[5].r.part0[10] , 
	\sa_ctrl[5].r.part0[9] , \sa_ctrl[5].r.part0[8] , 
	\sa_ctrl[5].r.part0[7] , \sa_ctrl[5].r.part0[6] , 
	\sa_ctrl[5].r.part0[5] , \sa_ctrl[5].r.part0[4] , 
	\sa_ctrl[5].r.part0[3] , \sa_ctrl[5].r.part0[2] , 
	\sa_ctrl[5].r.part0[1] , \sa_ctrl[5].r.part0[0] , 
	\sa_ctrl[4].r.part0[31] , \sa_ctrl[4].r.part0[30] , 
	\sa_ctrl[4].r.part0[29] , \sa_ctrl[4].r.part0[28] , 
	\sa_ctrl[4].r.part0[27] , \sa_ctrl[4].r.part0[26] , 
	\sa_ctrl[4].r.part0[25] , \sa_ctrl[4].r.part0[24] , 
	\sa_ctrl[4].r.part0[23] , \sa_ctrl[4].r.part0[22] , 
	\sa_ctrl[4].r.part0[21] , \sa_ctrl[4].r.part0[20] , 
	\sa_ctrl[4].r.part0[19] , \sa_ctrl[4].r.part0[18] , 
	\sa_ctrl[4].r.part0[17] , \sa_ctrl[4].r.part0[16] , 
	\sa_ctrl[4].r.part0[15] , \sa_ctrl[4].r.part0[14] , 
	\sa_ctrl[4].r.part0[13] , \sa_ctrl[4].r.part0[12] , 
	\sa_ctrl[4].r.part0[11] , \sa_ctrl[4].r.part0[10] , 
	\sa_ctrl[4].r.part0[9] , \sa_ctrl[4].r.part0[8] , 
	\sa_ctrl[4].r.part0[7] , \sa_ctrl[4].r.part0[6] , 
	\sa_ctrl[4].r.part0[5] , \sa_ctrl[4].r.part0[4] , 
	\sa_ctrl[4].r.part0[3] , \sa_ctrl[4].r.part0[2] , 
	\sa_ctrl[4].r.part0[1] , \sa_ctrl[4].r.part0[0] , 
	\sa_ctrl[3].r.part0[31] , \sa_ctrl[3].r.part0[30] , 
	\sa_ctrl[3].r.part0[29] , \sa_ctrl[3].r.part0[28] , 
	\sa_ctrl[3].r.part0[27] , \sa_ctrl[3].r.part0[26] , 
	\sa_ctrl[3].r.part0[25] , \sa_ctrl[3].r.part0[24] , 
	\sa_ctrl[3].r.part0[23] , \sa_ctrl[3].r.part0[22] , 
	\sa_ctrl[3].r.part0[21] , \sa_ctrl[3].r.part0[20] , 
	\sa_ctrl[3].r.part0[19] , \sa_ctrl[3].r.part0[18] , 
	\sa_ctrl[3].r.part0[17] , \sa_ctrl[3].r.part0[16] , 
	\sa_ctrl[3].r.part0[15] , \sa_ctrl[3].r.part0[14] , 
	\sa_ctrl[3].r.part0[13] , \sa_ctrl[3].r.part0[12] , 
	\sa_ctrl[3].r.part0[11] , \sa_ctrl[3].r.part0[10] , 
	\sa_ctrl[3].r.part0[9] , \sa_ctrl[3].r.part0[8] , 
	\sa_ctrl[3].r.part0[7] , \sa_ctrl[3].r.part0[6] , 
	\sa_ctrl[3].r.part0[5] , \sa_ctrl[3].r.part0[4] , 
	\sa_ctrl[3].r.part0[3] , \sa_ctrl[3].r.part0[2] , 
	\sa_ctrl[3].r.part0[1] , \sa_ctrl[3].r.part0[0] , 
	\sa_ctrl[2].r.part0[31] , \sa_ctrl[2].r.part0[30] , 
	\sa_ctrl[2].r.part0[29] , \sa_ctrl[2].r.part0[28] , 
	\sa_ctrl[2].r.part0[27] , \sa_ctrl[2].r.part0[26] , 
	\sa_ctrl[2].r.part0[25] , \sa_ctrl[2].r.part0[24] , 
	\sa_ctrl[2].r.part0[23] , \sa_ctrl[2].r.part0[22] , 
	\sa_ctrl[2].r.part0[21] , \sa_ctrl[2].r.part0[20] , 
	\sa_ctrl[2].r.part0[19] , \sa_ctrl[2].r.part0[18] , 
	\sa_ctrl[2].r.part0[17] , \sa_ctrl[2].r.part0[16] , 
	\sa_ctrl[2].r.part0[15] , \sa_ctrl[2].r.part0[14] , 
	\sa_ctrl[2].r.part0[13] , \sa_ctrl[2].r.part0[12] , 
	\sa_ctrl[2].r.part0[11] , \sa_ctrl[2].r.part0[10] , 
	\sa_ctrl[2].r.part0[9] , \sa_ctrl[2].r.part0[8] , 
	\sa_ctrl[2].r.part0[7] , \sa_ctrl[2].r.part0[6] , 
	\sa_ctrl[2].r.part0[5] , \sa_ctrl[2].r.part0[4] , 
	\sa_ctrl[2].r.part0[3] , \sa_ctrl[2].r.part0[2] , 
	\sa_ctrl[2].r.part0[1] , \sa_ctrl[2].r.part0[0] , 
	\sa_ctrl[1].r.part0[31] , \sa_ctrl[1].r.part0[30] , 
	\sa_ctrl[1].r.part0[29] , \sa_ctrl[1].r.part0[28] , 
	\sa_ctrl[1].r.part0[27] , \sa_ctrl[1].r.part0[26] , 
	\sa_ctrl[1].r.part0[25] , \sa_ctrl[1].r.part0[24] , 
	\sa_ctrl[1].r.part0[23] , \sa_ctrl[1].r.part0[22] , 
	\sa_ctrl[1].r.part0[21] , \sa_ctrl[1].r.part0[20] , 
	\sa_ctrl[1].r.part0[19] , \sa_ctrl[1].r.part0[18] , 
	\sa_ctrl[1].r.part0[17] , \sa_ctrl[1].r.part0[16] , 
	\sa_ctrl[1].r.part0[15] , \sa_ctrl[1].r.part0[14] , 
	\sa_ctrl[1].r.part0[13] , \sa_ctrl[1].r.part0[12] , 
	\sa_ctrl[1].r.part0[11] , \sa_ctrl[1].r.part0[10] , 
	\sa_ctrl[1].r.part0[9] , \sa_ctrl[1].r.part0[8] , 
	\sa_ctrl[1].r.part0[7] , \sa_ctrl[1].r.part0[6] , 
	\sa_ctrl[1].r.part0[5] , \sa_ctrl[1].r.part0[4] , 
	\sa_ctrl[1].r.part0[3] , \sa_ctrl[1].r.part0[2] , 
	\sa_ctrl[1].r.part0[1] , \sa_ctrl[1].r.part0[0] , 
	\sa_ctrl[0].r.part0[31] , \sa_ctrl[0].r.part0[30] , 
	\sa_ctrl[0].r.part0[29] , \sa_ctrl[0].r.part0[28] , 
	\sa_ctrl[0].r.part0[27] , \sa_ctrl[0].r.part0[26] , 
	\sa_ctrl[0].r.part0[25] , \sa_ctrl[0].r.part0[24] , 
	\sa_ctrl[0].r.part0[23] , \sa_ctrl[0].r.part0[22] , 
	\sa_ctrl[0].r.part0[21] , \sa_ctrl[0].r.part0[20] , 
	\sa_ctrl[0].r.part0[19] , \sa_ctrl[0].r.part0[18] , 
	\sa_ctrl[0].r.part0[17] , \sa_ctrl[0].r.part0[16] , 
	\sa_ctrl[0].r.part0[15] , \sa_ctrl[0].r.part0[14] , 
	\sa_ctrl[0].r.part0[13] , \sa_ctrl[0].r.part0[12] , 
	\sa_ctrl[0].r.part0[11] , \sa_ctrl[0].r.part0[10] , 
	\sa_ctrl[0].r.part0[9] , \sa_ctrl[0].r.part0[8] , 
	\sa_ctrl[0].r.part0[7] , \sa_ctrl[0].r.part0[6] , 
	\sa_ctrl[0].r.part0[5] , \sa_ctrl[0].r.part0[4] , 
	\sa_ctrl[0].r.part0[3] , \sa_ctrl[0].r.part0[2] , 
	\sa_ctrl[0].r.part0[1] , \sa_ctrl[0].r.part0[0] } ), 
	debug_kme_ib_tvalid, debug_kme_ib_tlast, debug_kme_ib_tid, 
	debug_kme_ib_tstrb, debug_kme_ib_tuser, debug_kme_ib_tdata, clk, 
	rst_n, ovstb, lvm, mlvm, .rbus_ring_i( {\rbus_ring_i.addr [15], 
	\rbus_ring_i.addr [14], \rbus_ring_i.addr [13], 
	\rbus_ring_i.addr [12], \rbus_ring_i.addr [11], 
	\rbus_ring_i.addr [10], \rbus_ring_i.addr [9], \rbus_ring_i.addr [8], 
	\rbus_ring_i.addr [7], \rbus_ring_i.addr [6], \rbus_ring_i.addr [5], 
	\rbus_ring_i.addr [4], \rbus_ring_i.addr [3], \rbus_ring_i.addr [2], 
	\rbus_ring_i.addr [1], \rbus_ring_i.addr [0], \rbus_ring_i.wr_strb , 
	\rbus_ring_i.wr_data [31], \rbus_ring_i.wr_data [30], 
	\rbus_ring_i.wr_data [29], \rbus_ring_i.wr_data [28], 
	\rbus_ring_i.wr_data [27], \rbus_ring_i.wr_data [26], 
	\rbus_ring_i.wr_data [25], \rbus_ring_i.wr_data [24], 
	\rbus_ring_i.wr_data [23], \rbus_ring_i.wr_data [22], 
	\rbus_ring_i.wr_data [21], \rbus_ring_i.wr_data [20], 
	\rbus_ring_i.wr_data [19], \rbus_ring_i.wr_data [18], 
	\rbus_ring_i.wr_data [17], \rbus_ring_i.wr_data [16], 
	\rbus_ring_i.wr_data [15], \rbus_ring_i.wr_data [14], 
	\rbus_ring_i.wr_data [13], \rbus_ring_i.wr_data [12], 
	\rbus_ring_i.wr_data [11], \rbus_ring_i.wr_data [10], 
	\rbus_ring_i.wr_data [9], \rbus_ring_i.wr_data [8], 
	\rbus_ring_i.wr_data [7], \rbus_ring_i.wr_data [6], 
	\rbus_ring_i.wr_data [5], \rbus_ring_i.wr_data [4], 
	\rbus_ring_i.wr_data [3], \rbus_ring_i.wr_data [2], 
	\rbus_ring_i.wr_data [1], \rbus_ring_i.wr_data [0], 
	\rbus_ring_i.rd_strb , \rbus_ring_i.rd_data [31], 
	\rbus_ring_i.rd_data [30], \rbus_ring_i.rd_data [29], 
	\rbus_ring_i.rd_data [28], \rbus_ring_i.rd_data [27], 
	\rbus_ring_i.rd_data [26], \rbus_ring_i.rd_data [25], 
	\rbus_ring_i.rd_data [24], \rbus_ring_i.rd_data [23], 
	\rbus_ring_i.rd_data [22], \rbus_ring_i.rd_data [21], 
	\rbus_ring_i.rd_data [20], \rbus_ring_i.rd_data [19], 
	\rbus_ring_i.rd_data [18], \rbus_ring_i.rd_data [17], 
	\rbus_ring_i.rd_data [16], \rbus_ring_i.rd_data [15], 
	\rbus_ring_i.rd_data [14], \rbus_ring_i.rd_data [13], 
	\rbus_ring_i.rd_data [12], \rbus_ring_i.rd_data [11], 
	\rbus_ring_i.rd_data [10], \rbus_ring_i.rd_data [9], 
	\rbus_ring_i.rd_data [8], \rbus_ring_i.rd_data [7], 
	\rbus_ring_i.rd_data [6], \rbus_ring_i.rd_data [5], 
	\rbus_ring_i.rd_data [4], \rbus_ring_i.rd_data [3], 
	\rbus_ring_i.rd_data [2], \rbus_ring_i.rd_data [1], 
	\rbus_ring_i.rd_data [0], \rbus_ring_i.ack , \rbus_ring_i.err_ack } ), 
	cfg_start_addr, cfg_end_addr, .kme_cceip0_ob_out_pre( {
	\kme_cceip0_ob_out_pre.tvalid , \kme_cceip0_ob_out_pre.tlast , 
	\kme_cceip0_ob_out_pre.tid [0], \kme_cceip0_ob_out_pre.tstrb [7], 
	\kme_cceip0_ob_out_pre.tstrb [6], \kme_cceip0_ob_out_pre.tstrb [5], 
	\kme_cceip0_ob_out_pre.tstrb [4], \kme_cceip0_ob_out_pre.tstrb [3], 
	\kme_cceip0_ob_out_pre.tstrb [2], \kme_cceip0_ob_out_pre.tstrb [1], 
	\kme_cceip0_ob_out_pre.tstrb [0], \kme_cceip0_ob_out_pre.tuser [7], 
	\kme_cceip0_ob_out_pre.tuser [6], \kme_cceip0_ob_out_pre.tuser [5], 
	\kme_cceip0_ob_out_pre.tuser [4], \kme_cceip0_ob_out_pre.tuser [3], 
	\kme_cceip0_ob_out_pre.tuser [2], \kme_cceip0_ob_out_pre.tuser [1], 
	\kme_cceip0_ob_out_pre.tuser [0], \kme_cceip0_ob_out_pre.tdata [63], 
	\kme_cceip0_ob_out_pre.tdata [62], \kme_cceip0_ob_out_pre.tdata [61], 
	\kme_cceip0_ob_out_pre.tdata [60], \kme_cceip0_ob_out_pre.tdata [59], 
	\kme_cceip0_ob_out_pre.tdata [58], \kme_cceip0_ob_out_pre.tdata [57], 
	\kme_cceip0_ob_out_pre.tdata [56], \kme_cceip0_ob_out_pre.tdata [55], 
	\kme_cceip0_ob_out_pre.tdata [54], \kme_cceip0_ob_out_pre.tdata [53], 
	\kme_cceip0_ob_out_pre.tdata [52], \kme_cceip0_ob_out_pre.tdata [51], 
	\kme_cceip0_ob_out_pre.tdata [50], \kme_cceip0_ob_out_pre.tdata [49], 
	\kme_cceip0_ob_out_pre.tdata [48], \kme_cceip0_ob_out_pre.tdata [47], 
	\kme_cceip0_ob_out_pre.tdata [46], \kme_cceip0_ob_out_pre.tdata [45], 
	\kme_cceip0_ob_out_pre.tdata [44], \kme_cceip0_ob_out_pre.tdata [43], 
	\kme_cceip0_ob_out_pre.tdata [42], \kme_cceip0_ob_out_pre.tdata [41], 
	\kme_cceip0_ob_out_pre.tdata [40], \kme_cceip0_ob_out_pre.tdata [39], 
	\kme_cceip0_ob_out_pre.tdata [38], \kme_cceip0_ob_out_pre.tdata [37], 
	\kme_cceip0_ob_out_pre.tdata [36], \kme_cceip0_ob_out_pre.tdata [35], 
	\kme_cceip0_ob_out_pre.tdata [34], \kme_cceip0_ob_out_pre.tdata [33], 
	\kme_cceip0_ob_out_pre.tdata [32], \kme_cceip0_ob_out_pre.tdata [31], 
	\kme_cceip0_ob_out_pre.tdata [30], \kme_cceip0_ob_out_pre.tdata [29], 
	\kme_cceip0_ob_out_pre.tdata [28], \kme_cceip0_ob_out_pre.tdata [27], 
	\kme_cceip0_ob_out_pre.tdata [26], \kme_cceip0_ob_out_pre.tdata [25], 
	\kme_cceip0_ob_out_pre.tdata [24], \kme_cceip0_ob_out_pre.tdata [23], 
	\kme_cceip0_ob_out_pre.tdata [22], \kme_cceip0_ob_out_pre.tdata [21], 
	\kme_cceip0_ob_out_pre.tdata [20], \kme_cceip0_ob_out_pre.tdata [19], 
	\kme_cceip0_ob_out_pre.tdata [18], \kme_cceip0_ob_out_pre.tdata [17], 
	\kme_cceip0_ob_out_pre.tdata [16], \kme_cceip0_ob_out_pre.tdata [15], 
	\kme_cceip0_ob_out_pre.tdata [14], \kme_cceip0_ob_out_pre.tdata [13], 
	\kme_cceip0_ob_out_pre.tdata [12], \kme_cceip0_ob_out_pre.tdata [11], 
	\kme_cceip0_ob_out_pre.tdata [10], \kme_cceip0_ob_out_pre.tdata [9], 
	\kme_cceip0_ob_out_pre.tdata [8], \kme_cceip0_ob_out_pre.tdata [7], 
	\kme_cceip0_ob_out_pre.tdata [6], \kme_cceip0_ob_out_pre.tdata [5], 
	\kme_cceip0_ob_out_pre.tdata [4], \kme_cceip0_ob_out_pre.tdata [3], 
	\kme_cceip0_ob_out_pre.tdata [2], \kme_cceip0_ob_out_pre.tdata [1], 
	\kme_cceip0_ob_out_pre.tdata [0]} ), .kme_cceip0_ob_in( {
	\kme_cceip0_ob_in.tready } ), .kme_cceip1_ob_out_pre( {
	\kme_cceip1_ob_out_pre.tvalid , \kme_cceip1_ob_out_pre.tlast , 
	\kme_cceip1_ob_out_pre.tid [0], \kme_cceip1_ob_out_pre.tstrb [7], 
	\kme_cceip1_ob_out_pre.tstrb [6], \kme_cceip1_ob_out_pre.tstrb [5], 
	\kme_cceip1_ob_out_pre.tstrb [4], \kme_cceip1_ob_out_pre.tstrb [3], 
	\kme_cceip1_ob_out_pre.tstrb [2], \kme_cceip1_ob_out_pre.tstrb [1], 
	\kme_cceip1_ob_out_pre.tstrb [0], \kme_cceip1_ob_out_pre.tuser [7], 
	\kme_cceip1_ob_out_pre.tuser [6], \kme_cceip1_ob_out_pre.tuser [5], 
	\kme_cceip1_ob_out_pre.tuser [4], \kme_cceip1_ob_out_pre.tuser [3], 
	\kme_cceip1_ob_out_pre.tuser [2], \kme_cceip1_ob_out_pre.tuser [1], 
	\kme_cceip1_ob_out_pre.tuser [0], \kme_cceip1_ob_out_pre.tdata [63], 
	\kme_cceip1_ob_out_pre.tdata [62], \kme_cceip1_ob_out_pre.tdata [61], 
	\kme_cceip1_ob_out_pre.tdata [60], \kme_cceip1_ob_out_pre.tdata [59], 
	\kme_cceip1_ob_out_pre.tdata [58], \kme_cceip1_ob_out_pre.tdata [57], 
	\kme_cceip1_ob_out_pre.tdata [56], \kme_cceip1_ob_out_pre.tdata [55], 
	\kme_cceip1_ob_out_pre.tdata [54], \kme_cceip1_ob_out_pre.tdata [53], 
	\kme_cceip1_ob_out_pre.tdata [52], \kme_cceip1_ob_out_pre.tdata [51], 
	\kme_cceip1_ob_out_pre.tdata [50], \kme_cceip1_ob_out_pre.tdata [49], 
	\kme_cceip1_ob_out_pre.tdata [48], \kme_cceip1_ob_out_pre.tdata [47], 
	\kme_cceip1_ob_out_pre.tdata [46], \kme_cceip1_ob_out_pre.tdata [45], 
	\kme_cceip1_ob_out_pre.tdata [44], \kme_cceip1_ob_out_pre.tdata [43], 
	\kme_cceip1_ob_out_pre.tdata [42], \kme_cceip1_ob_out_pre.tdata [41], 
	\kme_cceip1_ob_out_pre.tdata [40], \kme_cceip1_ob_out_pre.tdata [39], 
	\kme_cceip1_ob_out_pre.tdata [38], \kme_cceip1_ob_out_pre.tdata [37], 
	\kme_cceip1_ob_out_pre.tdata [36], \kme_cceip1_ob_out_pre.tdata [35], 
	\kme_cceip1_ob_out_pre.tdata [34], \kme_cceip1_ob_out_pre.tdata [33], 
	\kme_cceip1_ob_out_pre.tdata [32], \kme_cceip1_ob_out_pre.tdata [31], 
	\kme_cceip1_ob_out_pre.tdata [30], \kme_cceip1_ob_out_pre.tdata [29], 
	\kme_cceip1_ob_out_pre.tdata [28], \kme_cceip1_ob_out_pre.tdata [27], 
	\kme_cceip1_ob_out_pre.tdata [26], \kme_cceip1_ob_out_pre.tdata [25], 
	\kme_cceip1_ob_out_pre.tdata [24], \kme_cceip1_ob_out_pre.tdata [23], 
	\kme_cceip1_ob_out_pre.tdata [22], \kme_cceip1_ob_out_pre.tdata [21], 
	\kme_cceip1_ob_out_pre.tdata [20], \kme_cceip1_ob_out_pre.tdata [19], 
	\kme_cceip1_ob_out_pre.tdata [18], \kme_cceip1_ob_out_pre.tdata [17], 
	\kme_cceip1_ob_out_pre.tdata [16], \kme_cceip1_ob_out_pre.tdata [15], 
	\kme_cceip1_ob_out_pre.tdata [14], \kme_cceip1_ob_out_pre.tdata [13], 
	\kme_cceip1_ob_out_pre.tdata [12], \kme_cceip1_ob_out_pre.tdata [11], 
	\kme_cceip1_ob_out_pre.tdata [10], \kme_cceip1_ob_out_pre.tdata [9], 
	\kme_cceip1_ob_out_pre.tdata [8], \kme_cceip1_ob_out_pre.tdata [7], 
	\kme_cceip1_ob_out_pre.tdata [6], \kme_cceip1_ob_out_pre.tdata [5], 
	\kme_cceip1_ob_out_pre.tdata [4], \kme_cceip1_ob_out_pre.tdata [3], 
	\kme_cceip1_ob_out_pre.tdata [2], \kme_cceip1_ob_out_pre.tdata [1], 
	\kme_cceip1_ob_out_pre.tdata [0]} ), .kme_cceip1_ob_in( {
	\kme_cceip1_ob_in.tready } ), .kme_cceip2_ob_out_pre( {
	\kme_cceip2_ob_out_pre.tvalid , \kme_cceip2_ob_out_pre.tlast , 
	\kme_cceip2_ob_out_pre.tid [0], \kme_cceip2_ob_out_pre.tstrb [7], 
	\kme_cceip2_ob_out_pre.tstrb [6], \kme_cceip2_ob_out_pre.tstrb [5], 
	\kme_cceip2_ob_out_pre.tstrb [4], \kme_cceip2_ob_out_pre.tstrb [3], 
	\kme_cceip2_ob_out_pre.tstrb [2], \kme_cceip2_ob_out_pre.tstrb [1], 
	\kme_cceip2_ob_out_pre.tstrb [0], \kme_cceip2_ob_out_pre.tuser [7], 
	\kme_cceip2_ob_out_pre.tuser [6], \kme_cceip2_ob_out_pre.tuser [5], 
	\kme_cceip2_ob_out_pre.tuser [4], \kme_cceip2_ob_out_pre.tuser [3], 
	\kme_cceip2_ob_out_pre.tuser [2], \kme_cceip2_ob_out_pre.tuser [1], 
	\kme_cceip2_ob_out_pre.tuser [0], \kme_cceip2_ob_out_pre.tdata [63], 
	\kme_cceip2_ob_out_pre.tdata [62], \kme_cceip2_ob_out_pre.tdata [61], 
	\kme_cceip2_ob_out_pre.tdata [60], \kme_cceip2_ob_out_pre.tdata [59], 
	\kme_cceip2_ob_out_pre.tdata [58], \kme_cceip2_ob_out_pre.tdata [57], 
	\kme_cceip2_ob_out_pre.tdata [56], \kme_cceip2_ob_out_pre.tdata [55], 
	\kme_cceip2_ob_out_pre.tdata [54], \kme_cceip2_ob_out_pre.tdata [53], 
	\kme_cceip2_ob_out_pre.tdata [52], \kme_cceip2_ob_out_pre.tdata [51], 
	\kme_cceip2_ob_out_pre.tdata [50], \kme_cceip2_ob_out_pre.tdata [49], 
	\kme_cceip2_ob_out_pre.tdata [48], \kme_cceip2_ob_out_pre.tdata [47], 
	\kme_cceip2_ob_out_pre.tdata [46], \kme_cceip2_ob_out_pre.tdata [45], 
	\kme_cceip2_ob_out_pre.tdata [44], \kme_cceip2_ob_out_pre.tdata [43], 
	\kme_cceip2_ob_out_pre.tdata [42], \kme_cceip2_ob_out_pre.tdata [41], 
	\kme_cceip2_ob_out_pre.tdata [40], \kme_cceip2_ob_out_pre.tdata [39], 
	\kme_cceip2_ob_out_pre.tdata [38], \kme_cceip2_ob_out_pre.tdata [37], 
	\kme_cceip2_ob_out_pre.tdata [36], \kme_cceip2_ob_out_pre.tdata [35], 
	\kme_cceip2_ob_out_pre.tdata [34], \kme_cceip2_ob_out_pre.tdata [33], 
	\kme_cceip2_ob_out_pre.tdata [32], \kme_cceip2_ob_out_pre.tdata [31], 
	\kme_cceip2_ob_out_pre.tdata [30], \kme_cceip2_ob_out_pre.tdata [29], 
	\kme_cceip2_ob_out_pre.tdata [28], \kme_cceip2_ob_out_pre.tdata [27], 
	\kme_cceip2_ob_out_pre.tdata [26], \kme_cceip2_ob_out_pre.tdata [25], 
	\kme_cceip2_ob_out_pre.tdata [24], \kme_cceip2_ob_out_pre.tdata [23], 
	\kme_cceip2_ob_out_pre.tdata [22], \kme_cceip2_ob_out_pre.tdata [21], 
	\kme_cceip2_ob_out_pre.tdata [20], \kme_cceip2_ob_out_pre.tdata [19], 
	\kme_cceip2_ob_out_pre.tdata [18], \kme_cceip2_ob_out_pre.tdata [17], 
	\kme_cceip2_ob_out_pre.tdata [16], \kme_cceip2_ob_out_pre.tdata [15], 
	\kme_cceip2_ob_out_pre.tdata [14], \kme_cceip2_ob_out_pre.tdata [13], 
	\kme_cceip2_ob_out_pre.tdata [12], \kme_cceip2_ob_out_pre.tdata [11], 
	\kme_cceip2_ob_out_pre.tdata [10], \kme_cceip2_ob_out_pre.tdata [9], 
	\kme_cceip2_ob_out_pre.tdata [8], \kme_cceip2_ob_out_pre.tdata [7], 
	\kme_cceip2_ob_out_pre.tdata [6], \kme_cceip2_ob_out_pre.tdata [5], 
	\kme_cceip2_ob_out_pre.tdata [4], \kme_cceip2_ob_out_pre.tdata [3], 
	\kme_cceip2_ob_out_pre.tdata [2], \kme_cceip2_ob_out_pre.tdata [1], 
	\kme_cceip2_ob_out_pre.tdata [0]} ), .kme_cceip2_ob_in( {
	\kme_cceip2_ob_in.tready } ), .kme_cceip3_ob_out_pre( {
	\kme_cceip3_ob_out_pre.tvalid , \kme_cceip3_ob_out_pre.tlast , 
	\kme_cceip3_ob_out_pre.tid [0], \kme_cceip3_ob_out_pre.tstrb [7], 
	\kme_cceip3_ob_out_pre.tstrb [6], \kme_cceip3_ob_out_pre.tstrb [5], 
	\kme_cceip3_ob_out_pre.tstrb [4], \kme_cceip3_ob_out_pre.tstrb [3], 
	\kme_cceip3_ob_out_pre.tstrb [2], \kme_cceip3_ob_out_pre.tstrb [1], 
	\kme_cceip3_ob_out_pre.tstrb [0], \kme_cceip3_ob_out_pre.tuser [7], 
	\kme_cceip3_ob_out_pre.tuser [6], \kme_cceip3_ob_out_pre.tuser [5], 
	\kme_cceip3_ob_out_pre.tuser [4], \kme_cceip3_ob_out_pre.tuser [3], 
	\kme_cceip3_ob_out_pre.tuser [2], \kme_cceip3_ob_out_pre.tuser [1], 
	\kme_cceip3_ob_out_pre.tuser [0], \kme_cceip3_ob_out_pre.tdata [63], 
	\kme_cceip3_ob_out_pre.tdata [62], \kme_cceip3_ob_out_pre.tdata [61], 
	\kme_cceip3_ob_out_pre.tdata [60], \kme_cceip3_ob_out_pre.tdata [59], 
	\kme_cceip3_ob_out_pre.tdata [58], \kme_cceip3_ob_out_pre.tdata [57], 
	\kme_cceip3_ob_out_pre.tdata [56], \kme_cceip3_ob_out_pre.tdata [55], 
	\kme_cceip3_ob_out_pre.tdata [54], \kme_cceip3_ob_out_pre.tdata [53], 
	\kme_cceip3_ob_out_pre.tdata [52], \kme_cceip3_ob_out_pre.tdata [51], 
	\kme_cceip3_ob_out_pre.tdata [50], \kme_cceip3_ob_out_pre.tdata [49], 
	\kme_cceip3_ob_out_pre.tdata [48], \kme_cceip3_ob_out_pre.tdata [47], 
	\kme_cceip3_ob_out_pre.tdata [46], \kme_cceip3_ob_out_pre.tdata [45], 
	\kme_cceip3_ob_out_pre.tdata [44], \kme_cceip3_ob_out_pre.tdata [43], 
	\kme_cceip3_ob_out_pre.tdata [42], \kme_cceip3_ob_out_pre.tdata [41], 
	\kme_cceip3_ob_out_pre.tdata [40], \kme_cceip3_ob_out_pre.tdata [39], 
	\kme_cceip3_ob_out_pre.tdata [38], \kme_cceip3_ob_out_pre.tdata [37], 
	\kme_cceip3_ob_out_pre.tdata [36], \kme_cceip3_ob_out_pre.tdata [35], 
	\kme_cceip3_ob_out_pre.tdata [34], \kme_cceip3_ob_out_pre.tdata [33], 
	\kme_cceip3_ob_out_pre.tdata [32], \kme_cceip3_ob_out_pre.tdata [31], 
	\kme_cceip3_ob_out_pre.tdata [30], \kme_cceip3_ob_out_pre.tdata [29], 
	\kme_cceip3_ob_out_pre.tdata [28], \kme_cceip3_ob_out_pre.tdata [27], 
	\kme_cceip3_ob_out_pre.tdata [26], \kme_cceip3_ob_out_pre.tdata [25], 
	\kme_cceip3_ob_out_pre.tdata [24], \kme_cceip3_ob_out_pre.tdata [23], 
	\kme_cceip3_ob_out_pre.tdata [22], \kme_cceip3_ob_out_pre.tdata [21], 
	\kme_cceip3_ob_out_pre.tdata [20], \kme_cceip3_ob_out_pre.tdata [19], 
	\kme_cceip3_ob_out_pre.tdata [18], \kme_cceip3_ob_out_pre.tdata [17], 
	\kme_cceip3_ob_out_pre.tdata [16], \kme_cceip3_ob_out_pre.tdata [15], 
	\kme_cceip3_ob_out_pre.tdata [14], \kme_cceip3_ob_out_pre.tdata [13], 
	\kme_cceip3_ob_out_pre.tdata [12], \kme_cceip3_ob_out_pre.tdata [11], 
	\kme_cceip3_ob_out_pre.tdata [10], \kme_cceip3_ob_out_pre.tdata [9], 
	\kme_cceip3_ob_out_pre.tdata [8], \kme_cceip3_ob_out_pre.tdata [7], 
	\kme_cceip3_ob_out_pre.tdata [6], \kme_cceip3_ob_out_pre.tdata [5], 
	\kme_cceip3_ob_out_pre.tdata [4], \kme_cceip3_ob_out_pre.tdata [3], 
	\kme_cceip3_ob_out_pre.tdata [2], \kme_cceip3_ob_out_pre.tdata [1], 
	\kme_cceip3_ob_out_pre.tdata [0]} ), .kme_cceip3_ob_in( {
	\kme_cceip3_ob_in.tready } ), .kme_cddip0_ob_out_pre( {
	\kme_cddip0_ob_out_pre.tvalid , \kme_cddip0_ob_out_pre.tlast , 
	\kme_cddip0_ob_out_pre.tid [0], \kme_cddip0_ob_out_pre.tstrb [7], 
	\kme_cddip0_ob_out_pre.tstrb [6], \kme_cddip0_ob_out_pre.tstrb [5], 
	\kme_cddip0_ob_out_pre.tstrb [4], \kme_cddip0_ob_out_pre.tstrb [3], 
	\kme_cddip0_ob_out_pre.tstrb [2], \kme_cddip0_ob_out_pre.tstrb [1], 
	\kme_cddip0_ob_out_pre.tstrb [0], \kme_cddip0_ob_out_pre.tuser [7], 
	\kme_cddip0_ob_out_pre.tuser [6], \kme_cddip0_ob_out_pre.tuser [5], 
	\kme_cddip0_ob_out_pre.tuser [4], \kme_cddip0_ob_out_pre.tuser [3], 
	\kme_cddip0_ob_out_pre.tuser [2], \kme_cddip0_ob_out_pre.tuser [1], 
	\kme_cddip0_ob_out_pre.tuser [0], \kme_cddip0_ob_out_pre.tdata [63], 
	\kme_cddip0_ob_out_pre.tdata [62], \kme_cddip0_ob_out_pre.tdata [61], 
	\kme_cddip0_ob_out_pre.tdata [60], \kme_cddip0_ob_out_pre.tdata [59], 
	\kme_cddip0_ob_out_pre.tdata [58], \kme_cddip0_ob_out_pre.tdata [57], 
	\kme_cddip0_ob_out_pre.tdata [56], \kme_cddip0_ob_out_pre.tdata [55], 
	\kme_cddip0_ob_out_pre.tdata [54], \kme_cddip0_ob_out_pre.tdata [53], 
	\kme_cddip0_ob_out_pre.tdata [52], \kme_cddip0_ob_out_pre.tdata [51], 
	\kme_cddip0_ob_out_pre.tdata [50], \kme_cddip0_ob_out_pre.tdata [49], 
	\kme_cddip0_ob_out_pre.tdata [48], \kme_cddip0_ob_out_pre.tdata [47], 
	\kme_cddip0_ob_out_pre.tdata [46], \kme_cddip0_ob_out_pre.tdata [45], 
	\kme_cddip0_ob_out_pre.tdata [44], \kme_cddip0_ob_out_pre.tdata [43], 
	\kme_cddip0_ob_out_pre.tdata [42], \kme_cddip0_ob_out_pre.tdata [41], 
	\kme_cddip0_ob_out_pre.tdata [40], \kme_cddip0_ob_out_pre.tdata [39], 
	\kme_cddip0_ob_out_pre.tdata [38], \kme_cddip0_ob_out_pre.tdata [37], 
	\kme_cddip0_ob_out_pre.tdata [36], \kme_cddip0_ob_out_pre.tdata [35], 
	\kme_cddip0_ob_out_pre.tdata [34], \kme_cddip0_ob_out_pre.tdata [33], 
	\kme_cddip0_ob_out_pre.tdata [32], \kme_cddip0_ob_out_pre.tdata [31], 
	\kme_cddip0_ob_out_pre.tdata [30], \kme_cddip0_ob_out_pre.tdata [29], 
	\kme_cddip0_ob_out_pre.tdata [28], \kme_cddip0_ob_out_pre.tdata [27], 
	\kme_cddip0_ob_out_pre.tdata [26], \kme_cddip0_ob_out_pre.tdata [25], 
	\kme_cddip0_ob_out_pre.tdata [24], \kme_cddip0_ob_out_pre.tdata [23], 
	\kme_cddip0_ob_out_pre.tdata [22], \kme_cddip0_ob_out_pre.tdata [21], 
	\kme_cddip0_ob_out_pre.tdata [20], \kme_cddip0_ob_out_pre.tdata [19], 
	\kme_cddip0_ob_out_pre.tdata [18], \kme_cddip0_ob_out_pre.tdata [17], 
	\kme_cddip0_ob_out_pre.tdata [16], \kme_cddip0_ob_out_pre.tdata [15], 
	\kme_cddip0_ob_out_pre.tdata [14], \kme_cddip0_ob_out_pre.tdata [13], 
	\kme_cddip0_ob_out_pre.tdata [12], \kme_cddip0_ob_out_pre.tdata [11], 
	\kme_cddip0_ob_out_pre.tdata [10], \kme_cddip0_ob_out_pre.tdata [9], 
	\kme_cddip0_ob_out_pre.tdata [8], \kme_cddip0_ob_out_pre.tdata [7], 
	\kme_cddip0_ob_out_pre.tdata [6], \kme_cddip0_ob_out_pre.tdata [5], 
	\kme_cddip0_ob_out_pre.tdata [4], \kme_cddip0_ob_out_pre.tdata [3], 
	\kme_cddip0_ob_out_pre.tdata [2], \kme_cddip0_ob_out_pre.tdata [1], 
	\kme_cddip0_ob_out_pre.tdata [0]} ), .kme_cddip0_ob_in( {
	\kme_cddip0_ob_in.tready } ), .kme_cddip1_ob_out_pre( {
	\kme_cddip1_ob_out_pre.tvalid , \kme_cddip1_ob_out_pre.tlast , 
	\kme_cddip1_ob_out_pre.tid [0], \kme_cddip1_ob_out_pre.tstrb [7], 
	\kme_cddip1_ob_out_pre.tstrb [6], \kme_cddip1_ob_out_pre.tstrb [5], 
	\kme_cddip1_ob_out_pre.tstrb [4], \kme_cddip1_ob_out_pre.tstrb [3], 
	\kme_cddip1_ob_out_pre.tstrb [2], \kme_cddip1_ob_out_pre.tstrb [1], 
	\kme_cddip1_ob_out_pre.tstrb [0], \kme_cddip1_ob_out_pre.tuser [7], 
	\kme_cddip1_ob_out_pre.tuser [6], \kme_cddip1_ob_out_pre.tuser [5], 
	\kme_cddip1_ob_out_pre.tuser [4], \kme_cddip1_ob_out_pre.tuser [3], 
	\kme_cddip1_ob_out_pre.tuser [2], \kme_cddip1_ob_out_pre.tuser [1], 
	\kme_cddip1_ob_out_pre.tuser [0], \kme_cddip1_ob_out_pre.tdata [63], 
	\kme_cddip1_ob_out_pre.tdata [62], \kme_cddip1_ob_out_pre.tdata [61], 
	\kme_cddip1_ob_out_pre.tdata [60], \kme_cddip1_ob_out_pre.tdata [59], 
	\kme_cddip1_ob_out_pre.tdata [58], \kme_cddip1_ob_out_pre.tdata [57], 
	\kme_cddip1_ob_out_pre.tdata [56], \kme_cddip1_ob_out_pre.tdata [55], 
	\kme_cddip1_ob_out_pre.tdata [54], \kme_cddip1_ob_out_pre.tdata [53], 
	\kme_cddip1_ob_out_pre.tdata [52], \kme_cddip1_ob_out_pre.tdata [51], 
	\kme_cddip1_ob_out_pre.tdata [50], \kme_cddip1_ob_out_pre.tdata [49], 
	\kme_cddip1_ob_out_pre.tdata [48], \kme_cddip1_ob_out_pre.tdata [47], 
	\kme_cddip1_ob_out_pre.tdata [46], \kme_cddip1_ob_out_pre.tdata [45], 
	\kme_cddip1_ob_out_pre.tdata [44], \kme_cddip1_ob_out_pre.tdata [43], 
	\kme_cddip1_ob_out_pre.tdata [42], \kme_cddip1_ob_out_pre.tdata [41], 
	\kme_cddip1_ob_out_pre.tdata [40], \kme_cddip1_ob_out_pre.tdata [39], 
	\kme_cddip1_ob_out_pre.tdata [38], \kme_cddip1_ob_out_pre.tdata [37], 
	\kme_cddip1_ob_out_pre.tdata [36], \kme_cddip1_ob_out_pre.tdata [35], 
	\kme_cddip1_ob_out_pre.tdata [34], \kme_cddip1_ob_out_pre.tdata [33], 
	\kme_cddip1_ob_out_pre.tdata [32], \kme_cddip1_ob_out_pre.tdata [31], 
	\kme_cddip1_ob_out_pre.tdata [30], \kme_cddip1_ob_out_pre.tdata [29], 
	\kme_cddip1_ob_out_pre.tdata [28], \kme_cddip1_ob_out_pre.tdata [27], 
	\kme_cddip1_ob_out_pre.tdata [26], \kme_cddip1_ob_out_pre.tdata [25], 
	\kme_cddip1_ob_out_pre.tdata [24], \kme_cddip1_ob_out_pre.tdata [23], 
	\kme_cddip1_ob_out_pre.tdata [22], \kme_cddip1_ob_out_pre.tdata [21], 
	\kme_cddip1_ob_out_pre.tdata [20], \kme_cddip1_ob_out_pre.tdata [19], 
	\kme_cddip1_ob_out_pre.tdata [18], \kme_cddip1_ob_out_pre.tdata [17], 
	\kme_cddip1_ob_out_pre.tdata [16], \kme_cddip1_ob_out_pre.tdata [15], 
	\kme_cddip1_ob_out_pre.tdata [14], \kme_cddip1_ob_out_pre.tdata [13], 
	\kme_cddip1_ob_out_pre.tdata [12], \kme_cddip1_ob_out_pre.tdata [11], 
	\kme_cddip1_ob_out_pre.tdata [10], \kme_cddip1_ob_out_pre.tdata [9], 
	\kme_cddip1_ob_out_pre.tdata [8], \kme_cddip1_ob_out_pre.tdata [7], 
	\kme_cddip1_ob_out_pre.tdata [6], \kme_cddip1_ob_out_pre.tdata [5], 
	\kme_cddip1_ob_out_pre.tdata [4], \kme_cddip1_ob_out_pre.tdata [3], 
	\kme_cddip1_ob_out_pre.tdata [2], \kme_cddip1_ob_out_pre.tdata [1], 
	\kme_cddip1_ob_out_pre.tdata [0]} ), .kme_cddip1_ob_in( {
	\kme_cddip1_ob_in.tready } ), .kme_cddip2_ob_out_pre( {
	\kme_cddip2_ob_out_pre.tvalid , \kme_cddip2_ob_out_pre.tlast , 
	\kme_cddip2_ob_out_pre.tid [0], \kme_cddip2_ob_out_pre.tstrb [7], 
	\kme_cddip2_ob_out_pre.tstrb [6], \kme_cddip2_ob_out_pre.tstrb [5], 
	\kme_cddip2_ob_out_pre.tstrb [4], \kme_cddip2_ob_out_pre.tstrb [3], 
	\kme_cddip2_ob_out_pre.tstrb [2], \kme_cddip2_ob_out_pre.tstrb [1], 
	\kme_cddip2_ob_out_pre.tstrb [0], \kme_cddip2_ob_out_pre.tuser [7], 
	\kme_cddip2_ob_out_pre.tuser [6], \kme_cddip2_ob_out_pre.tuser [5], 
	\kme_cddip2_ob_out_pre.tuser [4], \kme_cddip2_ob_out_pre.tuser [3], 
	\kme_cddip2_ob_out_pre.tuser [2], \kme_cddip2_ob_out_pre.tuser [1], 
	\kme_cddip2_ob_out_pre.tuser [0], \kme_cddip2_ob_out_pre.tdata [63], 
	\kme_cddip2_ob_out_pre.tdata [62], \kme_cddip2_ob_out_pre.tdata [61], 
	\kme_cddip2_ob_out_pre.tdata [60], \kme_cddip2_ob_out_pre.tdata [59], 
	\kme_cddip2_ob_out_pre.tdata [58], \kme_cddip2_ob_out_pre.tdata [57], 
	\kme_cddip2_ob_out_pre.tdata [56], \kme_cddip2_ob_out_pre.tdata [55], 
	\kme_cddip2_ob_out_pre.tdata [54], \kme_cddip2_ob_out_pre.tdata [53], 
	\kme_cddip2_ob_out_pre.tdata [52], \kme_cddip2_ob_out_pre.tdata [51], 
	\kme_cddip2_ob_out_pre.tdata [50], \kme_cddip2_ob_out_pre.tdata [49], 
	\kme_cddip2_ob_out_pre.tdata [48], \kme_cddip2_ob_out_pre.tdata [47], 
	\kme_cddip2_ob_out_pre.tdata [46], \kme_cddip2_ob_out_pre.tdata [45], 
	\kme_cddip2_ob_out_pre.tdata [44], \kme_cddip2_ob_out_pre.tdata [43], 
	\kme_cddip2_ob_out_pre.tdata [42], \kme_cddip2_ob_out_pre.tdata [41], 
	\kme_cddip2_ob_out_pre.tdata [40], \kme_cddip2_ob_out_pre.tdata [39], 
	\kme_cddip2_ob_out_pre.tdata [38], \kme_cddip2_ob_out_pre.tdata [37], 
	\kme_cddip2_ob_out_pre.tdata [36], \kme_cddip2_ob_out_pre.tdata [35], 
	\kme_cddip2_ob_out_pre.tdata [34], \kme_cddip2_ob_out_pre.tdata [33], 
	\kme_cddip2_ob_out_pre.tdata [32], \kme_cddip2_ob_out_pre.tdata [31], 
	\kme_cddip2_ob_out_pre.tdata [30], \kme_cddip2_ob_out_pre.tdata [29], 
	\kme_cddip2_ob_out_pre.tdata [28], \kme_cddip2_ob_out_pre.tdata [27], 
	\kme_cddip2_ob_out_pre.tdata [26], \kme_cddip2_ob_out_pre.tdata [25], 
	\kme_cddip2_ob_out_pre.tdata [24], \kme_cddip2_ob_out_pre.tdata [23], 
	\kme_cddip2_ob_out_pre.tdata [22], \kme_cddip2_ob_out_pre.tdata [21], 
	\kme_cddip2_ob_out_pre.tdata [20], \kme_cddip2_ob_out_pre.tdata [19], 
	\kme_cddip2_ob_out_pre.tdata [18], \kme_cddip2_ob_out_pre.tdata [17], 
	\kme_cddip2_ob_out_pre.tdata [16], \kme_cddip2_ob_out_pre.tdata [15], 
	\kme_cddip2_ob_out_pre.tdata [14], \kme_cddip2_ob_out_pre.tdata [13], 
	\kme_cddip2_ob_out_pre.tdata [12], \kme_cddip2_ob_out_pre.tdata [11], 
	\kme_cddip2_ob_out_pre.tdata [10], \kme_cddip2_ob_out_pre.tdata [9], 
	\kme_cddip2_ob_out_pre.tdata [8], \kme_cddip2_ob_out_pre.tdata [7], 
	\kme_cddip2_ob_out_pre.tdata [6], \kme_cddip2_ob_out_pre.tdata [5], 
	\kme_cddip2_ob_out_pre.tdata [4], \kme_cddip2_ob_out_pre.tdata [3], 
	\kme_cddip2_ob_out_pre.tdata [2], \kme_cddip2_ob_out_pre.tdata [1], 
	\kme_cddip2_ob_out_pre.tdata [0]} ), .kme_cddip2_ob_in( {
	\kme_cddip2_ob_in.tready } ), .kme_cddip3_ob_out_pre( {
	\kme_cddip3_ob_out_pre.tvalid , \kme_cddip3_ob_out_pre.tlast , 
	\kme_cddip3_ob_out_pre.tid [0], \kme_cddip3_ob_out_pre.tstrb [7], 
	\kme_cddip3_ob_out_pre.tstrb [6], \kme_cddip3_ob_out_pre.tstrb [5], 
	\kme_cddip3_ob_out_pre.tstrb [4], \kme_cddip3_ob_out_pre.tstrb [3], 
	\kme_cddip3_ob_out_pre.tstrb [2], \kme_cddip3_ob_out_pre.tstrb [1], 
	\kme_cddip3_ob_out_pre.tstrb [0], \kme_cddip3_ob_out_pre.tuser [7], 
	\kme_cddip3_ob_out_pre.tuser [6], \kme_cddip3_ob_out_pre.tuser [5], 
	\kme_cddip3_ob_out_pre.tuser [4], \kme_cddip3_ob_out_pre.tuser [3], 
	\kme_cddip3_ob_out_pre.tuser [2], \kme_cddip3_ob_out_pre.tuser [1], 
	\kme_cddip3_ob_out_pre.tuser [0], \kme_cddip3_ob_out_pre.tdata [63], 
	\kme_cddip3_ob_out_pre.tdata [62], \kme_cddip3_ob_out_pre.tdata [61], 
	\kme_cddip3_ob_out_pre.tdata [60], \kme_cddip3_ob_out_pre.tdata [59], 
	\kme_cddip3_ob_out_pre.tdata [58], \kme_cddip3_ob_out_pre.tdata [57], 
	\kme_cddip3_ob_out_pre.tdata [56], \kme_cddip3_ob_out_pre.tdata [55], 
	\kme_cddip3_ob_out_pre.tdata [54], \kme_cddip3_ob_out_pre.tdata [53], 
	\kme_cddip3_ob_out_pre.tdata [52], \kme_cddip3_ob_out_pre.tdata [51], 
	\kme_cddip3_ob_out_pre.tdata [50], \kme_cddip3_ob_out_pre.tdata [49], 
	\kme_cddip3_ob_out_pre.tdata [48], \kme_cddip3_ob_out_pre.tdata [47], 
	\kme_cddip3_ob_out_pre.tdata [46], \kme_cddip3_ob_out_pre.tdata [45], 
	\kme_cddip3_ob_out_pre.tdata [44], \kme_cddip3_ob_out_pre.tdata [43], 
	\kme_cddip3_ob_out_pre.tdata [42], \kme_cddip3_ob_out_pre.tdata [41], 
	\kme_cddip3_ob_out_pre.tdata [40], \kme_cddip3_ob_out_pre.tdata [39], 
	\kme_cddip3_ob_out_pre.tdata [38], \kme_cddip3_ob_out_pre.tdata [37], 
	\kme_cddip3_ob_out_pre.tdata [36], \kme_cddip3_ob_out_pre.tdata [35], 
	\kme_cddip3_ob_out_pre.tdata [34], \kme_cddip3_ob_out_pre.tdata [33], 
	\kme_cddip3_ob_out_pre.tdata [32], \kme_cddip3_ob_out_pre.tdata [31], 
	\kme_cddip3_ob_out_pre.tdata [30], \kme_cddip3_ob_out_pre.tdata [29], 
	\kme_cddip3_ob_out_pre.tdata [28], \kme_cddip3_ob_out_pre.tdata [27], 
	\kme_cddip3_ob_out_pre.tdata [26], \kme_cddip3_ob_out_pre.tdata [25], 
	\kme_cddip3_ob_out_pre.tdata [24], \kme_cddip3_ob_out_pre.tdata [23], 
	\kme_cddip3_ob_out_pre.tdata [22], \kme_cddip3_ob_out_pre.tdata [21], 
	\kme_cddip3_ob_out_pre.tdata [20], \kme_cddip3_ob_out_pre.tdata [19], 
	\kme_cddip3_ob_out_pre.tdata [18], \kme_cddip3_ob_out_pre.tdata [17], 
	\kme_cddip3_ob_out_pre.tdata [16], \kme_cddip3_ob_out_pre.tdata [15], 
	\kme_cddip3_ob_out_pre.tdata [14], \kme_cddip3_ob_out_pre.tdata [13], 
	\kme_cddip3_ob_out_pre.tdata [12], \kme_cddip3_ob_out_pre.tdata [11], 
	\kme_cddip3_ob_out_pre.tdata [10], \kme_cddip3_ob_out_pre.tdata [9], 
	\kme_cddip3_ob_out_pre.tdata [8], \kme_cddip3_ob_out_pre.tdata [7], 
	\kme_cddip3_ob_out_pre.tdata [6], \kme_cddip3_ob_out_pre.tdata [5], 
	\kme_cddip3_ob_out_pre.tdata [4], \kme_cddip3_ob_out_pre.tdata [3], 
	\kme_cddip3_ob_out_pre.tdata [2], \kme_cddip3_ob_out_pre.tdata [1], 
	\kme_cddip3_ob_out_pre.tdata [0]} ), .kme_cddip3_ob_in( {
	\kme_cddip3_ob_in.tready } ), ckv_rd, ckv_addr, kim_rd, kim_addr, 
	cceip_encrypt_bimc_osync, cceip_encrypt_bimc_odat, cceip_encrypt_mbe, 
	cceip_validate_bimc_osync, cceip_validate_bimc_odat, 
	cceip_validate_mbe, cddip_decrypt_bimc_osync, 
	cddip_decrypt_bimc_odat, cddip_decrypt_mbe, axi_bimc_osync, 
	axi_bimc_odat, axi_mbe, seed0_invalidate, seed1_invalidate, 
	set_txc_bp_int, set_gcm_tag_fail_int, set_key_tlv_miscmp_int, 
	set_tlv_bip2_error_int, set_rsm_is_backpressuring, .idle_components( {
	\idle_components.r.part0 [31], \idle_components.r.part0 [30], 
	\idle_components.r.part0 [29], \idle_components.r.part0 [28], 
	\idle_components.r.part0 [27], \idle_components.r.part0 [26], 
	\idle_components.r.part0 [25], \idle_components.r.part0 [24], 
	\idle_components.r.part0 [23], \idle_components.r.part0 [22], 
	\idle_components.r.part0 [21], \idle_components.r.part0 [20], 
	\idle_components.r.part0 [19], \idle_components.r.part0 [18], 
	\idle_components.r.part0 [17], \idle_components.r.part0 [16], 
	\idle_components.r.part0 [15], \idle_components.r.part0 [14], 
	\idle_components.r.part0 [13], \idle_components.r.part0 [12], 
	\idle_components.r.part0 [11], \idle_components.r.part0 [10], 
	\idle_components.r.part0 [9], \idle_components.r.part0 [8], 
	\idle_components.r.part0 [7], \idle_components.r.part0 [6], 
	\idle_components.r.part0 [5], \idle_components.r.part0 [4], 
	\idle_components.r.part0 [3], \idle_components.r.part0 [2], 
	\idle_components.r.part0 [1], \idle_components.r.part0 [0]} ), 
	.sa_snapshot( {\sa_snapshot[31].r.part1[31] , 
	\sa_snapshot[31].r.part1[30] , \sa_snapshot[31].r.part1[29] , 
	\sa_snapshot[31].r.part1[28] , \sa_snapshot[31].r.part1[27] , 
	\sa_snapshot[31].r.part1[26] , \sa_snapshot[31].r.part1[25] , 
	\sa_snapshot[31].r.part1[24] , \sa_snapshot[31].r.part1[23] , 
	\sa_snapshot[31].r.part1[22] , \sa_snapshot[31].r.part1[21] , 
	\sa_snapshot[31].r.part1[20] , \sa_snapshot[31].r.part1[19] , 
	\sa_snapshot[31].r.part1[18] , \sa_snapshot[31].r.part1[17] , 
	\sa_snapshot[31].r.part1[16] , \sa_snapshot[31].r.part1[15] , 
	\sa_snapshot[31].r.part1[14] , \sa_snapshot[31].r.part1[13] , 
	\sa_snapshot[31].r.part1[12] , \sa_snapshot[31].r.part1[11] , 
	\sa_snapshot[31].r.part1[10] , \sa_snapshot[31].r.part1[9] , 
	\sa_snapshot[31].r.part1[8] , \sa_snapshot[31].r.part1[7] , 
	\sa_snapshot[31].r.part1[6] , \sa_snapshot[31].r.part1[5] , 
	\sa_snapshot[31].r.part1[4] , \sa_snapshot[31].r.part1[3] , 
	\sa_snapshot[31].r.part1[2] , \sa_snapshot[31].r.part1[1] , 
	\sa_snapshot[31].r.part1[0] , \sa_snapshot[31].r.part0[31] , 
	\sa_snapshot[31].r.part0[30] , \sa_snapshot[31].r.part0[29] , 
	\sa_snapshot[31].r.part0[28] , \sa_snapshot[31].r.part0[27] , 
	\sa_snapshot[31].r.part0[26] , \sa_snapshot[31].r.part0[25] , 
	\sa_snapshot[31].r.part0[24] , \sa_snapshot[31].r.part0[23] , 
	\sa_snapshot[31].r.part0[22] , \sa_snapshot[31].r.part0[21] , 
	\sa_snapshot[31].r.part0[20] , \sa_snapshot[31].r.part0[19] , 
	\sa_snapshot[31].r.part0[18] , \sa_snapshot[31].r.part0[17] , 
	\sa_snapshot[31].r.part0[16] , \sa_snapshot[31].r.part0[15] , 
	\sa_snapshot[31].r.part0[14] , \sa_snapshot[31].r.part0[13] , 
	\sa_snapshot[31].r.part0[12] , \sa_snapshot[31].r.part0[11] , 
	\sa_snapshot[31].r.part0[10] , \sa_snapshot[31].r.part0[9] , 
	\sa_snapshot[31].r.part0[8] , \sa_snapshot[31].r.part0[7] , 
	\sa_snapshot[31].r.part0[6] , \sa_snapshot[31].r.part0[5] , 
	\sa_snapshot[31].r.part0[4] , \sa_snapshot[31].r.part0[3] , 
	\sa_snapshot[31].r.part0[2] , \sa_snapshot[31].r.part0[1] , 
	\sa_snapshot[31].r.part0[0] , \sa_snapshot[30].r.part1[31] , 
	\sa_snapshot[30].r.part1[30] , \sa_snapshot[30].r.part1[29] , 
	\sa_snapshot[30].r.part1[28] , \sa_snapshot[30].r.part1[27] , 
	\sa_snapshot[30].r.part1[26] , \sa_snapshot[30].r.part1[25] , 
	\sa_snapshot[30].r.part1[24] , \sa_snapshot[30].r.part1[23] , 
	\sa_snapshot[30].r.part1[22] , \sa_snapshot[30].r.part1[21] , 
	\sa_snapshot[30].r.part1[20] , \sa_snapshot[30].r.part1[19] , 
	\sa_snapshot[30].r.part1[18] , \sa_snapshot[30].r.part1[17] , 
	\sa_snapshot[30].r.part1[16] , \sa_snapshot[30].r.part1[15] , 
	\sa_snapshot[30].r.part1[14] , \sa_snapshot[30].r.part1[13] , 
	\sa_snapshot[30].r.part1[12] , \sa_snapshot[30].r.part1[11] , 
	\sa_snapshot[30].r.part1[10] , \sa_snapshot[30].r.part1[9] , 
	\sa_snapshot[30].r.part1[8] , \sa_snapshot[30].r.part1[7] , 
	\sa_snapshot[30].r.part1[6] , \sa_snapshot[30].r.part1[5] , 
	\sa_snapshot[30].r.part1[4] , \sa_snapshot[30].r.part1[3] , 
	\sa_snapshot[30].r.part1[2] , \sa_snapshot[30].r.part1[1] , 
	\sa_snapshot[30].r.part1[0] , \sa_snapshot[30].r.part0[31] , 
	\sa_snapshot[30].r.part0[30] , \sa_snapshot[30].r.part0[29] , 
	\sa_snapshot[30].r.part0[28] , \sa_snapshot[30].r.part0[27] , 
	\sa_snapshot[30].r.part0[26] , \sa_snapshot[30].r.part0[25] , 
	\sa_snapshot[30].r.part0[24] , \sa_snapshot[30].r.part0[23] , 
	\sa_snapshot[30].r.part0[22] , \sa_snapshot[30].r.part0[21] , 
	\sa_snapshot[30].r.part0[20] , \sa_snapshot[30].r.part0[19] , 
	\sa_snapshot[30].r.part0[18] , \sa_snapshot[30].r.part0[17] , 
	\sa_snapshot[30].r.part0[16] , \sa_snapshot[30].r.part0[15] , 
	\sa_snapshot[30].r.part0[14] , \sa_snapshot[30].r.part0[13] , 
	\sa_snapshot[30].r.part0[12] , \sa_snapshot[30].r.part0[11] , 
	\sa_snapshot[30].r.part0[10] , \sa_snapshot[30].r.part0[9] , 
	\sa_snapshot[30].r.part0[8] , \sa_snapshot[30].r.part0[7] , 
	\sa_snapshot[30].r.part0[6] , \sa_snapshot[30].r.part0[5] , 
	\sa_snapshot[30].r.part0[4] , \sa_snapshot[30].r.part0[3] , 
	\sa_snapshot[30].r.part0[2] , \sa_snapshot[30].r.part0[1] , 
	\sa_snapshot[30].r.part0[0] , \sa_snapshot[29].r.part1[31] , 
	\sa_snapshot[29].r.part1[30] , \sa_snapshot[29].r.part1[29] , 
	\sa_snapshot[29].r.part1[28] , \sa_snapshot[29].r.part1[27] , 
	\sa_snapshot[29].r.part1[26] , \sa_snapshot[29].r.part1[25] , 
	\sa_snapshot[29].r.part1[24] , \sa_snapshot[29].r.part1[23] , 
	\sa_snapshot[29].r.part1[22] , \sa_snapshot[29].r.part1[21] , 
	\sa_snapshot[29].r.part1[20] , \sa_snapshot[29].r.part1[19] , 
	\sa_snapshot[29].r.part1[18] , \sa_snapshot[29].r.part1[17] , 
	\sa_snapshot[29].r.part1[16] , \sa_snapshot[29].r.part1[15] , 
	\sa_snapshot[29].r.part1[14] , \sa_snapshot[29].r.part1[13] , 
	\sa_snapshot[29].r.part1[12] , \sa_snapshot[29].r.part1[11] , 
	\sa_snapshot[29].r.part1[10] , \sa_snapshot[29].r.part1[9] , 
	\sa_snapshot[29].r.part1[8] , \sa_snapshot[29].r.part1[7] , 
	\sa_snapshot[29].r.part1[6] , \sa_snapshot[29].r.part1[5] , 
	\sa_snapshot[29].r.part1[4] , \sa_snapshot[29].r.part1[3] , 
	\sa_snapshot[29].r.part1[2] , \sa_snapshot[29].r.part1[1] , 
	\sa_snapshot[29].r.part1[0] , \sa_snapshot[29].r.part0[31] , 
	\sa_snapshot[29].r.part0[30] , \sa_snapshot[29].r.part0[29] , 
	\sa_snapshot[29].r.part0[28] , \sa_snapshot[29].r.part0[27] , 
	\sa_snapshot[29].r.part0[26] , \sa_snapshot[29].r.part0[25] , 
	\sa_snapshot[29].r.part0[24] , \sa_snapshot[29].r.part0[23] , 
	\sa_snapshot[29].r.part0[22] , \sa_snapshot[29].r.part0[21] , 
	\sa_snapshot[29].r.part0[20] , \sa_snapshot[29].r.part0[19] , 
	\sa_snapshot[29].r.part0[18] , \sa_snapshot[29].r.part0[17] , 
	\sa_snapshot[29].r.part0[16] , \sa_snapshot[29].r.part0[15] , 
	\sa_snapshot[29].r.part0[14] , \sa_snapshot[29].r.part0[13] , 
	\sa_snapshot[29].r.part0[12] , \sa_snapshot[29].r.part0[11] , 
	\sa_snapshot[29].r.part0[10] , \sa_snapshot[29].r.part0[9] , 
	\sa_snapshot[29].r.part0[8] , \sa_snapshot[29].r.part0[7] , 
	\sa_snapshot[29].r.part0[6] , \sa_snapshot[29].r.part0[5] , 
	\sa_snapshot[29].r.part0[4] , \sa_snapshot[29].r.part0[3] , 
	\sa_snapshot[29].r.part0[2] , \sa_snapshot[29].r.part0[1] , 
	\sa_snapshot[29].r.part0[0] , \sa_snapshot[28].r.part1[31] , 
	\sa_snapshot[28].r.part1[30] , \sa_snapshot[28].r.part1[29] , 
	\sa_snapshot[28].r.part1[28] , \sa_snapshot[28].r.part1[27] , 
	\sa_snapshot[28].r.part1[26] , \sa_snapshot[28].r.part1[25] , 
	\sa_snapshot[28].r.part1[24] , \sa_snapshot[28].r.part1[23] , 
	\sa_snapshot[28].r.part1[22] , \sa_snapshot[28].r.part1[21] , 
	\sa_snapshot[28].r.part1[20] , \sa_snapshot[28].r.part1[19] , 
	\sa_snapshot[28].r.part1[18] , \sa_snapshot[28].r.part1[17] , 
	\sa_snapshot[28].r.part1[16] , \sa_snapshot[28].r.part1[15] , 
	\sa_snapshot[28].r.part1[14] , \sa_snapshot[28].r.part1[13] , 
	\sa_snapshot[28].r.part1[12] , \sa_snapshot[28].r.part1[11] , 
	\sa_snapshot[28].r.part1[10] , \sa_snapshot[28].r.part1[9] , 
	\sa_snapshot[28].r.part1[8] , \sa_snapshot[28].r.part1[7] , 
	\sa_snapshot[28].r.part1[6] , \sa_snapshot[28].r.part1[5] , 
	\sa_snapshot[28].r.part1[4] , \sa_snapshot[28].r.part1[3] , 
	\sa_snapshot[28].r.part1[2] , \sa_snapshot[28].r.part1[1] , 
	\sa_snapshot[28].r.part1[0] , \sa_snapshot[28].r.part0[31] , 
	\sa_snapshot[28].r.part0[30] , \sa_snapshot[28].r.part0[29] , 
	\sa_snapshot[28].r.part0[28] , \sa_snapshot[28].r.part0[27] , 
	\sa_snapshot[28].r.part0[26] , \sa_snapshot[28].r.part0[25] , 
	\sa_snapshot[28].r.part0[24] , \sa_snapshot[28].r.part0[23] , 
	\sa_snapshot[28].r.part0[22] , \sa_snapshot[28].r.part0[21] , 
	\sa_snapshot[28].r.part0[20] , \sa_snapshot[28].r.part0[19] , 
	\sa_snapshot[28].r.part0[18] , \sa_snapshot[28].r.part0[17] , 
	\sa_snapshot[28].r.part0[16] , \sa_snapshot[28].r.part0[15] , 
	\sa_snapshot[28].r.part0[14] , \sa_snapshot[28].r.part0[13] , 
	\sa_snapshot[28].r.part0[12] , \sa_snapshot[28].r.part0[11] , 
	\sa_snapshot[28].r.part0[10] , \sa_snapshot[28].r.part0[9] , 
	\sa_snapshot[28].r.part0[8] , \sa_snapshot[28].r.part0[7] , 
	\sa_snapshot[28].r.part0[6] , \sa_snapshot[28].r.part0[5] , 
	\sa_snapshot[28].r.part0[4] , \sa_snapshot[28].r.part0[3] , 
	\sa_snapshot[28].r.part0[2] , \sa_snapshot[28].r.part0[1] , 
	\sa_snapshot[28].r.part0[0] , \sa_snapshot[27].r.part1[31] , 
	\sa_snapshot[27].r.part1[30] , \sa_snapshot[27].r.part1[29] , 
	\sa_snapshot[27].r.part1[28] , \sa_snapshot[27].r.part1[27] , 
	\sa_snapshot[27].r.part1[26] , \sa_snapshot[27].r.part1[25] , 
	\sa_snapshot[27].r.part1[24] , \sa_snapshot[27].r.part1[23] , 
	\sa_snapshot[27].r.part1[22] , \sa_snapshot[27].r.part1[21] , 
	\sa_snapshot[27].r.part1[20] , \sa_snapshot[27].r.part1[19] , 
	\sa_snapshot[27].r.part1[18] , \sa_snapshot[27].r.part1[17] , 
	\sa_snapshot[27].r.part1[16] , \sa_snapshot[27].r.part1[15] , 
	\sa_snapshot[27].r.part1[14] , \sa_snapshot[27].r.part1[13] , 
	\sa_snapshot[27].r.part1[12] , \sa_snapshot[27].r.part1[11] , 
	\sa_snapshot[27].r.part1[10] , \sa_snapshot[27].r.part1[9] , 
	\sa_snapshot[27].r.part1[8] , \sa_snapshot[27].r.part1[7] , 
	\sa_snapshot[27].r.part1[6] , \sa_snapshot[27].r.part1[5] , 
	\sa_snapshot[27].r.part1[4] , \sa_snapshot[27].r.part1[3] , 
	\sa_snapshot[27].r.part1[2] , \sa_snapshot[27].r.part1[1] , 
	\sa_snapshot[27].r.part1[0] , \sa_snapshot[27].r.part0[31] , 
	\sa_snapshot[27].r.part0[30] , \sa_snapshot[27].r.part0[29] , 
	\sa_snapshot[27].r.part0[28] , \sa_snapshot[27].r.part0[27] , 
	\sa_snapshot[27].r.part0[26] , \sa_snapshot[27].r.part0[25] , 
	\sa_snapshot[27].r.part0[24] , \sa_snapshot[27].r.part0[23] , 
	\sa_snapshot[27].r.part0[22] , \sa_snapshot[27].r.part0[21] , 
	\sa_snapshot[27].r.part0[20] , \sa_snapshot[27].r.part0[19] , 
	\sa_snapshot[27].r.part0[18] , \sa_snapshot[27].r.part0[17] , 
	\sa_snapshot[27].r.part0[16] , \sa_snapshot[27].r.part0[15] , 
	\sa_snapshot[27].r.part0[14] , \sa_snapshot[27].r.part0[13] , 
	\sa_snapshot[27].r.part0[12] , \sa_snapshot[27].r.part0[11] , 
	\sa_snapshot[27].r.part0[10] , \sa_snapshot[27].r.part0[9] , 
	\sa_snapshot[27].r.part0[8] , \sa_snapshot[27].r.part0[7] , 
	\sa_snapshot[27].r.part0[6] , \sa_snapshot[27].r.part0[5] , 
	\sa_snapshot[27].r.part0[4] , \sa_snapshot[27].r.part0[3] , 
	\sa_snapshot[27].r.part0[2] , \sa_snapshot[27].r.part0[1] , 
	\sa_snapshot[27].r.part0[0] , \sa_snapshot[26].r.part1[31] , 
	\sa_snapshot[26].r.part1[30] , \sa_snapshot[26].r.part1[29] , 
	\sa_snapshot[26].r.part1[28] , \sa_snapshot[26].r.part1[27] , 
	\sa_snapshot[26].r.part1[26] , \sa_snapshot[26].r.part1[25] , 
	\sa_snapshot[26].r.part1[24] , \sa_snapshot[26].r.part1[23] , 
	\sa_snapshot[26].r.part1[22] , \sa_snapshot[26].r.part1[21] , 
	\sa_snapshot[26].r.part1[20] , \sa_snapshot[26].r.part1[19] , 
	\sa_snapshot[26].r.part1[18] , \sa_snapshot[26].r.part1[17] , 
	\sa_snapshot[26].r.part1[16] , \sa_snapshot[26].r.part1[15] , 
	\sa_snapshot[26].r.part1[14] , \sa_snapshot[26].r.part1[13] , 
	\sa_snapshot[26].r.part1[12] , \sa_snapshot[26].r.part1[11] , 
	\sa_snapshot[26].r.part1[10] , \sa_snapshot[26].r.part1[9] , 
	\sa_snapshot[26].r.part1[8] , \sa_snapshot[26].r.part1[7] , 
	\sa_snapshot[26].r.part1[6] , \sa_snapshot[26].r.part1[5] , 
	\sa_snapshot[26].r.part1[4] , \sa_snapshot[26].r.part1[3] , 
	\sa_snapshot[26].r.part1[2] , \sa_snapshot[26].r.part1[1] , 
	\sa_snapshot[26].r.part1[0] , \sa_snapshot[26].r.part0[31] , 
	\sa_snapshot[26].r.part0[30] , \sa_snapshot[26].r.part0[29] , 
	\sa_snapshot[26].r.part0[28] , \sa_snapshot[26].r.part0[27] , 
	\sa_snapshot[26].r.part0[26] , \sa_snapshot[26].r.part0[25] , 
	\sa_snapshot[26].r.part0[24] , \sa_snapshot[26].r.part0[23] , 
	\sa_snapshot[26].r.part0[22] , \sa_snapshot[26].r.part0[21] , 
	\sa_snapshot[26].r.part0[20] , \sa_snapshot[26].r.part0[19] , 
	\sa_snapshot[26].r.part0[18] , \sa_snapshot[26].r.part0[17] , 
	\sa_snapshot[26].r.part0[16] , \sa_snapshot[26].r.part0[15] , 
	\sa_snapshot[26].r.part0[14] , \sa_snapshot[26].r.part0[13] , 
	\sa_snapshot[26].r.part0[12] , \sa_snapshot[26].r.part0[11] , 
	\sa_snapshot[26].r.part0[10] , \sa_snapshot[26].r.part0[9] , 
	\sa_snapshot[26].r.part0[8] , \sa_snapshot[26].r.part0[7] , 
	\sa_snapshot[26].r.part0[6] , \sa_snapshot[26].r.part0[5] , 
	\sa_snapshot[26].r.part0[4] , \sa_snapshot[26].r.part0[3] , 
	\sa_snapshot[26].r.part0[2] , \sa_snapshot[26].r.part0[1] , 
	\sa_snapshot[26].r.part0[0] , \sa_snapshot[25].r.part1[31] , 
	\sa_snapshot[25].r.part1[30] , \sa_snapshot[25].r.part1[29] , 
	\sa_snapshot[25].r.part1[28] , \sa_snapshot[25].r.part1[27] , 
	\sa_snapshot[25].r.part1[26] , \sa_snapshot[25].r.part1[25] , 
	\sa_snapshot[25].r.part1[24] , \sa_snapshot[25].r.part1[23] , 
	\sa_snapshot[25].r.part1[22] , \sa_snapshot[25].r.part1[21] , 
	\sa_snapshot[25].r.part1[20] , \sa_snapshot[25].r.part1[19] , 
	\sa_snapshot[25].r.part1[18] , \sa_snapshot[25].r.part1[17] , 
	\sa_snapshot[25].r.part1[16] , \sa_snapshot[25].r.part1[15] , 
	\sa_snapshot[25].r.part1[14] , \sa_snapshot[25].r.part1[13] , 
	\sa_snapshot[25].r.part1[12] , \sa_snapshot[25].r.part1[11] , 
	\sa_snapshot[25].r.part1[10] , \sa_snapshot[25].r.part1[9] , 
	\sa_snapshot[25].r.part1[8] , \sa_snapshot[25].r.part1[7] , 
	\sa_snapshot[25].r.part1[6] , \sa_snapshot[25].r.part1[5] , 
	\sa_snapshot[25].r.part1[4] , \sa_snapshot[25].r.part1[3] , 
	\sa_snapshot[25].r.part1[2] , \sa_snapshot[25].r.part1[1] , 
	\sa_snapshot[25].r.part1[0] , \sa_snapshot[25].r.part0[31] , 
	\sa_snapshot[25].r.part0[30] , \sa_snapshot[25].r.part0[29] , 
	\sa_snapshot[25].r.part0[28] , \sa_snapshot[25].r.part0[27] , 
	\sa_snapshot[25].r.part0[26] , \sa_snapshot[25].r.part0[25] , 
	\sa_snapshot[25].r.part0[24] , \sa_snapshot[25].r.part0[23] , 
	\sa_snapshot[25].r.part0[22] , \sa_snapshot[25].r.part0[21] , 
	\sa_snapshot[25].r.part0[20] , \sa_snapshot[25].r.part0[19] , 
	\sa_snapshot[25].r.part0[18] , \sa_snapshot[25].r.part0[17] , 
	\sa_snapshot[25].r.part0[16] , \sa_snapshot[25].r.part0[15] , 
	\sa_snapshot[25].r.part0[14] , \sa_snapshot[25].r.part0[13] , 
	\sa_snapshot[25].r.part0[12] , \sa_snapshot[25].r.part0[11] , 
	\sa_snapshot[25].r.part0[10] , \sa_snapshot[25].r.part0[9] , 
	\sa_snapshot[25].r.part0[8] , \sa_snapshot[25].r.part0[7] , 
	\sa_snapshot[25].r.part0[6] , \sa_snapshot[25].r.part0[5] , 
	\sa_snapshot[25].r.part0[4] , \sa_snapshot[25].r.part0[3] , 
	\sa_snapshot[25].r.part0[2] , \sa_snapshot[25].r.part0[1] , 
	\sa_snapshot[25].r.part0[0] , \sa_snapshot[24].r.part1[31] , 
	\sa_snapshot[24].r.part1[30] , \sa_snapshot[24].r.part1[29] , 
	\sa_snapshot[24].r.part1[28] , \sa_snapshot[24].r.part1[27] , 
	\sa_snapshot[24].r.part1[26] , \sa_snapshot[24].r.part1[25] , 
	\sa_snapshot[24].r.part1[24] , \sa_snapshot[24].r.part1[23] , 
	\sa_snapshot[24].r.part1[22] , \sa_snapshot[24].r.part1[21] , 
	\sa_snapshot[24].r.part1[20] , \sa_snapshot[24].r.part1[19] , 
	\sa_snapshot[24].r.part1[18] , \sa_snapshot[24].r.part1[17] , 
	\sa_snapshot[24].r.part1[16] , \sa_snapshot[24].r.part1[15] , 
	\sa_snapshot[24].r.part1[14] , \sa_snapshot[24].r.part1[13] , 
	\sa_snapshot[24].r.part1[12] , \sa_snapshot[24].r.part1[11] , 
	\sa_snapshot[24].r.part1[10] , \sa_snapshot[24].r.part1[9] , 
	\sa_snapshot[24].r.part1[8] , \sa_snapshot[24].r.part1[7] , 
	\sa_snapshot[24].r.part1[6] , \sa_snapshot[24].r.part1[5] , 
	\sa_snapshot[24].r.part1[4] , \sa_snapshot[24].r.part1[3] , 
	\sa_snapshot[24].r.part1[2] , \sa_snapshot[24].r.part1[1] , 
	\sa_snapshot[24].r.part1[0] , \sa_snapshot[24].r.part0[31] , 
	\sa_snapshot[24].r.part0[30] , \sa_snapshot[24].r.part0[29] , 
	\sa_snapshot[24].r.part0[28] , \sa_snapshot[24].r.part0[27] , 
	\sa_snapshot[24].r.part0[26] , \sa_snapshot[24].r.part0[25] , 
	\sa_snapshot[24].r.part0[24] , \sa_snapshot[24].r.part0[23] , 
	\sa_snapshot[24].r.part0[22] , \sa_snapshot[24].r.part0[21] , 
	\sa_snapshot[24].r.part0[20] , \sa_snapshot[24].r.part0[19] , 
	\sa_snapshot[24].r.part0[18] , \sa_snapshot[24].r.part0[17] , 
	\sa_snapshot[24].r.part0[16] , \sa_snapshot[24].r.part0[15] , 
	\sa_snapshot[24].r.part0[14] , \sa_snapshot[24].r.part0[13] , 
	\sa_snapshot[24].r.part0[12] , \sa_snapshot[24].r.part0[11] , 
	\sa_snapshot[24].r.part0[10] , \sa_snapshot[24].r.part0[9] , 
	\sa_snapshot[24].r.part0[8] , \sa_snapshot[24].r.part0[7] , 
	\sa_snapshot[24].r.part0[6] , \sa_snapshot[24].r.part0[5] , 
	\sa_snapshot[24].r.part0[4] , \sa_snapshot[24].r.part0[3] , 
	\sa_snapshot[24].r.part0[2] , \sa_snapshot[24].r.part0[1] , 
	\sa_snapshot[24].r.part0[0] , \sa_snapshot[23].r.part1[31] , 
	\sa_snapshot[23].r.part1[30] , \sa_snapshot[23].r.part1[29] , 
	\sa_snapshot[23].r.part1[28] , \sa_snapshot[23].r.part1[27] , 
	\sa_snapshot[23].r.part1[26] , \sa_snapshot[23].r.part1[25] , 
	\sa_snapshot[23].r.part1[24] , \sa_snapshot[23].r.part1[23] , 
	\sa_snapshot[23].r.part1[22] , \sa_snapshot[23].r.part1[21] , 
	\sa_snapshot[23].r.part1[20] , \sa_snapshot[23].r.part1[19] , 
	\sa_snapshot[23].r.part1[18] , \sa_snapshot[23].r.part1[17] , 
	\sa_snapshot[23].r.part1[16] , \sa_snapshot[23].r.part1[15] , 
	\sa_snapshot[23].r.part1[14] , \sa_snapshot[23].r.part1[13] , 
	\sa_snapshot[23].r.part1[12] , \sa_snapshot[23].r.part1[11] , 
	\sa_snapshot[23].r.part1[10] , \sa_snapshot[23].r.part1[9] , 
	\sa_snapshot[23].r.part1[8] , \sa_snapshot[23].r.part1[7] , 
	\sa_snapshot[23].r.part1[6] , \sa_snapshot[23].r.part1[5] , 
	\sa_snapshot[23].r.part1[4] , \sa_snapshot[23].r.part1[3] , 
	\sa_snapshot[23].r.part1[2] , \sa_snapshot[23].r.part1[1] , 
	\sa_snapshot[23].r.part1[0] , \sa_snapshot[23].r.part0[31] , 
	\sa_snapshot[23].r.part0[30] , \sa_snapshot[23].r.part0[29] , 
	\sa_snapshot[23].r.part0[28] , \sa_snapshot[23].r.part0[27] , 
	\sa_snapshot[23].r.part0[26] , \sa_snapshot[23].r.part0[25] , 
	\sa_snapshot[23].r.part0[24] , \sa_snapshot[23].r.part0[23] , 
	\sa_snapshot[23].r.part0[22] , \sa_snapshot[23].r.part0[21] , 
	\sa_snapshot[23].r.part0[20] , \sa_snapshot[23].r.part0[19] , 
	\sa_snapshot[23].r.part0[18] , \sa_snapshot[23].r.part0[17] , 
	\sa_snapshot[23].r.part0[16] , \sa_snapshot[23].r.part0[15] , 
	\sa_snapshot[23].r.part0[14] , \sa_snapshot[23].r.part0[13] , 
	\sa_snapshot[23].r.part0[12] , \sa_snapshot[23].r.part0[11] , 
	\sa_snapshot[23].r.part0[10] , \sa_snapshot[23].r.part0[9] , 
	\sa_snapshot[23].r.part0[8] , \sa_snapshot[23].r.part0[7] , 
	\sa_snapshot[23].r.part0[6] , \sa_snapshot[23].r.part0[5] , 
	\sa_snapshot[23].r.part0[4] , \sa_snapshot[23].r.part0[3] , 
	\sa_snapshot[23].r.part0[2] , \sa_snapshot[23].r.part0[1] , 
	\sa_snapshot[23].r.part0[0] , \sa_snapshot[22].r.part1[31] , 
	\sa_snapshot[22].r.part1[30] , \sa_snapshot[22].r.part1[29] , 
	\sa_snapshot[22].r.part1[28] , \sa_snapshot[22].r.part1[27] , 
	\sa_snapshot[22].r.part1[26] , \sa_snapshot[22].r.part1[25] , 
	\sa_snapshot[22].r.part1[24] , \sa_snapshot[22].r.part1[23] , 
	\sa_snapshot[22].r.part1[22] , \sa_snapshot[22].r.part1[21] , 
	\sa_snapshot[22].r.part1[20] , \sa_snapshot[22].r.part1[19] , 
	\sa_snapshot[22].r.part1[18] , \sa_snapshot[22].r.part1[17] , 
	\sa_snapshot[22].r.part1[16] , \sa_snapshot[22].r.part1[15] , 
	\sa_snapshot[22].r.part1[14] , \sa_snapshot[22].r.part1[13] , 
	\sa_snapshot[22].r.part1[12] , \sa_snapshot[22].r.part1[11] , 
	\sa_snapshot[22].r.part1[10] , \sa_snapshot[22].r.part1[9] , 
	\sa_snapshot[22].r.part1[8] , \sa_snapshot[22].r.part1[7] , 
	\sa_snapshot[22].r.part1[6] , \sa_snapshot[22].r.part1[5] , 
	\sa_snapshot[22].r.part1[4] , \sa_snapshot[22].r.part1[3] , 
	\sa_snapshot[22].r.part1[2] , \sa_snapshot[22].r.part1[1] , 
	\sa_snapshot[22].r.part1[0] , \sa_snapshot[22].r.part0[31] , 
	\sa_snapshot[22].r.part0[30] , \sa_snapshot[22].r.part0[29] , 
	\sa_snapshot[22].r.part0[28] , \sa_snapshot[22].r.part0[27] , 
	\sa_snapshot[22].r.part0[26] , \sa_snapshot[22].r.part0[25] , 
	\sa_snapshot[22].r.part0[24] , \sa_snapshot[22].r.part0[23] , 
	\sa_snapshot[22].r.part0[22] , \sa_snapshot[22].r.part0[21] , 
	\sa_snapshot[22].r.part0[20] , \sa_snapshot[22].r.part0[19] , 
	\sa_snapshot[22].r.part0[18] , \sa_snapshot[22].r.part0[17] , 
	\sa_snapshot[22].r.part0[16] , \sa_snapshot[22].r.part0[15] , 
	\sa_snapshot[22].r.part0[14] , \sa_snapshot[22].r.part0[13] , 
	\sa_snapshot[22].r.part0[12] , \sa_snapshot[22].r.part0[11] , 
	\sa_snapshot[22].r.part0[10] , \sa_snapshot[22].r.part0[9] , 
	\sa_snapshot[22].r.part0[8] , \sa_snapshot[22].r.part0[7] , 
	\sa_snapshot[22].r.part0[6] , \sa_snapshot[22].r.part0[5] , 
	\sa_snapshot[22].r.part0[4] , \sa_snapshot[22].r.part0[3] , 
	\sa_snapshot[22].r.part0[2] , \sa_snapshot[22].r.part0[1] , 
	\sa_snapshot[22].r.part0[0] , \sa_snapshot[21].r.part1[31] , 
	\sa_snapshot[21].r.part1[30] , \sa_snapshot[21].r.part1[29] , 
	\sa_snapshot[21].r.part1[28] , \sa_snapshot[21].r.part1[27] , 
	\sa_snapshot[21].r.part1[26] , \sa_snapshot[21].r.part1[25] , 
	\sa_snapshot[21].r.part1[24] , \sa_snapshot[21].r.part1[23] , 
	\sa_snapshot[21].r.part1[22] , \sa_snapshot[21].r.part1[21] , 
	\sa_snapshot[21].r.part1[20] , \sa_snapshot[21].r.part1[19] , 
	\sa_snapshot[21].r.part1[18] , \sa_snapshot[21].r.part1[17] , 
	\sa_snapshot[21].r.part1[16] , \sa_snapshot[21].r.part1[15] , 
	\sa_snapshot[21].r.part1[14] , \sa_snapshot[21].r.part1[13] , 
	\sa_snapshot[21].r.part1[12] , \sa_snapshot[21].r.part1[11] , 
	\sa_snapshot[21].r.part1[10] , \sa_snapshot[21].r.part1[9] , 
	\sa_snapshot[21].r.part1[8] , \sa_snapshot[21].r.part1[7] , 
	\sa_snapshot[21].r.part1[6] , \sa_snapshot[21].r.part1[5] , 
	\sa_snapshot[21].r.part1[4] , \sa_snapshot[21].r.part1[3] , 
	\sa_snapshot[21].r.part1[2] , \sa_snapshot[21].r.part1[1] , 
	\sa_snapshot[21].r.part1[0] , \sa_snapshot[21].r.part0[31] , 
	\sa_snapshot[21].r.part0[30] , \sa_snapshot[21].r.part0[29] , 
	\sa_snapshot[21].r.part0[28] , \sa_snapshot[21].r.part0[27] , 
	\sa_snapshot[21].r.part0[26] , \sa_snapshot[21].r.part0[25] , 
	\sa_snapshot[21].r.part0[24] , \sa_snapshot[21].r.part0[23] , 
	\sa_snapshot[21].r.part0[22] , \sa_snapshot[21].r.part0[21] , 
	\sa_snapshot[21].r.part0[20] , \sa_snapshot[21].r.part0[19] , 
	\sa_snapshot[21].r.part0[18] , \sa_snapshot[21].r.part0[17] , 
	\sa_snapshot[21].r.part0[16] , \sa_snapshot[21].r.part0[15] , 
	\sa_snapshot[21].r.part0[14] , \sa_snapshot[21].r.part0[13] , 
	\sa_snapshot[21].r.part0[12] , \sa_snapshot[21].r.part0[11] , 
	\sa_snapshot[21].r.part0[10] , \sa_snapshot[21].r.part0[9] , 
	\sa_snapshot[21].r.part0[8] , \sa_snapshot[21].r.part0[7] , 
	\sa_snapshot[21].r.part0[6] , \sa_snapshot[21].r.part0[5] , 
	\sa_snapshot[21].r.part0[4] , \sa_snapshot[21].r.part0[3] , 
	\sa_snapshot[21].r.part0[2] , \sa_snapshot[21].r.part0[1] , 
	\sa_snapshot[21].r.part0[0] , \sa_snapshot[20].r.part1[31] , 
	\sa_snapshot[20].r.part1[30] , \sa_snapshot[20].r.part1[29] , 
	\sa_snapshot[20].r.part1[28] , \sa_snapshot[20].r.part1[27] , 
	\sa_snapshot[20].r.part1[26] , \sa_snapshot[20].r.part1[25] , 
	\sa_snapshot[20].r.part1[24] , \sa_snapshot[20].r.part1[23] , 
	\sa_snapshot[20].r.part1[22] , \sa_snapshot[20].r.part1[21] , 
	\sa_snapshot[20].r.part1[20] , \sa_snapshot[20].r.part1[19] , 
	\sa_snapshot[20].r.part1[18] , \sa_snapshot[20].r.part1[17] , 
	\sa_snapshot[20].r.part1[16] , \sa_snapshot[20].r.part1[15] , 
	\sa_snapshot[20].r.part1[14] , \sa_snapshot[20].r.part1[13] , 
	\sa_snapshot[20].r.part1[12] , \sa_snapshot[20].r.part1[11] , 
	\sa_snapshot[20].r.part1[10] , \sa_snapshot[20].r.part1[9] , 
	\sa_snapshot[20].r.part1[8] , \sa_snapshot[20].r.part1[7] , 
	\sa_snapshot[20].r.part1[6] , \sa_snapshot[20].r.part1[5] , 
	\sa_snapshot[20].r.part1[4] , \sa_snapshot[20].r.part1[3] , 
	\sa_snapshot[20].r.part1[2] , \sa_snapshot[20].r.part1[1] , 
	\sa_snapshot[20].r.part1[0] , \sa_snapshot[20].r.part0[31] , 
	\sa_snapshot[20].r.part0[30] , \sa_snapshot[20].r.part0[29] , 
	\sa_snapshot[20].r.part0[28] , \sa_snapshot[20].r.part0[27] , 
	\sa_snapshot[20].r.part0[26] , \sa_snapshot[20].r.part0[25] , 
	\sa_snapshot[20].r.part0[24] , \sa_snapshot[20].r.part0[23] , 
	\sa_snapshot[20].r.part0[22] , \sa_snapshot[20].r.part0[21] , 
	\sa_snapshot[20].r.part0[20] , \sa_snapshot[20].r.part0[19] , 
	\sa_snapshot[20].r.part0[18] , \sa_snapshot[20].r.part0[17] , 
	\sa_snapshot[20].r.part0[16] , \sa_snapshot[20].r.part0[15] , 
	\sa_snapshot[20].r.part0[14] , \sa_snapshot[20].r.part0[13] , 
	\sa_snapshot[20].r.part0[12] , \sa_snapshot[20].r.part0[11] , 
	\sa_snapshot[20].r.part0[10] , \sa_snapshot[20].r.part0[9] , 
	\sa_snapshot[20].r.part0[8] , \sa_snapshot[20].r.part0[7] , 
	\sa_snapshot[20].r.part0[6] , \sa_snapshot[20].r.part0[5] , 
	\sa_snapshot[20].r.part0[4] , \sa_snapshot[20].r.part0[3] , 
	\sa_snapshot[20].r.part0[2] , \sa_snapshot[20].r.part0[1] , 
	\sa_snapshot[20].r.part0[0] , \sa_snapshot[19].r.part1[31] , 
	\sa_snapshot[19].r.part1[30] , \sa_snapshot[19].r.part1[29] , 
	\sa_snapshot[19].r.part1[28] , \sa_snapshot[19].r.part1[27] , 
	\sa_snapshot[19].r.part1[26] , \sa_snapshot[19].r.part1[25] , 
	\sa_snapshot[19].r.part1[24] , \sa_snapshot[19].r.part1[23] , 
	\sa_snapshot[19].r.part1[22] , \sa_snapshot[19].r.part1[21] , 
	\sa_snapshot[19].r.part1[20] , \sa_snapshot[19].r.part1[19] , 
	\sa_snapshot[19].r.part1[18] , \sa_snapshot[19].r.part1[17] , 
	\sa_snapshot[19].r.part1[16] , \sa_snapshot[19].r.part1[15] , 
	\sa_snapshot[19].r.part1[14] , \sa_snapshot[19].r.part1[13] , 
	\sa_snapshot[19].r.part1[12] , \sa_snapshot[19].r.part1[11] , 
	\sa_snapshot[19].r.part1[10] , \sa_snapshot[19].r.part1[9] , 
	\sa_snapshot[19].r.part1[8] , \sa_snapshot[19].r.part1[7] , 
	\sa_snapshot[19].r.part1[6] , \sa_snapshot[19].r.part1[5] , 
	\sa_snapshot[19].r.part1[4] , \sa_snapshot[19].r.part1[3] , 
	\sa_snapshot[19].r.part1[2] , \sa_snapshot[19].r.part1[1] , 
	\sa_snapshot[19].r.part1[0] , \sa_snapshot[19].r.part0[31] , 
	\sa_snapshot[19].r.part0[30] , \sa_snapshot[19].r.part0[29] , 
	\sa_snapshot[19].r.part0[28] , \sa_snapshot[19].r.part0[27] , 
	\sa_snapshot[19].r.part0[26] , \sa_snapshot[19].r.part0[25] , 
	\sa_snapshot[19].r.part0[24] , \sa_snapshot[19].r.part0[23] , 
	\sa_snapshot[19].r.part0[22] , \sa_snapshot[19].r.part0[21] , 
	\sa_snapshot[19].r.part0[20] , \sa_snapshot[19].r.part0[19] , 
	\sa_snapshot[19].r.part0[18] , \sa_snapshot[19].r.part0[17] , 
	\sa_snapshot[19].r.part0[16] , \sa_snapshot[19].r.part0[15] , 
	\sa_snapshot[19].r.part0[14] , \sa_snapshot[19].r.part0[13] , 
	\sa_snapshot[19].r.part0[12] , \sa_snapshot[19].r.part0[11] , 
	\sa_snapshot[19].r.part0[10] , \sa_snapshot[19].r.part0[9] , 
	\sa_snapshot[19].r.part0[8] , \sa_snapshot[19].r.part0[7] , 
	\sa_snapshot[19].r.part0[6] , \sa_snapshot[19].r.part0[5] , 
	\sa_snapshot[19].r.part0[4] , \sa_snapshot[19].r.part0[3] , 
	\sa_snapshot[19].r.part0[2] , \sa_snapshot[19].r.part0[1] , 
	\sa_snapshot[19].r.part0[0] , \sa_snapshot[18].r.part1[31] , 
	\sa_snapshot[18].r.part1[30] , \sa_snapshot[18].r.part1[29] , 
	\sa_snapshot[18].r.part1[28] , \sa_snapshot[18].r.part1[27] , 
	\sa_snapshot[18].r.part1[26] , \sa_snapshot[18].r.part1[25] , 
	\sa_snapshot[18].r.part1[24] , \sa_snapshot[18].r.part1[23] , 
	\sa_snapshot[18].r.part1[22] , \sa_snapshot[18].r.part1[21] , 
	\sa_snapshot[18].r.part1[20] , \sa_snapshot[18].r.part1[19] , 
	\sa_snapshot[18].r.part1[18] , \sa_snapshot[18].r.part1[17] , 
	\sa_snapshot[18].r.part1[16] , \sa_snapshot[18].r.part1[15] , 
	\sa_snapshot[18].r.part1[14] , \sa_snapshot[18].r.part1[13] , 
	\sa_snapshot[18].r.part1[12] , \sa_snapshot[18].r.part1[11] , 
	\sa_snapshot[18].r.part1[10] , \sa_snapshot[18].r.part1[9] , 
	\sa_snapshot[18].r.part1[8] , \sa_snapshot[18].r.part1[7] , 
	\sa_snapshot[18].r.part1[6] , \sa_snapshot[18].r.part1[5] , 
	\sa_snapshot[18].r.part1[4] , \sa_snapshot[18].r.part1[3] , 
	\sa_snapshot[18].r.part1[2] , \sa_snapshot[18].r.part1[1] , 
	\sa_snapshot[18].r.part1[0] , \sa_snapshot[18].r.part0[31] , 
	\sa_snapshot[18].r.part0[30] , \sa_snapshot[18].r.part0[29] , 
	\sa_snapshot[18].r.part0[28] , \sa_snapshot[18].r.part0[27] , 
	\sa_snapshot[18].r.part0[26] , \sa_snapshot[18].r.part0[25] , 
	\sa_snapshot[18].r.part0[24] , \sa_snapshot[18].r.part0[23] , 
	\sa_snapshot[18].r.part0[22] , \sa_snapshot[18].r.part0[21] , 
	\sa_snapshot[18].r.part0[20] , \sa_snapshot[18].r.part0[19] , 
	\sa_snapshot[18].r.part0[18] , \sa_snapshot[18].r.part0[17] , 
	\sa_snapshot[18].r.part0[16] , \sa_snapshot[18].r.part0[15] , 
	\sa_snapshot[18].r.part0[14] , \sa_snapshot[18].r.part0[13] , 
	\sa_snapshot[18].r.part0[12] , \sa_snapshot[18].r.part0[11] , 
	\sa_snapshot[18].r.part0[10] , \sa_snapshot[18].r.part0[9] , 
	\sa_snapshot[18].r.part0[8] , \sa_snapshot[18].r.part0[7] , 
	\sa_snapshot[18].r.part0[6] , \sa_snapshot[18].r.part0[5] , 
	\sa_snapshot[18].r.part0[4] , \sa_snapshot[18].r.part0[3] , 
	\sa_snapshot[18].r.part0[2] , \sa_snapshot[18].r.part0[1] , 
	\sa_snapshot[18].r.part0[0] , \sa_snapshot[17].r.part1[31] , 
	\sa_snapshot[17].r.part1[30] , \sa_snapshot[17].r.part1[29] , 
	\sa_snapshot[17].r.part1[28] , \sa_snapshot[17].r.part1[27] , 
	\sa_snapshot[17].r.part1[26] , \sa_snapshot[17].r.part1[25] , 
	\sa_snapshot[17].r.part1[24] , \sa_snapshot[17].r.part1[23] , 
	\sa_snapshot[17].r.part1[22] , \sa_snapshot[17].r.part1[21] , 
	\sa_snapshot[17].r.part1[20] , \sa_snapshot[17].r.part1[19] , 
	\sa_snapshot[17].r.part1[18] , \sa_snapshot[17].r.part1[17] , 
	\sa_snapshot[17].r.part1[16] , \sa_snapshot[17].r.part1[15] , 
	\sa_snapshot[17].r.part1[14] , \sa_snapshot[17].r.part1[13] , 
	\sa_snapshot[17].r.part1[12] , \sa_snapshot[17].r.part1[11] , 
	\sa_snapshot[17].r.part1[10] , \sa_snapshot[17].r.part1[9] , 
	\sa_snapshot[17].r.part1[8] , \sa_snapshot[17].r.part1[7] , 
	\sa_snapshot[17].r.part1[6] , \sa_snapshot[17].r.part1[5] , 
	\sa_snapshot[17].r.part1[4] , \sa_snapshot[17].r.part1[3] , 
	\sa_snapshot[17].r.part1[2] , \sa_snapshot[17].r.part1[1] , 
	\sa_snapshot[17].r.part1[0] , \sa_snapshot[17].r.part0[31] , 
	\sa_snapshot[17].r.part0[30] , \sa_snapshot[17].r.part0[29] , 
	\sa_snapshot[17].r.part0[28] , \sa_snapshot[17].r.part0[27] , 
	\sa_snapshot[17].r.part0[26] , \sa_snapshot[17].r.part0[25] , 
	\sa_snapshot[17].r.part0[24] , \sa_snapshot[17].r.part0[23] , 
	\sa_snapshot[17].r.part0[22] , \sa_snapshot[17].r.part0[21] , 
	\sa_snapshot[17].r.part0[20] , \sa_snapshot[17].r.part0[19] , 
	\sa_snapshot[17].r.part0[18] , \sa_snapshot[17].r.part0[17] , 
	\sa_snapshot[17].r.part0[16] , \sa_snapshot[17].r.part0[15] , 
	\sa_snapshot[17].r.part0[14] , \sa_snapshot[17].r.part0[13] , 
	\sa_snapshot[17].r.part0[12] , \sa_snapshot[17].r.part0[11] , 
	\sa_snapshot[17].r.part0[10] , \sa_snapshot[17].r.part0[9] , 
	\sa_snapshot[17].r.part0[8] , \sa_snapshot[17].r.part0[7] , 
	\sa_snapshot[17].r.part0[6] , \sa_snapshot[17].r.part0[5] , 
	\sa_snapshot[17].r.part0[4] , \sa_snapshot[17].r.part0[3] , 
	\sa_snapshot[17].r.part0[2] , \sa_snapshot[17].r.part0[1] , 
	\sa_snapshot[17].r.part0[0] , \sa_snapshot[16].r.part1[31] , 
	\sa_snapshot[16].r.part1[30] , \sa_snapshot[16].r.part1[29] , 
	\sa_snapshot[16].r.part1[28] , \sa_snapshot[16].r.part1[27] , 
	\sa_snapshot[16].r.part1[26] , \sa_snapshot[16].r.part1[25] , 
	\sa_snapshot[16].r.part1[24] , \sa_snapshot[16].r.part1[23] , 
	\sa_snapshot[16].r.part1[22] , \sa_snapshot[16].r.part1[21] , 
	\sa_snapshot[16].r.part1[20] , \sa_snapshot[16].r.part1[19] , 
	\sa_snapshot[16].r.part1[18] , \sa_snapshot[16].r.part1[17] , 
	\sa_snapshot[16].r.part1[16] , \sa_snapshot[16].r.part1[15] , 
	\sa_snapshot[16].r.part1[14] , \sa_snapshot[16].r.part1[13] , 
	\sa_snapshot[16].r.part1[12] , \sa_snapshot[16].r.part1[11] , 
	\sa_snapshot[16].r.part1[10] , \sa_snapshot[16].r.part1[9] , 
	\sa_snapshot[16].r.part1[8] , \sa_snapshot[16].r.part1[7] , 
	\sa_snapshot[16].r.part1[6] , \sa_snapshot[16].r.part1[5] , 
	\sa_snapshot[16].r.part1[4] , \sa_snapshot[16].r.part1[3] , 
	\sa_snapshot[16].r.part1[2] , \sa_snapshot[16].r.part1[1] , 
	\sa_snapshot[16].r.part1[0] , \sa_snapshot[16].r.part0[31] , 
	\sa_snapshot[16].r.part0[30] , \sa_snapshot[16].r.part0[29] , 
	\sa_snapshot[16].r.part0[28] , \sa_snapshot[16].r.part0[27] , 
	\sa_snapshot[16].r.part0[26] , \sa_snapshot[16].r.part0[25] , 
	\sa_snapshot[16].r.part0[24] , \sa_snapshot[16].r.part0[23] , 
	\sa_snapshot[16].r.part0[22] , \sa_snapshot[16].r.part0[21] , 
	\sa_snapshot[16].r.part0[20] , \sa_snapshot[16].r.part0[19] , 
	\sa_snapshot[16].r.part0[18] , \sa_snapshot[16].r.part0[17] , 
	\sa_snapshot[16].r.part0[16] , \sa_snapshot[16].r.part0[15] , 
	\sa_snapshot[16].r.part0[14] , \sa_snapshot[16].r.part0[13] , 
	\sa_snapshot[16].r.part0[12] , \sa_snapshot[16].r.part0[11] , 
	\sa_snapshot[16].r.part0[10] , \sa_snapshot[16].r.part0[9] , 
	\sa_snapshot[16].r.part0[8] , \sa_snapshot[16].r.part0[7] , 
	\sa_snapshot[16].r.part0[6] , \sa_snapshot[16].r.part0[5] , 
	\sa_snapshot[16].r.part0[4] , \sa_snapshot[16].r.part0[3] , 
	\sa_snapshot[16].r.part0[2] , \sa_snapshot[16].r.part0[1] , 
	\sa_snapshot[16].r.part0[0] , \sa_snapshot[15].r.part1[31] , 
	\sa_snapshot[15].r.part1[30] , \sa_snapshot[15].r.part1[29] , 
	\sa_snapshot[15].r.part1[28] , \sa_snapshot[15].r.part1[27] , 
	\sa_snapshot[15].r.part1[26] , \sa_snapshot[15].r.part1[25] , 
	\sa_snapshot[15].r.part1[24] , \sa_snapshot[15].r.part1[23] , 
	\sa_snapshot[15].r.part1[22] , \sa_snapshot[15].r.part1[21] , 
	\sa_snapshot[15].r.part1[20] , \sa_snapshot[15].r.part1[19] , 
	\sa_snapshot[15].r.part1[18] , \sa_snapshot[15].r.part1[17] , 
	\sa_snapshot[15].r.part1[16] , \sa_snapshot[15].r.part1[15] , 
	\sa_snapshot[15].r.part1[14] , \sa_snapshot[15].r.part1[13] , 
	\sa_snapshot[15].r.part1[12] , \sa_snapshot[15].r.part1[11] , 
	\sa_snapshot[15].r.part1[10] , \sa_snapshot[15].r.part1[9] , 
	\sa_snapshot[15].r.part1[8] , \sa_snapshot[15].r.part1[7] , 
	\sa_snapshot[15].r.part1[6] , \sa_snapshot[15].r.part1[5] , 
	\sa_snapshot[15].r.part1[4] , \sa_snapshot[15].r.part1[3] , 
	\sa_snapshot[15].r.part1[2] , \sa_snapshot[15].r.part1[1] , 
	\sa_snapshot[15].r.part1[0] , \sa_snapshot[15].r.part0[31] , 
	\sa_snapshot[15].r.part0[30] , \sa_snapshot[15].r.part0[29] , 
	\sa_snapshot[15].r.part0[28] , \sa_snapshot[15].r.part0[27] , 
	\sa_snapshot[15].r.part0[26] , \sa_snapshot[15].r.part0[25] , 
	\sa_snapshot[15].r.part0[24] , \sa_snapshot[15].r.part0[23] , 
	\sa_snapshot[15].r.part0[22] , \sa_snapshot[15].r.part0[21] , 
	\sa_snapshot[15].r.part0[20] , \sa_snapshot[15].r.part0[19] , 
	\sa_snapshot[15].r.part0[18] , \sa_snapshot[15].r.part0[17] , 
	\sa_snapshot[15].r.part0[16] , \sa_snapshot[15].r.part0[15] , 
	\sa_snapshot[15].r.part0[14] , \sa_snapshot[15].r.part0[13] , 
	\sa_snapshot[15].r.part0[12] , \sa_snapshot[15].r.part0[11] , 
	\sa_snapshot[15].r.part0[10] , \sa_snapshot[15].r.part0[9] , 
	\sa_snapshot[15].r.part0[8] , \sa_snapshot[15].r.part0[7] , 
	\sa_snapshot[15].r.part0[6] , \sa_snapshot[15].r.part0[5] , 
	\sa_snapshot[15].r.part0[4] , \sa_snapshot[15].r.part0[3] , 
	\sa_snapshot[15].r.part0[2] , \sa_snapshot[15].r.part0[1] , 
	\sa_snapshot[15].r.part0[0] , \sa_snapshot[14].r.part1[31] , 
	\sa_snapshot[14].r.part1[30] , \sa_snapshot[14].r.part1[29] , 
	\sa_snapshot[14].r.part1[28] , \sa_snapshot[14].r.part1[27] , 
	\sa_snapshot[14].r.part1[26] , \sa_snapshot[14].r.part1[25] , 
	\sa_snapshot[14].r.part1[24] , \sa_snapshot[14].r.part1[23] , 
	\sa_snapshot[14].r.part1[22] , \sa_snapshot[14].r.part1[21] , 
	\sa_snapshot[14].r.part1[20] , \sa_snapshot[14].r.part1[19] , 
	\sa_snapshot[14].r.part1[18] , \sa_snapshot[14].r.part1[17] , 
	\sa_snapshot[14].r.part1[16] , \sa_snapshot[14].r.part1[15] , 
	\sa_snapshot[14].r.part1[14] , \sa_snapshot[14].r.part1[13] , 
	\sa_snapshot[14].r.part1[12] , \sa_snapshot[14].r.part1[11] , 
	\sa_snapshot[14].r.part1[10] , \sa_snapshot[14].r.part1[9] , 
	\sa_snapshot[14].r.part1[8] , \sa_snapshot[14].r.part1[7] , 
	\sa_snapshot[14].r.part1[6] , \sa_snapshot[14].r.part1[5] , 
	\sa_snapshot[14].r.part1[4] , \sa_snapshot[14].r.part1[3] , 
	\sa_snapshot[14].r.part1[2] , \sa_snapshot[14].r.part1[1] , 
	\sa_snapshot[14].r.part1[0] , \sa_snapshot[14].r.part0[31] , 
	\sa_snapshot[14].r.part0[30] , \sa_snapshot[14].r.part0[29] , 
	\sa_snapshot[14].r.part0[28] , \sa_snapshot[14].r.part0[27] , 
	\sa_snapshot[14].r.part0[26] , \sa_snapshot[14].r.part0[25] , 
	\sa_snapshot[14].r.part0[24] , \sa_snapshot[14].r.part0[23] , 
	\sa_snapshot[14].r.part0[22] , \sa_snapshot[14].r.part0[21] , 
	\sa_snapshot[14].r.part0[20] , \sa_snapshot[14].r.part0[19] , 
	\sa_snapshot[14].r.part0[18] , \sa_snapshot[14].r.part0[17] , 
	\sa_snapshot[14].r.part0[16] , \sa_snapshot[14].r.part0[15] , 
	\sa_snapshot[14].r.part0[14] , \sa_snapshot[14].r.part0[13] , 
	\sa_snapshot[14].r.part0[12] , \sa_snapshot[14].r.part0[11] , 
	\sa_snapshot[14].r.part0[10] , \sa_snapshot[14].r.part0[9] , 
	\sa_snapshot[14].r.part0[8] , \sa_snapshot[14].r.part0[7] , 
	\sa_snapshot[14].r.part0[6] , \sa_snapshot[14].r.part0[5] , 
	\sa_snapshot[14].r.part0[4] , \sa_snapshot[14].r.part0[3] , 
	\sa_snapshot[14].r.part0[2] , \sa_snapshot[14].r.part0[1] , 
	\sa_snapshot[14].r.part0[0] , \sa_snapshot[13].r.part1[31] , 
	\sa_snapshot[13].r.part1[30] , \sa_snapshot[13].r.part1[29] , 
	\sa_snapshot[13].r.part1[28] , \sa_snapshot[13].r.part1[27] , 
	\sa_snapshot[13].r.part1[26] , \sa_snapshot[13].r.part1[25] , 
	\sa_snapshot[13].r.part1[24] , \sa_snapshot[13].r.part1[23] , 
	\sa_snapshot[13].r.part1[22] , \sa_snapshot[13].r.part1[21] , 
	\sa_snapshot[13].r.part1[20] , \sa_snapshot[13].r.part1[19] , 
	\sa_snapshot[13].r.part1[18] , \sa_snapshot[13].r.part1[17] , 
	\sa_snapshot[13].r.part1[16] , \sa_snapshot[13].r.part1[15] , 
	\sa_snapshot[13].r.part1[14] , \sa_snapshot[13].r.part1[13] , 
	\sa_snapshot[13].r.part1[12] , \sa_snapshot[13].r.part1[11] , 
	\sa_snapshot[13].r.part1[10] , \sa_snapshot[13].r.part1[9] , 
	\sa_snapshot[13].r.part1[8] , \sa_snapshot[13].r.part1[7] , 
	\sa_snapshot[13].r.part1[6] , \sa_snapshot[13].r.part1[5] , 
	\sa_snapshot[13].r.part1[4] , \sa_snapshot[13].r.part1[3] , 
	\sa_snapshot[13].r.part1[2] , \sa_snapshot[13].r.part1[1] , 
	\sa_snapshot[13].r.part1[0] , \sa_snapshot[13].r.part0[31] , 
	\sa_snapshot[13].r.part0[30] , \sa_snapshot[13].r.part0[29] , 
	\sa_snapshot[13].r.part0[28] , \sa_snapshot[13].r.part0[27] , 
	\sa_snapshot[13].r.part0[26] , \sa_snapshot[13].r.part0[25] , 
	\sa_snapshot[13].r.part0[24] , \sa_snapshot[13].r.part0[23] , 
	\sa_snapshot[13].r.part0[22] , \sa_snapshot[13].r.part0[21] , 
	\sa_snapshot[13].r.part0[20] , \sa_snapshot[13].r.part0[19] , 
	\sa_snapshot[13].r.part0[18] , \sa_snapshot[13].r.part0[17] , 
	\sa_snapshot[13].r.part0[16] , \sa_snapshot[13].r.part0[15] , 
	\sa_snapshot[13].r.part0[14] , \sa_snapshot[13].r.part0[13] , 
	\sa_snapshot[13].r.part0[12] , \sa_snapshot[13].r.part0[11] , 
	\sa_snapshot[13].r.part0[10] , \sa_snapshot[13].r.part0[9] , 
	\sa_snapshot[13].r.part0[8] , \sa_snapshot[13].r.part0[7] , 
	\sa_snapshot[13].r.part0[6] , \sa_snapshot[13].r.part0[5] , 
	\sa_snapshot[13].r.part0[4] , \sa_snapshot[13].r.part0[3] , 
	\sa_snapshot[13].r.part0[2] , \sa_snapshot[13].r.part0[1] , 
	\sa_snapshot[13].r.part0[0] , \sa_snapshot[12].r.part1[31] , 
	\sa_snapshot[12].r.part1[30] , \sa_snapshot[12].r.part1[29] , 
	\sa_snapshot[12].r.part1[28] , \sa_snapshot[12].r.part1[27] , 
	\sa_snapshot[12].r.part1[26] , \sa_snapshot[12].r.part1[25] , 
	\sa_snapshot[12].r.part1[24] , \sa_snapshot[12].r.part1[23] , 
	\sa_snapshot[12].r.part1[22] , \sa_snapshot[12].r.part1[21] , 
	\sa_snapshot[12].r.part1[20] , \sa_snapshot[12].r.part1[19] , 
	\sa_snapshot[12].r.part1[18] , \sa_snapshot[12].r.part1[17] , 
	\sa_snapshot[12].r.part1[16] , \sa_snapshot[12].r.part1[15] , 
	\sa_snapshot[12].r.part1[14] , \sa_snapshot[12].r.part1[13] , 
	\sa_snapshot[12].r.part1[12] , \sa_snapshot[12].r.part1[11] , 
	\sa_snapshot[12].r.part1[10] , \sa_snapshot[12].r.part1[9] , 
	\sa_snapshot[12].r.part1[8] , \sa_snapshot[12].r.part1[7] , 
	\sa_snapshot[12].r.part1[6] , \sa_snapshot[12].r.part1[5] , 
	\sa_snapshot[12].r.part1[4] , \sa_snapshot[12].r.part1[3] , 
	\sa_snapshot[12].r.part1[2] , \sa_snapshot[12].r.part1[1] , 
	\sa_snapshot[12].r.part1[0] , \sa_snapshot[12].r.part0[31] , 
	\sa_snapshot[12].r.part0[30] , \sa_snapshot[12].r.part0[29] , 
	\sa_snapshot[12].r.part0[28] , \sa_snapshot[12].r.part0[27] , 
	\sa_snapshot[12].r.part0[26] , \sa_snapshot[12].r.part0[25] , 
	\sa_snapshot[12].r.part0[24] , \sa_snapshot[12].r.part0[23] , 
	\sa_snapshot[12].r.part0[22] , \sa_snapshot[12].r.part0[21] , 
	\sa_snapshot[12].r.part0[20] , \sa_snapshot[12].r.part0[19] , 
	\sa_snapshot[12].r.part0[18] , \sa_snapshot[12].r.part0[17] , 
	\sa_snapshot[12].r.part0[16] , \sa_snapshot[12].r.part0[15] , 
	\sa_snapshot[12].r.part0[14] , \sa_snapshot[12].r.part0[13] , 
	\sa_snapshot[12].r.part0[12] , \sa_snapshot[12].r.part0[11] , 
	\sa_snapshot[12].r.part0[10] , \sa_snapshot[12].r.part0[9] , 
	\sa_snapshot[12].r.part0[8] , \sa_snapshot[12].r.part0[7] , 
	\sa_snapshot[12].r.part0[6] , \sa_snapshot[12].r.part0[5] , 
	\sa_snapshot[12].r.part0[4] , \sa_snapshot[12].r.part0[3] , 
	\sa_snapshot[12].r.part0[2] , \sa_snapshot[12].r.part0[1] , 
	\sa_snapshot[12].r.part0[0] , \sa_snapshot[11].r.part1[31] , 
	\sa_snapshot[11].r.part1[30] , \sa_snapshot[11].r.part1[29] , 
	\sa_snapshot[11].r.part1[28] , \sa_snapshot[11].r.part1[27] , 
	\sa_snapshot[11].r.part1[26] , \sa_snapshot[11].r.part1[25] , 
	\sa_snapshot[11].r.part1[24] , \sa_snapshot[11].r.part1[23] , 
	\sa_snapshot[11].r.part1[22] , \sa_snapshot[11].r.part1[21] , 
	\sa_snapshot[11].r.part1[20] , \sa_snapshot[11].r.part1[19] , 
	\sa_snapshot[11].r.part1[18] , \sa_snapshot[11].r.part1[17] , 
	\sa_snapshot[11].r.part1[16] , \sa_snapshot[11].r.part1[15] , 
	\sa_snapshot[11].r.part1[14] , \sa_snapshot[11].r.part1[13] , 
	\sa_snapshot[11].r.part1[12] , \sa_snapshot[11].r.part1[11] , 
	\sa_snapshot[11].r.part1[10] , \sa_snapshot[11].r.part1[9] , 
	\sa_snapshot[11].r.part1[8] , \sa_snapshot[11].r.part1[7] , 
	\sa_snapshot[11].r.part1[6] , \sa_snapshot[11].r.part1[5] , 
	\sa_snapshot[11].r.part1[4] , \sa_snapshot[11].r.part1[3] , 
	\sa_snapshot[11].r.part1[2] , \sa_snapshot[11].r.part1[1] , 
	\sa_snapshot[11].r.part1[0] , \sa_snapshot[11].r.part0[31] , 
	\sa_snapshot[11].r.part0[30] , \sa_snapshot[11].r.part0[29] , 
	\sa_snapshot[11].r.part0[28] , \sa_snapshot[11].r.part0[27] , 
	\sa_snapshot[11].r.part0[26] , \sa_snapshot[11].r.part0[25] , 
	\sa_snapshot[11].r.part0[24] , \sa_snapshot[11].r.part0[23] , 
	\sa_snapshot[11].r.part0[22] , \sa_snapshot[11].r.part0[21] , 
	\sa_snapshot[11].r.part0[20] , \sa_snapshot[11].r.part0[19] , 
	\sa_snapshot[11].r.part0[18] , \sa_snapshot[11].r.part0[17] , 
	\sa_snapshot[11].r.part0[16] , \sa_snapshot[11].r.part0[15] , 
	\sa_snapshot[11].r.part0[14] , \sa_snapshot[11].r.part0[13] , 
	\sa_snapshot[11].r.part0[12] , \sa_snapshot[11].r.part0[11] , 
	\sa_snapshot[11].r.part0[10] , \sa_snapshot[11].r.part0[9] , 
	\sa_snapshot[11].r.part0[8] , \sa_snapshot[11].r.part0[7] , 
	\sa_snapshot[11].r.part0[6] , \sa_snapshot[11].r.part0[5] , 
	\sa_snapshot[11].r.part0[4] , \sa_snapshot[11].r.part0[3] , 
	\sa_snapshot[11].r.part0[2] , \sa_snapshot[11].r.part0[1] , 
	\sa_snapshot[11].r.part0[0] , \sa_snapshot[10].r.part1[31] , 
	\sa_snapshot[10].r.part1[30] , \sa_snapshot[10].r.part1[29] , 
	\sa_snapshot[10].r.part1[28] , \sa_snapshot[10].r.part1[27] , 
	\sa_snapshot[10].r.part1[26] , \sa_snapshot[10].r.part1[25] , 
	\sa_snapshot[10].r.part1[24] , \sa_snapshot[10].r.part1[23] , 
	\sa_snapshot[10].r.part1[22] , \sa_snapshot[10].r.part1[21] , 
	\sa_snapshot[10].r.part1[20] , \sa_snapshot[10].r.part1[19] , 
	\sa_snapshot[10].r.part1[18] , \sa_snapshot[10].r.part1[17] , 
	\sa_snapshot[10].r.part1[16] , \sa_snapshot[10].r.part1[15] , 
	\sa_snapshot[10].r.part1[14] , \sa_snapshot[10].r.part1[13] , 
	\sa_snapshot[10].r.part1[12] , \sa_snapshot[10].r.part1[11] , 
	\sa_snapshot[10].r.part1[10] , \sa_snapshot[10].r.part1[9] , 
	\sa_snapshot[10].r.part1[8] , \sa_snapshot[10].r.part1[7] , 
	\sa_snapshot[10].r.part1[6] , \sa_snapshot[10].r.part1[5] , 
	\sa_snapshot[10].r.part1[4] , \sa_snapshot[10].r.part1[3] , 
	\sa_snapshot[10].r.part1[2] , \sa_snapshot[10].r.part1[1] , 
	\sa_snapshot[10].r.part1[0] , \sa_snapshot[10].r.part0[31] , 
	\sa_snapshot[10].r.part0[30] , \sa_snapshot[10].r.part0[29] , 
	\sa_snapshot[10].r.part0[28] , \sa_snapshot[10].r.part0[27] , 
	\sa_snapshot[10].r.part0[26] , \sa_snapshot[10].r.part0[25] , 
	\sa_snapshot[10].r.part0[24] , \sa_snapshot[10].r.part0[23] , 
	\sa_snapshot[10].r.part0[22] , \sa_snapshot[10].r.part0[21] , 
	\sa_snapshot[10].r.part0[20] , \sa_snapshot[10].r.part0[19] , 
	\sa_snapshot[10].r.part0[18] , \sa_snapshot[10].r.part0[17] , 
	\sa_snapshot[10].r.part0[16] , \sa_snapshot[10].r.part0[15] , 
	\sa_snapshot[10].r.part0[14] , \sa_snapshot[10].r.part0[13] , 
	\sa_snapshot[10].r.part0[12] , \sa_snapshot[10].r.part0[11] , 
	\sa_snapshot[10].r.part0[10] , \sa_snapshot[10].r.part0[9] , 
	\sa_snapshot[10].r.part0[8] , \sa_snapshot[10].r.part0[7] , 
	\sa_snapshot[10].r.part0[6] , \sa_snapshot[10].r.part0[5] , 
	\sa_snapshot[10].r.part0[4] , \sa_snapshot[10].r.part0[3] , 
	\sa_snapshot[10].r.part0[2] , \sa_snapshot[10].r.part0[1] , 
	\sa_snapshot[10].r.part0[0] , \sa_snapshot[9].r.part1[31] , 
	\sa_snapshot[9].r.part1[30] , \sa_snapshot[9].r.part1[29] , 
	\sa_snapshot[9].r.part1[28] , \sa_snapshot[9].r.part1[27] , 
	\sa_snapshot[9].r.part1[26] , \sa_snapshot[9].r.part1[25] , 
	\sa_snapshot[9].r.part1[24] , \sa_snapshot[9].r.part1[23] , 
	\sa_snapshot[9].r.part1[22] , \sa_snapshot[9].r.part1[21] , 
	\sa_snapshot[9].r.part1[20] , \sa_snapshot[9].r.part1[19] , 
	\sa_snapshot[9].r.part1[18] , \sa_snapshot[9].r.part1[17] , 
	\sa_snapshot[9].r.part1[16] , \sa_snapshot[9].r.part1[15] , 
	\sa_snapshot[9].r.part1[14] , \sa_snapshot[9].r.part1[13] , 
	\sa_snapshot[9].r.part1[12] , \sa_snapshot[9].r.part1[11] , 
	\sa_snapshot[9].r.part1[10] , \sa_snapshot[9].r.part1[9] , 
	\sa_snapshot[9].r.part1[8] , \sa_snapshot[9].r.part1[7] , 
	\sa_snapshot[9].r.part1[6] , \sa_snapshot[9].r.part1[5] , 
	\sa_snapshot[9].r.part1[4] , \sa_snapshot[9].r.part1[3] , 
	\sa_snapshot[9].r.part1[2] , \sa_snapshot[9].r.part1[1] , 
	\sa_snapshot[9].r.part1[0] , \sa_snapshot[9].r.part0[31] , 
	\sa_snapshot[9].r.part0[30] , \sa_snapshot[9].r.part0[29] , 
	\sa_snapshot[9].r.part0[28] , \sa_snapshot[9].r.part0[27] , 
	\sa_snapshot[9].r.part0[26] , \sa_snapshot[9].r.part0[25] , 
	\sa_snapshot[9].r.part0[24] , \sa_snapshot[9].r.part0[23] , 
	\sa_snapshot[9].r.part0[22] , \sa_snapshot[9].r.part0[21] , 
	\sa_snapshot[9].r.part0[20] , \sa_snapshot[9].r.part0[19] , 
	\sa_snapshot[9].r.part0[18] , \sa_snapshot[9].r.part0[17] , 
	\sa_snapshot[9].r.part0[16] , \sa_snapshot[9].r.part0[15] , 
	\sa_snapshot[9].r.part0[14] , \sa_snapshot[9].r.part0[13] , 
	\sa_snapshot[9].r.part0[12] , \sa_snapshot[9].r.part0[11] , 
	\sa_snapshot[9].r.part0[10] , \sa_snapshot[9].r.part0[9] , 
	\sa_snapshot[9].r.part0[8] , \sa_snapshot[9].r.part0[7] , 
	\sa_snapshot[9].r.part0[6] , \sa_snapshot[9].r.part0[5] , 
	\sa_snapshot[9].r.part0[4] , \sa_snapshot[9].r.part0[3] , 
	\sa_snapshot[9].r.part0[2] , \sa_snapshot[9].r.part0[1] , 
	\sa_snapshot[9].r.part0[0] , \sa_snapshot[8].r.part1[31] , 
	\sa_snapshot[8].r.part1[30] , \sa_snapshot[8].r.part1[29] , 
	\sa_snapshot[8].r.part1[28] , \sa_snapshot[8].r.part1[27] , 
	\sa_snapshot[8].r.part1[26] , \sa_snapshot[8].r.part1[25] , 
	\sa_snapshot[8].r.part1[24] , \sa_snapshot[8].r.part1[23] , 
	\sa_snapshot[8].r.part1[22] , \sa_snapshot[8].r.part1[21] , 
	\sa_snapshot[8].r.part1[20] , \sa_snapshot[8].r.part1[19] , 
	\sa_snapshot[8].r.part1[18] , \sa_snapshot[8].r.part1[17] , 
	\sa_snapshot[8].r.part1[16] , \sa_snapshot[8].r.part1[15] , 
	\sa_snapshot[8].r.part1[14] , \sa_snapshot[8].r.part1[13] , 
	\sa_snapshot[8].r.part1[12] , \sa_snapshot[8].r.part1[11] , 
	\sa_snapshot[8].r.part1[10] , \sa_snapshot[8].r.part1[9] , 
	\sa_snapshot[8].r.part1[8] , \sa_snapshot[8].r.part1[7] , 
	\sa_snapshot[8].r.part1[6] , \sa_snapshot[8].r.part1[5] , 
	\sa_snapshot[8].r.part1[4] , \sa_snapshot[8].r.part1[3] , 
	\sa_snapshot[8].r.part1[2] , \sa_snapshot[8].r.part1[1] , 
	\sa_snapshot[8].r.part1[0] , \sa_snapshot[8].r.part0[31] , 
	\sa_snapshot[8].r.part0[30] , \sa_snapshot[8].r.part0[29] , 
	\sa_snapshot[8].r.part0[28] , \sa_snapshot[8].r.part0[27] , 
	\sa_snapshot[8].r.part0[26] , \sa_snapshot[8].r.part0[25] , 
	\sa_snapshot[8].r.part0[24] , \sa_snapshot[8].r.part0[23] , 
	\sa_snapshot[8].r.part0[22] , \sa_snapshot[8].r.part0[21] , 
	\sa_snapshot[8].r.part0[20] , \sa_snapshot[8].r.part0[19] , 
	\sa_snapshot[8].r.part0[18] , \sa_snapshot[8].r.part0[17] , 
	\sa_snapshot[8].r.part0[16] , \sa_snapshot[8].r.part0[15] , 
	\sa_snapshot[8].r.part0[14] , \sa_snapshot[8].r.part0[13] , 
	\sa_snapshot[8].r.part0[12] , \sa_snapshot[8].r.part0[11] , 
	\sa_snapshot[8].r.part0[10] , \sa_snapshot[8].r.part0[9] , 
	\sa_snapshot[8].r.part0[8] , \sa_snapshot[8].r.part0[7] , 
	\sa_snapshot[8].r.part0[6] , \sa_snapshot[8].r.part0[5] , 
	\sa_snapshot[8].r.part0[4] , \sa_snapshot[8].r.part0[3] , 
	\sa_snapshot[8].r.part0[2] , \sa_snapshot[8].r.part0[1] , 
	\sa_snapshot[8].r.part0[0] , \sa_snapshot[7].r.part1[31] , 
	\sa_snapshot[7].r.part1[30] , \sa_snapshot[7].r.part1[29] , 
	\sa_snapshot[7].r.part1[28] , \sa_snapshot[7].r.part1[27] , 
	\sa_snapshot[7].r.part1[26] , \sa_snapshot[7].r.part1[25] , 
	\sa_snapshot[7].r.part1[24] , \sa_snapshot[7].r.part1[23] , 
	\sa_snapshot[7].r.part1[22] , \sa_snapshot[7].r.part1[21] , 
	\sa_snapshot[7].r.part1[20] , \sa_snapshot[7].r.part1[19] , 
	\sa_snapshot[7].r.part1[18] , \sa_snapshot[7].r.part1[17] , 
	\sa_snapshot[7].r.part1[16] , \sa_snapshot[7].r.part1[15] , 
	\sa_snapshot[7].r.part1[14] , \sa_snapshot[7].r.part1[13] , 
	\sa_snapshot[7].r.part1[12] , \sa_snapshot[7].r.part1[11] , 
	\sa_snapshot[7].r.part1[10] , \sa_snapshot[7].r.part1[9] , 
	\sa_snapshot[7].r.part1[8] , \sa_snapshot[7].r.part1[7] , 
	\sa_snapshot[7].r.part1[6] , \sa_snapshot[7].r.part1[5] , 
	\sa_snapshot[7].r.part1[4] , \sa_snapshot[7].r.part1[3] , 
	\sa_snapshot[7].r.part1[2] , \sa_snapshot[7].r.part1[1] , 
	\sa_snapshot[7].r.part1[0] , \sa_snapshot[7].r.part0[31] , 
	\sa_snapshot[7].r.part0[30] , \sa_snapshot[7].r.part0[29] , 
	\sa_snapshot[7].r.part0[28] , \sa_snapshot[7].r.part0[27] , 
	\sa_snapshot[7].r.part0[26] , \sa_snapshot[7].r.part0[25] , 
	\sa_snapshot[7].r.part0[24] , \sa_snapshot[7].r.part0[23] , 
	\sa_snapshot[7].r.part0[22] , \sa_snapshot[7].r.part0[21] , 
	\sa_snapshot[7].r.part0[20] , \sa_snapshot[7].r.part0[19] , 
	\sa_snapshot[7].r.part0[18] , \sa_snapshot[7].r.part0[17] , 
	\sa_snapshot[7].r.part0[16] , \sa_snapshot[7].r.part0[15] , 
	\sa_snapshot[7].r.part0[14] , \sa_snapshot[7].r.part0[13] , 
	\sa_snapshot[7].r.part0[12] , \sa_snapshot[7].r.part0[11] , 
	\sa_snapshot[7].r.part0[10] , \sa_snapshot[7].r.part0[9] , 
	\sa_snapshot[7].r.part0[8] , \sa_snapshot[7].r.part0[7] , 
	\sa_snapshot[7].r.part0[6] , \sa_snapshot[7].r.part0[5] , 
	\sa_snapshot[7].r.part0[4] , \sa_snapshot[7].r.part0[3] , 
	\sa_snapshot[7].r.part0[2] , \sa_snapshot[7].r.part0[1] , 
	\sa_snapshot[7].r.part0[0] , \sa_snapshot[6].r.part1[31] , 
	\sa_snapshot[6].r.part1[30] , \sa_snapshot[6].r.part1[29] , 
	\sa_snapshot[6].r.part1[28] , \sa_snapshot[6].r.part1[27] , 
	\sa_snapshot[6].r.part1[26] , \sa_snapshot[6].r.part1[25] , 
	\sa_snapshot[6].r.part1[24] , \sa_snapshot[6].r.part1[23] , 
	\sa_snapshot[6].r.part1[22] , \sa_snapshot[6].r.part1[21] , 
	\sa_snapshot[6].r.part1[20] , \sa_snapshot[6].r.part1[19] , 
	\sa_snapshot[6].r.part1[18] , \sa_snapshot[6].r.part1[17] , 
	\sa_snapshot[6].r.part1[16] , \sa_snapshot[6].r.part1[15] , 
	\sa_snapshot[6].r.part1[14] , \sa_snapshot[6].r.part1[13] , 
	\sa_snapshot[6].r.part1[12] , \sa_snapshot[6].r.part1[11] , 
	\sa_snapshot[6].r.part1[10] , \sa_snapshot[6].r.part1[9] , 
	\sa_snapshot[6].r.part1[8] , \sa_snapshot[6].r.part1[7] , 
	\sa_snapshot[6].r.part1[6] , \sa_snapshot[6].r.part1[5] , 
	\sa_snapshot[6].r.part1[4] , \sa_snapshot[6].r.part1[3] , 
	\sa_snapshot[6].r.part1[2] , \sa_snapshot[6].r.part1[1] , 
	\sa_snapshot[6].r.part1[0] , \sa_snapshot[6].r.part0[31] , 
	\sa_snapshot[6].r.part0[30] , \sa_snapshot[6].r.part0[29] , 
	\sa_snapshot[6].r.part0[28] , \sa_snapshot[6].r.part0[27] , 
	\sa_snapshot[6].r.part0[26] , \sa_snapshot[6].r.part0[25] , 
	\sa_snapshot[6].r.part0[24] , \sa_snapshot[6].r.part0[23] , 
	\sa_snapshot[6].r.part0[22] , \sa_snapshot[6].r.part0[21] , 
	\sa_snapshot[6].r.part0[20] , \sa_snapshot[6].r.part0[19] , 
	\sa_snapshot[6].r.part0[18] , \sa_snapshot[6].r.part0[17] , 
	\sa_snapshot[6].r.part0[16] , \sa_snapshot[6].r.part0[15] , 
	\sa_snapshot[6].r.part0[14] , \sa_snapshot[6].r.part0[13] , 
	\sa_snapshot[6].r.part0[12] , \sa_snapshot[6].r.part0[11] , 
	\sa_snapshot[6].r.part0[10] , \sa_snapshot[6].r.part0[9] , 
	\sa_snapshot[6].r.part0[8] , \sa_snapshot[6].r.part0[7] , 
	\sa_snapshot[6].r.part0[6] , \sa_snapshot[6].r.part0[5] , 
	\sa_snapshot[6].r.part0[4] , \sa_snapshot[6].r.part0[3] , 
	\sa_snapshot[6].r.part0[2] , \sa_snapshot[6].r.part0[1] , 
	\sa_snapshot[6].r.part0[0] , \sa_snapshot[5].r.part1[31] , 
	\sa_snapshot[5].r.part1[30] , \sa_snapshot[5].r.part1[29] , 
	\sa_snapshot[5].r.part1[28] , \sa_snapshot[5].r.part1[27] , 
	\sa_snapshot[5].r.part1[26] , \sa_snapshot[5].r.part1[25] , 
	\sa_snapshot[5].r.part1[24] , \sa_snapshot[5].r.part1[23] , 
	\sa_snapshot[5].r.part1[22] , \sa_snapshot[5].r.part1[21] , 
	\sa_snapshot[5].r.part1[20] , \sa_snapshot[5].r.part1[19] , 
	\sa_snapshot[5].r.part1[18] , \sa_snapshot[5].r.part1[17] , 
	\sa_snapshot[5].r.part1[16] , \sa_snapshot[5].r.part1[15] , 
	\sa_snapshot[5].r.part1[14] , \sa_snapshot[5].r.part1[13] , 
	\sa_snapshot[5].r.part1[12] , \sa_snapshot[5].r.part1[11] , 
	\sa_snapshot[5].r.part1[10] , \sa_snapshot[5].r.part1[9] , 
	\sa_snapshot[5].r.part1[8] , \sa_snapshot[5].r.part1[7] , 
	\sa_snapshot[5].r.part1[6] , \sa_snapshot[5].r.part1[5] , 
	\sa_snapshot[5].r.part1[4] , \sa_snapshot[5].r.part1[3] , 
	\sa_snapshot[5].r.part1[2] , \sa_snapshot[5].r.part1[1] , 
	\sa_snapshot[5].r.part1[0] , \sa_snapshot[5].r.part0[31] , 
	\sa_snapshot[5].r.part0[30] , \sa_snapshot[5].r.part0[29] , 
	\sa_snapshot[5].r.part0[28] , \sa_snapshot[5].r.part0[27] , 
	\sa_snapshot[5].r.part0[26] , \sa_snapshot[5].r.part0[25] , 
	\sa_snapshot[5].r.part0[24] , \sa_snapshot[5].r.part0[23] , 
	\sa_snapshot[5].r.part0[22] , \sa_snapshot[5].r.part0[21] , 
	\sa_snapshot[5].r.part0[20] , \sa_snapshot[5].r.part0[19] , 
	\sa_snapshot[5].r.part0[18] , \sa_snapshot[5].r.part0[17] , 
	\sa_snapshot[5].r.part0[16] , \sa_snapshot[5].r.part0[15] , 
	\sa_snapshot[5].r.part0[14] , \sa_snapshot[5].r.part0[13] , 
	\sa_snapshot[5].r.part0[12] , \sa_snapshot[5].r.part0[11] , 
	\sa_snapshot[5].r.part0[10] , \sa_snapshot[5].r.part0[9] , 
	\sa_snapshot[5].r.part0[8] , \sa_snapshot[5].r.part0[7] , 
	\sa_snapshot[5].r.part0[6] , \sa_snapshot[5].r.part0[5] , 
	\sa_snapshot[5].r.part0[4] , \sa_snapshot[5].r.part0[3] , 
	\sa_snapshot[5].r.part0[2] , \sa_snapshot[5].r.part0[1] , 
	\sa_snapshot[5].r.part0[0] , \sa_snapshot[4].r.part1[31] , 
	\sa_snapshot[4].r.part1[30] , \sa_snapshot[4].r.part1[29] , 
	\sa_snapshot[4].r.part1[28] , \sa_snapshot[4].r.part1[27] , 
	\sa_snapshot[4].r.part1[26] , \sa_snapshot[4].r.part1[25] , 
	\sa_snapshot[4].r.part1[24] , \sa_snapshot[4].r.part1[23] , 
	\sa_snapshot[4].r.part1[22] , \sa_snapshot[4].r.part1[21] , 
	\sa_snapshot[4].r.part1[20] , \sa_snapshot[4].r.part1[19] , 
	\sa_snapshot[4].r.part1[18] , \sa_snapshot[4].r.part1[17] , 
	\sa_snapshot[4].r.part1[16] , \sa_snapshot[4].r.part1[15] , 
	\sa_snapshot[4].r.part1[14] , \sa_snapshot[4].r.part1[13] , 
	\sa_snapshot[4].r.part1[12] , \sa_snapshot[4].r.part1[11] , 
	\sa_snapshot[4].r.part1[10] , \sa_snapshot[4].r.part1[9] , 
	\sa_snapshot[4].r.part1[8] , \sa_snapshot[4].r.part1[7] , 
	\sa_snapshot[4].r.part1[6] , \sa_snapshot[4].r.part1[5] , 
	\sa_snapshot[4].r.part1[4] , \sa_snapshot[4].r.part1[3] , 
	\sa_snapshot[4].r.part1[2] , \sa_snapshot[4].r.part1[1] , 
	\sa_snapshot[4].r.part1[0] , \sa_snapshot[4].r.part0[31] , 
	\sa_snapshot[4].r.part0[30] , \sa_snapshot[4].r.part0[29] , 
	\sa_snapshot[4].r.part0[28] , \sa_snapshot[4].r.part0[27] , 
	\sa_snapshot[4].r.part0[26] , \sa_snapshot[4].r.part0[25] , 
	\sa_snapshot[4].r.part0[24] , \sa_snapshot[4].r.part0[23] , 
	\sa_snapshot[4].r.part0[22] , \sa_snapshot[4].r.part0[21] , 
	\sa_snapshot[4].r.part0[20] , \sa_snapshot[4].r.part0[19] , 
	\sa_snapshot[4].r.part0[18] , \sa_snapshot[4].r.part0[17] , 
	\sa_snapshot[4].r.part0[16] , \sa_snapshot[4].r.part0[15] , 
	\sa_snapshot[4].r.part0[14] , \sa_snapshot[4].r.part0[13] , 
	\sa_snapshot[4].r.part0[12] , \sa_snapshot[4].r.part0[11] , 
	\sa_snapshot[4].r.part0[10] , \sa_snapshot[4].r.part0[9] , 
	\sa_snapshot[4].r.part0[8] , \sa_snapshot[4].r.part0[7] , 
	\sa_snapshot[4].r.part0[6] , \sa_snapshot[4].r.part0[5] , 
	\sa_snapshot[4].r.part0[4] , \sa_snapshot[4].r.part0[3] , 
	\sa_snapshot[4].r.part0[2] , \sa_snapshot[4].r.part0[1] , 
	\sa_snapshot[4].r.part0[0] , \sa_snapshot[3].r.part1[31] , 
	\sa_snapshot[3].r.part1[30] , \sa_snapshot[3].r.part1[29] , 
	\sa_snapshot[3].r.part1[28] , \sa_snapshot[3].r.part1[27] , 
	\sa_snapshot[3].r.part1[26] , \sa_snapshot[3].r.part1[25] , 
	\sa_snapshot[3].r.part1[24] , \sa_snapshot[3].r.part1[23] , 
	\sa_snapshot[3].r.part1[22] , \sa_snapshot[3].r.part1[21] , 
	\sa_snapshot[3].r.part1[20] , \sa_snapshot[3].r.part1[19] , 
	\sa_snapshot[3].r.part1[18] , \sa_snapshot[3].r.part1[17] , 
	\sa_snapshot[3].r.part1[16] , \sa_snapshot[3].r.part1[15] , 
	\sa_snapshot[3].r.part1[14] , \sa_snapshot[3].r.part1[13] , 
	\sa_snapshot[3].r.part1[12] , \sa_snapshot[3].r.part1[11] , 
	\sa_snapshot[3].r.part1[10] , \sa_snapshot[3].r.part1[9] , 
	\sa_snapshot[3].r.part1[8] , \sa_snapshot[3].r.part1[7] , 
	\sa_snapshot[3].r.part1[6] , \sa_snapshot[3].r.part1[5] , 
	\sa_snapshot[3].r.part1[4] , \sa_snapshot[3].r.part1[3] , 
	\sa_snapshot[3].r.part1[2] , \sa_snapshot[3].r.part1[1] , 
	\sa_snapshot[3].r.part1[0] , \sa_snapshot[3].r.part0[31] , 
	\sa_snapshot[3].r.part0[30] , \sa_snapshot[3].r.part0[29] , 
	\sa_snapshot[3].r.part0[28] , \sa_snapshot[3].r.part0[27] , 
	\sa_snapshot[3].r.part0[26] , \sa_snapshot[3].r.part0[25] , 
	\sa_snapshot[3].r.part0[24] , \sa_snapshot[3].r.part0[23] , 
	\sa_snapshot[3].r.part0[22] , \sa_snapshot[3].r.part0[21] , 
	\sa_snapshot[3].r.part0[20] , \sa_snapshot[3].r.part0[19] , 
	\sa_snapshot[3].r.part0[18] , \sa_snapshot[3].r.part0[17] , 
	\sa_snapshot[3].r.part0[16] , \sa_snapshot[3].r.part0[15] , 
	\sa_snapshot[3].r.part0[14] , \sa_snapshot[3].r.part0[13] , 
	\sa_snapshot[3].r.part0[12] , \sa_snapshot[3].r.part0[11] , 
	\sa_snapshot[3].r.part0[10] , \sa_snapshot[3].r.part0[9] , 
	\sa_snapshot[3].r.part0[8] , \sa_snapshot[3].r.part0[7] , 
	\sa_snapshot[3].r.part0[6] , \sa_snapshot[3].r.part0[5] , 
	\sa_snapshot[3].r.part0[4] , \sa_snapshot[3].r.part0[3] , 
	\sa_snapshot[3].r.part0[2] , \sa_snapshot[3].r.part0[1] , 
	\sa_snapshot[3].r.part0[0] , \sa_snapshot[2].r.part1[31] , 
	\sa_snapshot[2].r.part1[30] , \sa_snapshot[2].r.part1[29] , 
	\sa_snapshot[2].r.part1[28] , \sa_snapshot[2].r.part1[27] , 
	\sa_snapshot[2].r.part1[26] , \sa_snapshot[2].r.part1[25] , 
	\sa_snapshot[2].r.part1[24] , \sa_snapshot[2].r.part1[23] , 
	\sa_snapshot[2].r.part1[22] , \sa_snapshot[2].r.part1[21] , 
	\sa_snapshot[2].r.part1[20] , \sa_snapshot[2].r.part1[19] , 
	\sa_snapshot[2].r.part1[18] , \sa_snapshot[2].r.part1[17] , 
	\sa_snapshot[2].r.part1[16] , \sa_snapshot[2].r.part1[15] , 
	\sa_snapshot[2].r.part1[14] , \sa_snapshot[2].r.part1[13] , 
	\sa_snapshot[2].r.part1[12] , \sa_snapshot[2].r.part1[11] , 
	\sa_snapshot[2].r.part1[10] , \sa_snapshot[2].r.part1[9] , 
	\sa_snapshot[2].r.part1[8] , \sa_snapshot[2].r.part1[7] , 
	\sa_snapshot[2].r.part1[6] , \sa_snapshot[2].r.part1[5] , 
	\sa_snapshot[2].r.part1[4] , \sa_snapshot[2].r.part1[3] , 
	\sa_snapshot[2].r.part1[2] , \sa_snapshot[2].r.part1[1] , 
	\sa_snapshot[2].r.part1[0] , \sa_snapshot[2].r.part0[31] , 
	\sa_snapshot[2].r.part0[30] , \sa_snapshot[2].r.part0[29] , 
	\sa_snapshot[2].r.part0[28] , \sa_snapshot[2].r.part0[27] , 
	\sa_snapshot[2].r.part0[26] , \sa_snapshot[2].r.part0[25] , 
	\sa_snapshot[2].r.part0[24] , \sa_snapshot[2].r.part0[23] , 
	\sa_snapshot[2].r.part0[22] , \sa_snapshot[2].r.part0[21] , 
	\sa_snapshot[2].r.part0[20] , \sa_snapshot[2].r.part0[19] , 
	\sa_snapshot[2].r.part0[18] , \sa_snapshot[2].r.part0[17] , 
	\sa_snapshot[2].r.part0[16] , \sa_snapshot[2].r.part0[15] , 
	\sa_snapshot[2].r.part0[14] , \sa_snapshot[2].r.part0[13] , 
	\sa_snapshot[2].r.part0[12] , \sa_snapshot[2].r.part0[11] , 
	\sa_snapshot[2].r.part0[10] , \sa_snapshot[2].r.part0[9] , 
	\sa_snapshot[2].r.part0[8] , \sa_snapshot[2].r.part0[7] , 
	\sa_snapshot[2].r.part0[6] , \sa_snapshot[2].r.part0[5] , 
	\sa_snapshot[2].r.part0[4] , \sa_snapshot[2].r.part0[3] , 
	\sa_snapshot[2].r.part0[2] , \sa_snapshot[2].r.part0[1] , 
	\sa_snapshot[2].r.part0[0] , \sa_snapshot[1].r.part1[31] , 
	\sa_snapshot[1].r.part1[30] , \sa_snapshot[1].r.part1[29] , 
	\sa_snapshot[1].r.part1[28] , \sa_snapshot[1].r.part1[27] , 
	\sa_snapshot[1].r.part1[26] , \sa_snapshot[1].r.part1[25] , 
	\sa_snapshot[1].r.part1[24] , \sa_snapshot[1].r.part1[23] , 
	\sa_snapshot[1].r.part1[22] , \sa_snapshot[1].r.part1[21] , 
	\sa_snapshot[1].r.part1[20] , \sa_snapshot[1].r.part1[19] , 
	\sa_snapshot[1].r.part1[18] , \sa_snapshot[1].r.part1[17] , 
	\sa_snapshot[1].r.part1[16] , \sa_snapshot[1].r.part1[15] , 
	\sa_snapshot[1].r.part1[14] , \sa_snapshot[1].r.part1[13] , 
	\sa_snapshot[1].r.part1[12] , \sa_snapshot[1].r.part1[11] , 
	\sa_snapshot[1].r.part1[10] , \sa_snapshot[1].r.part1[9] , 
	\sa_snapshot[1].r.part1[8] , \sa_snapshot[1].r.part1[7] , 
	\sa_snapshot[1].r.part1[6] , \sa_snapshot[1].r.part1[5] , 
	\sa_snapshot[1].r.part1[4] , \sa_snapshot[1].r.part1[3] , 
	\sa_snapshot[1].r.part1[2] , \sa_snapshot[1].r.part1[1] , 
	\sa_snapshot[1].r.part1[0] , \sa_snapshot[1].r.part0[31] , 
	\sa_snapshot[1].r.part0[30] , \sa_snapshot[1].r.part0[29] , 
	\sa_snapshot[1].r.part0[28] , \sa_snapshot[1].r.part0[27] , 
	\sa_snapshot[1].r.part0[26] , \sa_snapshot[1].r.part0[25] , 
	\sa_snapshot[1].r.part0[24] , \sa_snapshot[1].r.part0[23] , 
	\sa_snapshot[1].r.part0[22] , \sa_snapshot[1].r.part0[21] , 
	\sa_snapshot[1].r.part0[20] , \sa_snapshot[1].r.part0[19] , 
	\sa_snapshot[1].r.part0[18] , \sa_snapshot[1].r.part0[17] , 
	\sa_snapshot[1].r.part0[16] , \sa_snapshot[1].r.part0[15] , 
	\sa_snapshot[1].r.part0[14] , \sa_snapshot[1].r.part0[13] , 
	\sa_snapshot[1].r.part0[12] , \sa_snapshot[1].r.part0[11] , 
	\sa_snapshot[1].r.part0[10] , \sa_snapshot[1].r.part0[9] , 
	\sa_snapshot[1].r.part0[8] , \sa_snapshot[1].r.part0[7] , 
	\sa_snapshot[1].r.part0[6] , \sa_snapshot[1].r.part0[5] , 
	\sa_snapshot[1].r.part0[4] , \sa_snapshot[1].r.part0[3] , 
	\sa_snapshot[1].r.part0[2] , \sa_snapshot[1].r.part0[1] , 
	\sa_snapshot[1].r.part0[0] , \sa_snapshot[0].r.part1[31] , 
	\sa_snapshot[0].r.part1[30] , \sa_snapshot[0].r.part1[29] , 
	\sa_snapshot[0].r.part1[28] , \sa_snapshot[0].r.part1[27] , 
	\sa_snapshot[0].r.part1[26] , \sa_snapshot[0].r.part1[25] , 
	\sa_snapshot[0].r.part1[24] , \sa_snapshot[0].r.part1[23] , 
	\sa_snapshot[0].r.part1[22] , \sa_snapshot[0].r.part1[21] , 
	\sa_snapshot[0].r.part1[20] , \sa_snapshot[0].r.part1[19] , 
	\sa_snapshot[0].r.part1[18] , \sa_snapshot[0].r.part1[17] , 
	\sa_snapshot[0].r.part1[16] , \sa_snapshot[0].r.part1[15] , 
	\sa_snapshot[0].r.part1[14] , \sa_snapshot[0].r.part1[13] , 
	\sa_snapshot[0].r.part1[12] , \sa_snapshot[0].r.part1[11] , 
	\sa_snapshot[0].r.part1[10] , \sa_snapshot[0].r.part1[9] , 
	\sa_snapshot[0].r.part1[8] , \sa_snapshot[0].r.part1[7] , 
	\sa_snapshot[0].r.part1[6] , \sa_snapshot[0].r.part1[5] , 
	\sa_snapshot[0].r.part1[4] , \sa_snapshot[0].r.part1[3] , 
	\sa_snapshot[0].r.part1[2] , \sa_snapshot[0].r.part1[1] , 
	\sa_snapshot[0].r.part1[0] , \sa_snapshot[0].r.part0[31] , 
	\sa_snapshot[0].r.part0[30] , \sa_snapshot[0].r.part0[29] , 
	\sa_snapshot[0].r.part0[28] , \sa_snapshot[0].r.part0[27] , 
	\sa_snapshot[0].r.part0[26] , \sa_snapshot[0].r.part0[25] , 
	\sa_snapshot[0].r.part0[24] , \sa_snapshot[0].r.part0[23] , 
	\sa_snapshot[0].r.part0[22] , \sa_snapshot[0].r.part0[21] , 
	\sa_snapshot[0].r.part0[20] , \sa_snapshot[0].r.part0[19] , 
	\sa_snapshot[0].r.part0[18] , \sa_snapshot[0].r.part0[17] , 
	\sa_snapshot[0].r.part0[16] , \sa_snapshot[0].r.part0[15] , 
	\sa_snapshot[0].r.part0[14] , \sa_snapshot[0].r.part0[13] , 
	\sa_snapshot[0].r.part0[12] , \sa_snapshot[0].r.part0[11] , 
	\sa_snapshot[0].r.part0[10] , \sa_snapshot[0].r.part0[9] , 
	\sa_snapshot[0].r.part0[8] , \sa_snapshot[0].r.part0[7] , 
	\sa_snapshot[0].r.part0[6] , \sa_snapshot[0].r.part0[5] , 
	\sa_snapshot[0].r.part0[4] , \sa_snapshot[0].r.part0[3] , 
	\sa_snapshot[0].r.part0[2] , \sa_snapshot[0].r.part0[1] , 
	\sa_snapshot[0].r.part0[0] } ), .sa_count( {
	\sa_count[31].r.part1[31] , \sa_count[31].r.part1[30] , 
	\sa_count[31].r.part1[29] , \sa_count[31].r.part1[28] , 
	\sa_count[31].r.part1[27] , \sa_count[31].r.part1[26] , 
	\sa_count[31].r.part1[25] , \sa_count[31].r.part1[24] , 
	\sa_count[31].r.part1[23] , \sa_count[31].r.part1[22] , 
	\sa_count[31].r.part1[21] , \sa_count[31].r.part1[20] , 
	\sa_count[31].r.part1[19] , \sa_count[31].r.part1[18] , 
	\sa_count[31].r.part1[17] , \sa_count[31].r.part1[16] , 
	\sa_count[31].r.part1[15] , \sa_count[31].r.part1[14] , 
	\sa_count[31].r.part1[13] , \sa_count[31].r.part1[12] , 
	\sa_count[31].r.part1[11] , \sa_count[31].r.part1[10] , 
	\sa_count[31].r.part1[9] , \sa_count[31].r.part1[8] , 
	\sa_count[31].r.part1[7] , \sa_count[31].r.part1[6] , 
	\sa_count[31].r.part1[5] , \sa_count[31].r.part1[4] , 
	\sa_count[31].r.part1[3] , \sa_count[31].r.part1[2] , 
	\sa_count[31].r.part1[1] , \sa_count[31].r.part1[0] , 
	\sa_count[31].r.part0[31] , \sa_count[31].r.part0[30] , 
	\sa_count[31].r.part0[29] , \sa_count[31].r.part0[28] , 
	\sa_count[31].r.part0[27] , \sa_count[31].r.part0[26] , 
	\sa_count[31].r.part0[25] , \sa_count[31].r.part0[24] , 
	\sa_count[31].r.part0[23] , \sa_count[31].r.part0[22] , 
	\sa_count[31].r.part0[21] , \sa_count[31].r.part0[20] , 
	\sa_count[31].r.part0[19] , \sa_count[31].r.part0[18] , 
	\sa_count[31].r.part0[17] , \sa_count[31].r.part0[16] , 
	\sa_count[31].r.part0[15] , \sa_count[31].r.part0[14] , 
	\sa_count[31].r.part0[13] , \sa_count[31].r.part0[12] , 
	\sa_count[31].r.part0[11] , \sa_count[31].r.part0[10] , 
	\sa_count[31].r.part0[9] , \sa_count[31].r.part0[8] , 
	\sa_count[31].r.part0[7] , \sa_count[31].r.part0[6] , 
	\sa_count[31].r.part0[5] , \sa_count[31].r.part0[4] , 
	\sa_count[31].r.part0[3] , \sa_count[31].r.part0[2] , 
	\sa_count[31].r.part0[1] , \sa_count[31].r.part0[0] , 
	\sa_count[30].r.part1[31] , \sa_count[30].r.part1[30] , 
	\sa_count[30].r.part1[29] , \sa_count[30].r.part1[28] , 
	\sa_count[30].r.part1[27] , \sa_count[30].r.part1[26] , 
	\sa_count[30].r.part1[25] , \sa_count[30].r.part1[24] , 
	\sa_count[30].r.part1[23] , \sa_count[30].r.part1[22] , 
	\sa_count[30].r.part1[21] , \sa_count[30].r.part1[20] , 
	\sa_count[30].r.part1[19] , \sa_count[30].r.part1[18] , 
	\sa_count[30].r.part1[17] , \sa_count[30].r.part1[16] , 
	\sa_count[30].r.part1[15] , \sa_count[30].r.part1[14] , 
	\sa_count[30].r.part1[13] , \sa_count[30].r.part1[12] , 
	\sa_count[30].r.part1[11] , \sa_count[30].r.part1[10] , 
	\sa_count[30].r.part1[9] , \sa_count[30].r.part1[8] , 
	\sa_count[30].r.part1[7] , \sa_count[30].r.part1[6] , 
	\sa_count[30].r.part1[5] , \sa_count[30].r.part1[4] , 
	\sa_count[30].r.part1[3] , \sa_count[30].r.part1[2] , 
	\sa_count[30].r.part1[1] , \sa_count[30].r.part1[0] , 
	\sa_count[30].r.part0[31] , \sa_count[30].r.part0[30] , 
	\sa_count[30].r.part0[29] , \sa_count[30].r.part0[28] , 
	\sa_count[30].r.part0[27] , \sa_count[30].r.part0[26] , 
	\sa_count[30].r.part0[25] , \sa_count[30].r.part0[24] , 
	\sa_count[30].r.part0[23] , \sa_count[30].r.part0[22] , 
	\sa_count[30].r.part0[21] , \sa_count[30].r.part0[20] , 
	\sa_count[30].r.part0[19] , \sa_count[30].r.part0[18] , 
	\sa_count[30].r.part0[17] , \sa_count[30].r.part0[16] , 
	\sa_count[30].r.part0[15] , \sa_count[30].r.part0[14] , 
	\sa_count[30].r.part0[13] , \sa_count[30].r.part0[12] , 
	\sa_count[30].r.part0[11] , \sa_count[30].r.part0[10] , 
	\sa_count[30].r.part0[9] , \sa_count[30].r.part0[8] , 
	\sa_count[30].r.part0[7] , \sa_count[30].r.part0[6] , 
	\sa_count[30].r.part0[5] , \sa_count[30].r.part0[4] , 
	\sa_count[30].r.part0[3] , \sa_count[30].r.part0[2] , 
	\sa_count[30].r.part0[1] , \sa_count[30].r.part0[0] , 
	\sa_count[29].r.part1[31] , \sa_count[29].r.part1[30] , 
	\sa_count[29].r.part1[29] , \sa_count[29].r.part1[28] , 
	\sa_count[29].r.part1[27] , \sa_count[29].r.part1[26] , 
	\sa_count[29].r.part1[25] , \sa_count[29].r.part1[24] , 
	\sa_count[29].r.part1[23] , \sa_count[29].r.part1[22] , 
	\sa_count[29].r.part1[21] , \sa_count[29].r.part1[20] , 
	\sa_count[29].r.part1[19] , \sa_count[29].r.part1[18] , 
	\sa_count[29].r.part1[17] , \sa_count[29].r.part1[16] , 
	\sa_count[29].r.part1[15] , \sa_count[29].r.part1[14] , 
	\sa_count[29].r.part1[13] , \sa_count[29].r.part1[12] , 
	\sa_count[29].r.part1[11] , \sa_count[29].r.part1[10] , 
	\sa_count[29].r.part1[9] , \sa_count[29].r.part1[8] , 
	\sa_count[29].r.part1[7] , \sa_count[29].r.part1[6] , 
	\sa_count[29].r.part1[5] , \sa_count[29].r.part1[4] , 
	\sa_count[29].r.part1[3] , \sa_count[29].r.part1[2] , 
	\sa_count[29].r.part1[1] , \sa_count[29].r.part1[0] , 
	\sa_count[29].r.part0[31] , \sa_count[29].r.part0[30] , 
	\sa_count[29].r.part0[29] , \sa_count[29].r.part0[28] , 
	\sa_count[29].r.part0[27] , \sa_count[29].r.part0[26] , 
	\sa_count[29].r.part0[25] , \sa_count[29].r.part0[24] , 
	\sa_count[29].r.part0[23] , \sa_count[29].r.part0[22] , 
	\sa_count[29].r.part0[21] , \sa_count[29].r.part0[20] , 
	\sa_count[29].r.part0[19] , \sa_count[29].r.part0[18] , 
	\sa_count[29].r.part0[17] , \sa_count[29].r.part0[16] , 
	\sa_count[29].r.part0[15] , \sa_count[29].r.part0[14] , 
	\sa_count[29].r.part0[13] , \sa_count[29].r.part0[12] , 
	\sa_count[29].r.part0[11] , \sa_count[29].r.part0[10] , 
	\sa_count[29].r.part0[9] , \sa_count[29].r.part0[8] , 
	\sa_count[29].r.part0[7] , \sa_count[29].r.part0[6] , 
	\sa_count[29].r.part0[5] , \sa_count[29].r.part0[4] , 
	\sa_count[29].r.part0[3] , \sa_count[29].r.part0[2] , 
	\sa_count[29].r.part0[1] , \sa_count[29].r.part0[0] , 
	\sa_count[28].r.part1[31] , \sa_count[28].r.part1[30] , 
	\sa_count[28].r.part1[29] , \sa_count[28].r.part1[28] , 
	\sa_count[28].r.part1[27] , \sa_count[28].r.part1[26] , 
	\sa_count[28].r.part1[25] , \sa_count[28].r.part1[24] , 
	\sa_count[28].r.part1[23] , \sa_count[28].r.part1[22] , 
	\sa_count[28].r.part1[21] , \sa_count[28].r.part1[20] , 
	\sa_count[28].r.part1[19] , \sa_count[28].r.part1[18] , 
	\sa_count[28].r.part1[17] , \sa_count[28].r.part1[16] , 
	\sa_count[28].r.part1[15] , \sa_count[28].r.part1[14] , 
	\sa_count[28].r.part1[13] , \sa_count[28].r.part1[12] , 
	\sa_count[28].r.part1[11] , \sa_count[28].r.part1[10] , 
	\sa_count[28].r.part1[9] , \sa_count[28].r.part1[8] , 
	\sa_count[28].r.part1[7] , \sa_count[28].r.part1[6] , 
	\sa_count[28].r.part1[5] , \sa_count[28].r.part1[4] , 
	\sa_count[28].r.part1[3] , \sa_count[28].r.part1[2] , 
	\sa_count[28].r.part1[1] , \sa_count[28].r.part1[0] , 
	\sa_count[28].r.part0[31] , \sa_count[28].r.part0[30] , 
	\sa_count[28].r.part0[29] , \sa_count[28].r.part0[28] , 
	\sa_count[28].r.part0[27] , \sa_count[28].r.part0[26] , 
	\sa_count[28].r.part0[25] , \sa_count[28].r.part0[24] , 
	\sa_count[28].r.part0[23] , \sa_count[28].r.part0[22] , 
	\sa_count[28].r.part0[21] , \sa_count[28].r.part0[20] , 
	\sa_count[28].r.part0[19] , \sa_count[28].r.part0[18] , 
	\sa_count[28].r.part0[17] , \sa_count[28].r.part0[16] , 
	\sa_count[28].r.part0[15] , \sa_count[28].r.part0[14] , 
	\sa_count[28].r.part0[13] , \sa_count[28].r.part0[12] , 
	\sa_count[28].r.part0[11] , \sa_count[28].r.part0[10] , 
	\sa_count[28].r.part0[9] , \sa_count[28].r.part0[8] , 
	\sa_count[28].r.part0[7] , \sa_count[28].r.part0[6] , 
	\sa_count[28].r.part0[5] , \sa_count[28].r.part0[4] , 
	\sa_count[28].r.part0[3] , \sa_count[28].r.part0[2] , 
	\sa_count[28].r.part0[1] , \sa_count[28].r.part0[0] , 
	\sa_count[27].r.part1[31] , \sa_count[27].r.part1[30] , 
	\sa_count[27].r.part1[29] , \sa_count[27].r.part1[28] , 
	\sa_count[27].r.part1[27] , \sa_count[27].r.part1[26] , 
	\sa_count[27].r.part1[25] , \sa_count[27].r.part1[24] , 
	\sa_count[27].r.part1[23] , \sa_count[27].r.part1[22] , 
	\sa_count[27].r.part1[21] , \sa_count[27].r.part1[20] , 
	\sa_count[27].r.part1[19] , \sa_count[27].r.part1[18] , 
	\sa_count[27].r.part1[17] , \sa_count[27].r.part1[16] , 
	\sa_count[27].r.part1[15] , \sa_count[27].r.part1[14] , 
	\sa_count[27].r.part1[13] , \sa_count[27].r.part1[12] , 
	\sa_count[27].r.part1[11] , \sa_count[27].r.part1[10] , 
	\sa_count[27].r.part1[9] , \sa_count[27].r.part1[8] , 
	\sa_count[27].r.part1[7] , \sa_count[27].r.part1[6] , 
	\sa_count[27].r.part1[5] , \sa_count[27].r.part1[4] , 
	\sa_count[27].r.part1[3] , \sa_count[27].r.part1[2] , 
	\sa_count[27].r.part1[1] , \sa_count[27].r.part1[0] , 
	\sa_count[27].r.part0[31] , \sa_count[27].r.part0[30] , 
	\sa_count[27].r.part0[29] , \sa_count[27].r.part0[28] , 
	\sa_count[27].r.part0[27] , \sa_count[27].r.part0[26] , 
	\sa_count[27].r.part0[25] , \sa_count[27].r.part0[24] , 
	\sa_count[27].r.part0[23] , \sa_count[27].r.part0[22] , 
	\sa_count[27].r.part0[21] , \sa_count[27].r.part0[20] , 
	\sa_count[27].r.part0[19] , \sa_count[27].r.part0[18] , 
	\sa_count[27].r.part0[17] , \sa_count[27].r.part0[16] , 
	\sa_count[27].r.part0[15] , \sa_count[27].r.part0[14] , 
	\sa_count[27].r.part0[13] , \sa_count[27].r.part0[12] , 
	\sa_count[27].r.part0[11] , \sa_count[27].r.part0[10] , 
	\sa_count[27].r.part0[9] , \sa_count[27].r.part0[8] , 
	\sa_count[27].r.part0[7] , \sa_count[27].r.part0[6] , 
	\sa_count[27].r.part0[5] , \sa_count[27].r.part0[4] , 
	\sa_count[27].r.part0[3] , \sa_count[27].r.part0[2] , 
	\sa_count[27].r.part0[1] , \sa_count[27].r.part0[0] , 
	\sa_count[26].r.part1[31] , \sa_count[26].r.part1[30] , 
	\sa_count[26].r.part1[29] , \sa_count[26].r.part1[28] , 
	\sa_count[26].r.part1[27] , \sa_count[26].r.part1[26] , 
	\sa_count[26].r.part1[25] , \sa_count[26].r.part1[24] , 
	\sa_count[26].r.part1[23] , \sa_count[26].r.part1[22] , 
	\sa_count[26].r.part1[21] , \sa_count[26].r.part1[20] , 
	\sa_count[26].r.part1[19] , \sa_count[26].r.part1[18] , 
	\sa_count[26].r.part1[17] , \sa_count[26].r.part1[16] , 
	\sa_count[26].r.part1[15] , \sa_count[26].r.part1[14] , 
	\sa_count[26].r.part1[13] , \sa_count[26].r.part1[12] , 
	\sa_count[26].r.part1[11] , \sa_count[26].r.part1[10] , 
	\sa_count[26].r.part1[9] , \sa_count[26].r.part1[8] , 
	\sa_count[26].r.part1[7] , \sa_count[26].r.part1[6] , 
	\sa_count[26].r.part1[5] , \sa_count[26].r.part1[4] , 
	\sa_count[26].r.part1[3] , \sa_count[26].r.part1[2] , 
	\sa_count[26].r.part1[1] , \sa_count[26].r.part1[0] , 
	\sa_count[26].r.part0[31] , \sa_count[26].r.part0[30] , 
	\sa_count[26].r.part0[29] , \sa_count[26].r.part0[28] , 
	\sa_count[26].r.part0[27] , \sa_count[26].r.part0[26] , 
	\sa_count[26].r.part0[25] , \sa_count[26].r.part0[24] , 
	\sa_count[26].r.part0[23] , \sa_count[26].r.part0[22] , 
	\sa_count[26].r.part0[21] , \sa_count[26].r.part0[20] , 
	\sa_count[26].r.part0[19] , \sa_count[26].r.part0[18] , 
	\sa_count[26].r.part0[17] , \sa_count[26].r.part0[16] , 
	\sa_count[26].r.part0[15] , \sa_count[26].r.part0[14] , 
	\sa_count[26].r.part0[13] , \sa_count[26].r.part0[12] , 
	\sa_count[26].r.part0[11] , \sa_count[26].r.part0[10] , 
	\sa_count[26].r.part0[9] , \sa_count[26].r.part0[8] , 
	\sa_count[26].r.part0[7] , \sa_count[26].r.part0[6] , 
	\sa_count[26].r.part0[5] , \sa_count[26].r.part0[4] , 
	\sa_count[26].r.part0[3] , \sa_count[26].r.part0[2] , 
	\sa_count[26].r.part0[1] , \sa_count[26].r.part0[0] , 
	\sa_count[25].r.part1[31] , \sa_count[25].r.part1[30] , 
	\sa_count[25].r.part1[29] , \sa_count[25].r.part1[28] , 
	\sa_count[25].r.part1[27] , \sa_count[25].r.part1[26] , 
	\sa_count[25].r.part1[25] , \sa_count[25].r.part1[24] , 
	\sa_count[25].r.part1[23] , \sa_count[25].r.part1[22] , 
	\sa_count[25].r.part1[21] , \sa_count[25].r.part1[20] , 
	\sa_count[25].r.part1[19] , \sa_count[25].r.part1[18] , 
	\sa_count[25].r.part1[17] , \sa_count[25].r.part1[16] , 
	\sa_count[25].r.part1[15] , \sa_count[25].r.part1[14] , 
	\sa_count[25].r.part1[13] , \sa_count[25].r.part1[12] , 
	\sa_count[25].r.part1[11] , \sa_count[25].r.part1[10] , 
	\sa_count[25].r.part1[9] , \sa_count[25].r.part1[8] , 
	\sa_count[25].r.part1[7] , \sa_count[25].r.part1[6] , 
	\sa_count[25].r.part1[5] , \sa_count[25].r.part1[4] , 
	\sa_count[25].r.part1[3] , \sa_count[25].r.part1[2] , 
	\sa_count[25].r.part1[1] , \sa_count[25].r.part1[0] , 
	\sa_count[25].r.part0[31] , \sa_count[25].r.part0[30] , 
	\sa_count[25].r.part0[29] , \sa_count[25].r.part0[28] , 
	\sa_count[25].r.part0[27] , \sa_count[25].r.part0[26] , 
	\sa_count[25].r.part0[25] , \sa_count[25].r.part0[24] , 
	\sa_count[25].r.part0[23] , \sa_count[25].r.part0[22] , 
	\sa_count[25].r.part0[21] , \sa_count[25].r.part0[20] , 
	\sa_count[25].r.part0[19] , \sa_count[25].r.part0[18] , 
	\sa_count[25].r.part0[17] , \sa_count[25].r.part0[16] , 
	\sa_count[25].r.part0[15] , \sa_count[25].r.part0[14] , 
	\sa_count[25].r.part0[13] , \sa_count[25].r.part0[12] , 
	\sa_count[25].r.part0[11] , \sa_count[25].r.part0[10] , 
	\sa_count[25].r.part0[9] , \sa_count[25].r.part0[8] , 
	\sa_count[25].r.part0[7] , \sa_count[25].r.part0[6] , 
	\sa_count[25].r.part0[5] , \sa_count[25].r.part0[4] , 
	\sa_count[25].r.part0[3] , \sa_count[25].r.part0[2] , 
	\sa_count[25].r.part0[1] , \sa_count[25].r.part0[0] , 
	\sa_count[24].r.part1[31] , \sa_count[24].r.part1[30] , 
	\sa_count[24].r.part1[29] , \sa_count[24].r.part1[28] , 
	\sa_count[24].r.part1[27] , \sa_count[24].r.part1[26] , 
	\sa_count[24].r.part1[25] , \sa_count[24].r.part1[24] , 
	\sa_count[24].r.part1[23] , \sa_count[24].r.part1[22] , 
	\sa_count[24].r.part1[21] , \sa_count[24].r.part1[20] , 
	\sa_count[24].r.part1[19] , \sa_count[24].r.part1[18] , 
	\sa_count[24].r.part1[17] , \sa_count[24].r.part1[16] , 
	\sa_count[24].r.part1[15] , \sa_count[24].r.part1[14] , 
	\sa_count[24].r.part1[13] , \sa_count[24].r.part1[12] , 
	\sa_count[24].r.part1[11] , \sa_count[24].r.part1[10] , 
	\sa_count[24].r.part1[9] , \sa_count[24].r.part1[8] , 
	\sa_count[24].r.part1[7] , \sa_count[24].r.part1[6] , 
	\sa_count[24].r.part1[5] , \sa_count[24].r.part1[4] , 
	\sa_count[24].r.part1[3] , \sa_count[24].r.part1[2] , 
	\sa_count[24].r.part1[1] , \sa_count[24].r.part1[0] , 
	\sa_count[24].r.part0[31] , \sa_count[24].r.part0[30] , 
	\sa_count[24].r.part0[29] , \sa_count[24].r.part0[28] , 
	\sa_count[24].r.part0[27] , \sa_count[24].r.part0[26] , 
	\sa_count[24].r.part0[25] , \sa_count[24].r.part0[24] , 
	\sa_count[24].r.part0[23] , \sa_count[24].r.part0[22] , 
	\sa_count[24].r.part0[21] , \sa_count[24].r.part0[20] , 
	\sa_count[24].r.part0[19] , \sa_count[24].r.part0[18] , 
	\sa_count[24].r.part0[17] , \sa_count[24].r.part0[16] , 
	\sa_count[24].r.part0[15] , \sa_count[24].r.part0[14] , 
	\sa_count[24].r.part0[13] , \sa_count[24].r.part0[12] , 
	\sa_count[24].r.part0[11] , \sa_count[24].r.part0[10] , 
	\sa_count[24].r.part0[9] , \sa_count[24].r.part0[8] , 
	\sa_count[24].r.part0[7] , \sa_count[24].r.part0[6] , 
	\sa_count[24].r.part0[5] , \sa_count[24].r.part0[4] , 
	\sa_count[24].r.part0[3] , \sa_count[24].r.part0[2] , 
	\sa_count[24].r.part0[1] , \sa_count[24].r.part0[0] , 
	\sa_count[23].r.part1[31] , \sa_count[23].r.part1[30] , 
	\sa_count[23].r.part1[29] , \sa_count[23].r.part1[28] , 
	\sa_count[23].r.part1[27] , \sa_count[23].r.part1[26] , 
	\sa_count[23].r.part1[25] , \sa_count[23].r.part1[24] , 
	\sa_count[23].r.part1[23] , \sa_count[23].r.part1[22] , 
	\sa_count[23].r.part1[21] , \sa_count[23].r.part1[20] , 
	\sa_count[23].r.part1[19] , \sa_count[23].r.part1[18] , 
	\sa_count[23].r.part1[17] , \sa_count[23].r.part1[16] , 
	\sa_count[23].r.part1[15] , \sa_count[23].r.part1[14] , 
	\sa_count[23].r.part1[13] , \sa_count[23].r.part1[12] , 
	\sa_count[23].r.part1[11] , \sa_count[23].r.part1[10] , 
	\sa_count[23].r.part1[9] , \sa_count[23].r.part1[8] , 
	\sa_count[23].r.part1[7] , \sa_count[23].r.part1[6] , 
	\sa_count[23].r.part1[5] , \sa_count[23].r.part1[4] , 
	\sa_count[23].r.part1[3] , \sa_count[23].r.part1[2] , 
	\sa_count[23].r.part1[1] , \sa_count[23].r.part1[0] , 
	\sa_count[23].r.part0[31] , \sa_count[23].r.part0[30] , 
	\sa_count[23].r.part0[29] , \sa_count[23].r.part0[28] , 
	\sa_count[23].r.part0[27] , \sa_count[23].r.part0[26] , 
	\sa_count[23].r.part0[25] , \sa_count[23].r.part0[24] , 
	\sa_count[23].r.part0[23] , \sa_count[23].r.part0[22] , 
	\sa_count[23].r.part0[21] , \sa_count[23].r.part0[20] , 
	\sa_count[23].r.part0[19] , \sa_count[23].r.part0[18] , 
	\sa_count[23].r.part0[17] , \sa_count[23].r.part0[16] , 
	\sa_count[23].r.part0[15] , \sa_count[23].r.part0[14] , 
	\sa_count[23].r.part0[13] , \sa_count[23].r.part0[12] , 
	\sa_count[23].r.part0[11] , \sa_count[23].r.part0[10] , 
	\sa_count[23].r.part0[9] , \sa_count[23].r.part0[8] , 
	\sa_count[23].r.part0[7] , \sa_count[23].r.part0[6] , 
	\sa_count[23].r.part0[5] , \sa_count[23].r.part0[4] , 
	\sa_count[23].r.part0[3] , \sa_count[23].r.part0[2] , 
	\sa_count[23].r.part0[1] , \sa_count[23].r.part0[0] , 
	\sa_count[22].r.part1[31] , \sa_count[22].r.part1[30] , 
	\sa_count[22].r.part1[29] , \sa_count[22].r.part1[28] , 
	\sa_count[22].r.part1[27] , \sa_count[22].r.part1[26] , 
	\sa_count[22].r.part1[25] , \sa_count[22].r.part1[24] , 
	\sa_count[22].r.part1[23] , \sa_count[22].r.part1[22] , 
	\sa_count[22].r.part1[21] , \sa_count[22].r.part1[20] , 
	\sa_count[22].r.part1[19] , \sa_count[22].r.part1[18] , 
	\sa_count[22].r.part1[17] , \sa_count[22].r.part1[16] , 
	\sa_count[22].r.part1[15] , \sa_count[22].r.part1[14] , 
	\sa_count[22].r.part1[13] , \sa_count[22].r.part1[12] , 
	\sa_count[22].r.part1[11] , \sa_count[22].r.part1[10] , 
	\sa_count[22].r.part1[9] , \sa_count[22].r.part1[8] , 
	\sa_count[22].r.part1[7] , \sa_count[22].r.part1[6] , 
	\sa_count[22].r.part1[5] , \sa_count[22].r.part1[4] , 
	\sa_count[22].r.part1[3] , \sa_count[22].r.part1[2] , 
	\sa_count[22].r.part1[1] , \sa_count[22].r.part1[0] , 
	\sa_count[22].r.part0[31] , \sa_count[22].r.part0[30] , 
	\sa_count[22].r.part0[29] , \sa_count[22].r.part0[28] , 
	\sa_count[22].r.part0[27] , \sa_count[22].r.part0[26] , 
	\sa_count[22].r.part0[25] , \sa_count[22].r.part0[24] , 
	\sa_count[22].r.part0[23] , \sa_count[22].r.part0[22] , 
	\sa_count[22].r.part0[21] , \sa_count[22].r.part0[20] , 
	\sa_count[22].r.part0[19] , \sa_count[22].r.part0[18] , 
	\sa_count[22].r.part0[17] , \sa_count[22].r.part0[16] , 
	\sa_count[22].r.part0[15] , \sa_count[22].r.part0[14] , 
	\sa_count[22].r.part0[13] , \sa_count[22].r.part0[12] , 
	\sa_count[22].r.part0[11] , \sa_count[22].r.part0[10] , 
	\sa_count[22].r.part0[9] , \sa_count[22].r.part0[8] , 
	\sa_count[22].r.part0[7] , \sa_count[22].r.part0[6] , 
	\sa_count[22].r.part0[5] , \sa_count[22].r.part0[4] , 
	\sa_count[22].r.part0[3] , \sa_count[22].r.part0[2] , 
	\sa_count[22].r.part0[1] , \sa_count[22].r.part0[0] , 
	\sa_count[21].r.part1[31] , \sa_count[21].r.part1[30] , 
	\sa_count[21].r.part1[29] , \sa_count[21].r.part1[28] , 
	\sa_count[21].r.part1[27] , \sa_count[21].r.part1[26] , 
	\sa_count[21].r.part1[25] , \sa_count[21].r.part1[24] , 
	\sa_count[21].r.part1[23] , \sa_count[21].r.part1[22] , 
	\sa_count[21].r.part1[21] , \sa_count[21].r.part1[20] , 
	\sa_count[21].r.part1[19] , \sa_count[21].r.part1[18] , 
	\sa_count[21].r.part1[17] , \sa_count[21].r.part1[16] , 
	\sa_count[21].r.part1[15] , \sa_count[21].r.part1[14] , 
	\sa_count[21].r.part1[13] , \sa_count[21].r.part1[12] , 
	\sa_count[21].r.part1[11] , \sa_count[21].r.part1[10] , 
	\sa_count[21].r.part1[9] , \sa_count[21].r.part1[8] , 
	\sa_count[21].r.part1[7] , \sa_count[21].r.part1[6] , 
	\sa_count[21].r.part1[5] , \sa_count[21].r.part1[4] , 
	\sa_count[21].r.part1[3] , \sa_count[21].r.part1[2] , 
	\sa_count[21].r.part1[1] , \sa_count[21].r.part1[0] , 
	\sa_count[21].r.part0[31] , \sa_count[21].r.part0[30] , 
	\sa_count[21].r.part0[29] , \sa_count[21].r.part0[28] , 
	\sa_count[21].r.part0[27] , \sa_count[21].r.part0[26] , 
	\sa_count[21].r.part0[25] , \sa_count[21].r.part0[24] , 
	\sa_count[21].r.part0[23] , \sa_count[21].r.part0[22] , 
	\sa_count[21].r.part0[21] , \sa_count[21].r.part0[20] , 
	\sa_count[21].r.part0[19] , \sa_count[21].r.part0[18] , 
	\sa_count[21].r.part0[17] , \sa_count[21].r.part0[16] , 
	\sa_count[21].r.part0[15] , \sa_count[21].r.part0[14] , 
	\sa_count[21].r.part0[13] , \sa_count[21].r.part0[12] , 
	\sa_count[21].r.part0[11] , \sa_count[21].r.part0[10] , 
	\sa_count[21].r.part0[9] , \sa_count[21].r.part0[8] , 
	\sa_count[21].r.part0[7] , \sa_count[21].r.part0[6] , 
	\sa_count[21].r.part0[5] , \sa_count[21].r.part0[4] , 
	\sa_count[21].r.part0[3] , \sa_count[21].r.part0[2] , 
	\sa_count[21].r.part0[1] , \sa_count[21].r.part0[0] , 
	\sa_count[20].r.part1[31] , \sa_count[20].r.part1[30] , 
	\sa_count[20].r.part1[29] , \sa_count[20].r.part1[28] , 
	\sa_count[20].r.part1[27] , \sa_count[20].r.part1[26] , 
	\sa_count[20].r.part1[25] , \sa_count[20].r.part1[24] , 
	\sa_count[20].r.part1[23] , \sa_count[20].r.part1[22] , 
	\sa_count[20].r.part1[21] , \sa_count[20].r.part1[20] , 
	\sa_count[20].r.part1[19] , \sa_count[20].r.part1[18] , 
	\sa_count[20].r.part1[17] , \sa_count[20].r.part1[16] , 
	\sa_count[20].r.part1[15] , \sa_count[20].r.part1[14] , 
	\sa_count[20].r.part1[13] , \sa_count[20].r.part1[12] , 
	\sa_count[20].r.part1[11] , \sa_count[20].r.part1[10] , 
	\sa_count[20].r.part1[9] , \sa_count[20].r.part1[8] , 
	\sa_count[20].r.part1[7] , \sa_count[20].r.part1[6] , 
	\sa_count[20].r.part1[5] , \sa_count[20].r.part1[4] , 
	\sa_count[20].r.part1[3] , \sa_count[20].r.part1[2] , 
	\sa_count[20].r.part1[1] , \sa_count[20].r.part1[0] , 
	\sa_count[20].r.part0[31] , \sa_count[20].r.part0[30] , 
	\sa_count[20].r.part0[29] , \sa_count[20].r.part0[28] , 
	\sa_count[20].r.part0[27] , \sa_count[20].r.part0[26] , 
	\sa_count[20].r.part0[25] , \sa_count[20].r.part0[24] , 
	\sa_count[20].r.part0[23] , \sa_count[20].r.part0[22] , 
	\sa_count[20].r.part0[21] , \sa_count[20].r.part0[20] , 
	\sa_count[20].r.part0[19] , \sa_count[20].r.part0[18] , 
	\sa_count[20].r.part0[17] , \sa_count[20].r.part0[16] , 
	\sa_count[20].r.part0[15] , \sa_count[20].r.part0[14] , 
	\sa_count[20].r.part0[13] , \sa_count[20].r.part0[12] , 
	\sa_count[20].r.part0[11] , \sa_count[20].r.part0[10] , 
	\sa_count[20].r.part0[9] , \sa_count[20].r.part0[8] , 
	\sa_count[20].r.part0[7] , \sa_count[20].r.part0[6] , 
	\sa_count[20].r.part0[5] , \sa_count[20].r.part0[4] , 
	\sa_count[20].r.part0[3] , \sa_count[20].r.part0[2] , 
	\sa_count[20].r.part0[1] , \sa_count[20].r.part0[0] , 
	\sa_count[19].r.part1[31] , \sa_count[19].r.part1[30] , 
	\sa_count[19].r.part1[29] , \sa_count[19].r.part1[28] , 
	\sa_count[19].r.part1[27] , \sa_count[19].r.part1[26] , 
	\sa_count[19].r.part1[25] , \sa_count[19].r.part1[24] , 
	\sa_count[19].r.part1[23] , \sa_count[19].r.part1[22] , 
	\sa_count[19].r.part1[21] , \sa_count[19].r.part1[20] , 
	\sa_count[19].r.part1[19] , \sa_count[19].r.part1[18] , 
	\sa_count[19].r.part1[17] , \sa_count[19].r.part1[16] , 
	\sa_count[19].r.part1[15] , \sa_count[19].r.part1[14] , 
	\sa_count[19].r.part1[13] , \sa_count[19].r.part1[12] , 
	\sa_count[19].r.part1[11] , \sa_count[19].r.part1[10] , 
	\sa_count[19].r.part1[9] , \sa_count[19].r.part1[8] , 
	\sa_count[19].r.part1[7] , \sa_count[19].r.part1[6] , 
	\sa_count[19].r.part1[5] , \sa_count[19].r.part1[4] , 
	\sa_count[19].r.part1[3] , \sa_count[19].r.part1[2] , 
	\sa_count[19].r.part1[1] , \sa_count[19].r.part1[0] , 
	\sa_count[19].r.part0[31] , \sa_count[19].r.part0[30] , 
	\sa_count[19].r.part0[29] , \sa_count[19].r.part0[28] , 
	\sa_count[19].r.part0[27] , \sa_count[19].r.part0[26] , 
	\sa_count[19].r.part0[25] , \sa_count[19].r.part0[24] , 
	\sa_count[19].r.part0[23] , \sa_count[19].r.part0[22] , 
	\sa_count[19].r.part0[21] , \sa_count[19].r.part0[20] , 
	\sa_count[19].r.part0[19] , \sa_count[19].r.part0[18] , 
	\sa_count[19].r.part0[17] , \sa_count[19].r.part0[16] , 
	\sa_count[19].r.part0[15] , \sa_count[19].r.part0[14] , 
	\sa_count[19].r.part0[13] , \sa_count[19].r.part0[12] , 
	\sa_count[19].r.part0[11] , \sa_count[19].r.part0[10] , 
	\sa_count[19].r.part0[9] , \sa_count[19].r.part0[8] , 
	\sa_count[19].r.part0[7] , \sa_count[19].r.part0[6] , 
	\sa_count[19].r.part0[5] , \sa_count[19].r.part0[4] , 
	\sa_count[19].r.part0[3] , \sa_count[19].r.part0[2] , 
	\sa_count[19].r.part0[1] , \sa_count[19].r.part0[0] , 
	\sa_count[18].r.part1[31] , \sa_count[18].r.part1[30] , 
	\sa_count[18].r.part1[29] , \sa_count[18].r.part1[28] , 
	\sa_count[18].r.part1[27] , \sa_count[18].r.part1[26] , 
	\sa_count[18].r.part1[25] , \sa_count[18].r.part1[24] , 
	\sa_count[18].r.part1[23] , \sa_count[18].r.part1[22] , 
	\sa_count[18].r.part1[21] , \sa_count[18].r.part1[20] , 
	\sa_count[18].r.part1[19] , \sa_count[18].r.part1[18] , 
	\sa_count[18].r.part1[17] , \sa_count[18].r.part1[16] , 
	\sa_count[18].r.part1[15] , \sa_count[18].r.part1[14] , 
	\sa_count[18].r.part1[13] , \sa_count[18].r.part1[12] , 
	\sa_count[18].r.part1[11] , \sa_count[18].r.part1[10] , 
	\sa_count[18].r.part1[9] , \sa_count[18].r.part1[8] , 
	\sa_count[18].r.part1[7] , \sa_count[18].r.part1[6] , 
	\sa_count[18].r.part1[5] , \sa_count[18].r.part1[4] , 
	\sa_count[18].r.part1[3] , \sa_count[18].r.part1[2] , 
	\sa_count[18].r.part1[1] , \sa_count[18].r.part1[0] , 
	\sa_count[18].r.part0[31] , \sa_count[18].r.part0[30] , 
	\sa_count[18].r.part0[29] , \sa_count[18].r.part0[28] , 
	\sa_count[18].r.part0[27] , \sa_count[18].r.part0[26] , 
	\sa_count[18].r.part0[25] , \sa_count[18].r.part0[24] , 
	\sa_count[18].r.part0[23] , \sa_count[18].r.part0[22] , 
	\sa_count[18].r.part0[21] , \sa_count[18].r.part0[20] , 
	\sa_count[18].r.part0[19] , \sa_count[18].r.part0[18] , 
	\sa_count[18].r.part0[17] , \sa_count[18].r.part0[16] , 
	\sa_count[18].r.part0[15] , \sa_count[18].r.part0[14] , 
	\sa_count[18].r.part0[13] , \sa_count[18].r.part0[12] , 
	\sa_count[18].r.part0[11] , \sa_count[18].r.part0[10] , 
	\sa_count[18].r.part0[9] , \sa_count[18].r.part0[8] , 
	\sa_count[18].r.part0[7] , \sa_count[18].r.part0[6] , 
	\sa_count[18].r.part0[5] , \sa_count[18].r.part0[4] , 
	\sa_count[18].r.part0[3] , \sa_count[18].r.part0[2] , 
	\sa_count[18].r.part0[1] , \sa_count[18].r.part0[0] , 
	\sa_count[17].r.part1[31] , \sa_count[17].r.part1[30] , 
	\sa_count[17].r.part1[29] , \sa_count[17].r.part1[28] , 
	\sa_count[17].r.part1[27] , \sa_count[17].r.part1[26] , 
	\sa_count[17].r.part1[25] , \sa_count[17].r.part1[24] , 
	\sa_count[17].r.part1[23] , \sa_count[17].r.part1[22] , 
	\sa_count[17].r.part1[21] , \sa_count[17].r.part1[20] , 
	\sa_count[17].r.part1[19] , \sa_count[17].r.part1[18] , 
	\sa_count[17].r.part1[17] , \sa_count[17].r.part1[16] , 
	\sa_count[17].r.part1[15] , \sa_count[17].r.part1[14] , 
	\sa_count[17].r.part1[13] , \sa_count[17].r.part1[12] , 
	\sa_count[17].r.part1[11] , \sa_count[17].r.part1[10] , 
	\sa_count[17].r.part1[9] , \sa_count[17].r.part1[8] , 
	\sa_count[17].r.part1[7] , \sa_count[17].r.part1[6] , 
	\sa_count[17].r.part1[5] , \sa_count[17].r.part1[4] , 
	\sa_count[17].r.part1[3] , \sa_count[17].r.part1[2] , 
	\sa_count[17].r.part1[1] , \sa_count[17].r.part1[0] , 
	\sa_count[17].r.part0[31] , \sa_count[17].r.part0[30] , 
	\sa_count[17].r.part0[29] , \sa_count[17].r.part0[28] , 
	\sa_count[17].r.part0[27] , \sa_count[17].r.part0[26] , 
	\sa_count[17].r.part0[25] , \sa_count[17].r.part0[24] , 
	\sa_count[17].r.part0[23] , \sa_count[17].r.part0[22] , 
	\sa_count[17].r.part0[21] , \sa_count[17].r.part0[20] , 
	\sa_count[17].r.part0[19] , \sa_count[17].r.part0[18] , 
	\sa_count[17].r.part0[17] , \sa_count[17].r.part0[16] , 
	\sa_count[17].r.part0[15] , \sa_count[17].r.part0[14] , 
	\sa_count[17].r.part0[13] , \sa_count[17].r.part0[12] , 
	\sa_count[17].r.part0[11] , \sa_count[17].r.part0[10] , 
	\sa_count[17].r.part0[9] , \sa_count[17].r.part0[8] , 
	\sa_count[17].r.part0[7] , \sa_count[17].r.part0[6] , 
	\sa_count[17].r.part0[5] , \sa_count[17].r.part0[4] , 
	\sa_count[17].r.part0[3] , \sa_count[17].r.part0[2] , 
	\sa_count[17].r.part0[1] , \sa_count[17].r.part0[0] , 
	\sa_count[16].r.part1[31] , \sa_count[16].r.part1[30] , 
	\sa_count[16].r.part1[29] , \sa_count[16].r.part1[28] , 
	\sa_count[16].r.part1[27] , \sa_count[16].r.part1[26] , 
	\sa_count[16].r.part1[25] , \sa_count[16].r.part1[24] , 
	\sa_count[16].r.part1[23] , \sa_count[16].r.part1[22] , 
	\sa_count[16].r.part1[21] , \sa_count[16].r.part1[20] , 
	\sa_count[16].r.part1[19] , \sa_count[16].r.part1[18] , 
	\sa_count[16].r.part1[17] , \sa_count[16].r.part1[16] , 
	\sa_count[16].r.part1[15] , \sa_count[16].r.part1[14] , 
	\sa_count[16].r.part1[13] , \sa_count[16].r.part1[12] , 
	\sa_count[16].r.part1[11] , \sa_count[16].r.part1[10] , 
	\sa_count[16].r.part1[9] , \sa_count[16].r.part1[8] , 
	\sa_count[16].r.part1[7] , \sa_count[16].r.part1[6] , 
	\sa_count[16].r.part1[5] , \sa_count[16].r.part1[4] , 
	\sa_count[16].r.part1[3] , \sa_count[16].r.part1[2] , 
	\sa_count[16].r.part1[1] , \sa_count[16].r.part1[0] , 
	\sa_count[16].r.part0[31] , \sa_count[16].r.part0[30] , 
	\sa_count[16].r.part0[29] , \sa_count[16].r.part0[28] , 
	\sa_count[16].r.part0[27] , \sa_count[16].r.part0[26] , 
	\sa_count[16].r.part0[25] , \sa_count[16].r.part0[24] , 
	\sa_count[16].r.part0[23] , \sa_count[16].r.part0[22] , 
	\sa_count[16].r.part0[21] , \sa_count[16].r.part0[20] , 
	\sa_count[16].r.part0[19] , \sa_count[16].r.part0[18] , 
	\sa_count[16].r.part0[17] , \sa_count[16].r.part0[16] , 
	\sa_count[16].r.part0[15] , \sa_count[16].r.part0[14] , 
	\sa_count[16].r.part0[13] , \sa_count[16].r.part0[12] , 
	\sa_count[16].r.part0[11] , \sa_count[16].r.part0[10] , 
	\sa_count[16].r.part0[9] , \sa_count[16].r.part0[8] , 
	\sa_count[16].r.part0[7] , \sa_count[16].r.part0[6] , 
	\sa_count[16].r.part0[5] , \sa_count[16].r.part0[4] , 
	\sa_count[16].r.part0[3] , \sa_count[16].r.part0[2] , 
	\sa_count[16].r.part0[1] , \sa_count[16].r.part0[0] , 
	\sa_count[15].r.part1[31] , \sa_count[15].r.part1[30] , 
	\sa_count[15].r.part1[29] , \sa_count[15].r.part1[28] , 
	\sa_count[15].r.part1[27] , \sa_count[15].r.part1[26] , 
	\sa_count[15].r.part1[25] , \sa_count[15].r.part1[24] , 
	\sa_count[15].r.part1[23] , \sa_count[15].r.part1[22] , 
	\sa_count[15].r.part1[21] , \sa_count[15].r.part1[20] , 
	\sa_count[15].r.part1[19] , \sa_count[15].r.part1[18] , 
	\sa_count[15].r.part1[17] , \sa_count[15].r.part1[16] , 
	\sa_count[15].r.part1[15] , \sa_count[15].r.part1[14] , 
	\sa_count[15].r.part1[13] , \sa_count[15].r.part1[12] , 
	\sa_count[15].r.part1[11] , \sa_count[15].r.part1[10] , 
	\sa_count[15].r.part1[9] , \sa_count[15].r.part1[8] , 
	\sa_count[15].r.part1[7] , \sa_count[15].r.part1[6] , 
	\sa_count[15].r.part1[5] , \sa_count[15].r.part1[4] , 
	\sa_count[15].r.part1[3] , \sa_count[15].r.part1[2] , 
	\sa_count[15].r.part1[1] , \sa_count[15].r.part1[0] , 
	\sa_count[15].r.part0[31] , \sa_count[15].r.part0[30] , 
	\sa_count[15].r.part0[29] , \sa_count[15].r.part0[28] , 
	\sa_count[15].r.part0[27] , \sa_count[15].r.part0[26] , 
	\sa_count[15].r.part0[25] , \sa_count[15].r.part0[24] , 
	\sa_count[15].r.part0[23] , \sa_count[15].r.part0[22] , 
	\sa_count[15].r.part0[21] , \sa_count[15].r.part0[20] , 
	\sa_count[15].r.part0[19] , \sa_count[15].r.part0[18] , 
	\sa_count[15].r.part0[17] , \sa_count[15].r.part0[16] , 
	\sa_count[15].r.part0[15] , \sa_count[15].r.part0[14] , 
	\sa_count[15].r.part0[13] , \sa_count[15].r.part0[12] , 
	\sa_count[15].r.part0[11] , \sa_count[15].r.part0[10] , 
	\sa_count[15].r.part0[9] , \sa_count[15].r.part0[8] , 
	\sa_count[15].r.part0[7] , \sa_count[15].r.part0[6] , 
	\sa_count[15].r.part0[5] , \sa_count[15].r.part0[4] , 
	\sa_count[15].r.part0[3] , \sa_count[15].r.part0[2] , 
	\sa_count[15].r.part0[1] , \sa_count[15].r.part0[0] , 
	\sa_count[14].r.part1[31] , \sa_count[14].r.part1[30] , 
	\sa_count[14].r.part1[29] , \sa_count[14].r.part1[28] , 
	\sa_count[14].r.part1[27] , \sa_count[14].r.part1[26] , 
	\sa_count[14].r.part1[25] , \sa_count[14].r.part1[24] , 
	\sa_count[14].r.part1[23] , \sa_count[14].r.part1[22] , 
	\sa_count[14].r.part1[21] , \sa_count[14].r.part1[20] , 
	\sa_count[14].r.part1[19] , \sa_count[14].r.part1[18] , 
	\sa_count[14].r.part1[17] , \sa_count[14].r.part1[16] , 
	\sa_count[14].r.part1[15] , \sa_count[14].r.part1[14] , 
	\sa_count[14].r.part1[13] , \sa_count[14].r.part1[12] , 
	\sa_count[14].r.part1[11] , \sa_count[14].r.part1[10] , 
	\sa_count[14].r.part1[9] , \sa_count[14].r.part1[8] , 
	\sa_count[14].r.part1[7] , \sa_count[14].r.part1[6] , 
	\sa_count[14].r.part1[5] , \sa_count[14].r.part1[4] , 
	\sa_count[14].r.part1[3] , \sa_count[14].r.part1[2] , 
	\sa_count[14].r.part1[1] , \sa_count[14].r.part1[0] , 
	\sa_count[14].r.part0[31] , \sa_count[14].r.part0[30] , 
	\sa_count[14].r.part0[29] , \sa_count[14].r.part0[28] , 
	\sa_count[14].r.part0[27] , \sa_count[14].r.part0[26] , 
	\sa_count[14].r.part0[25] , \sa_count[14].r.part0[24] , 
	\sa_count[14].r.part0[23] , \sa_count[14].r.part0[22] , 
	\sa_count[14].r.part0[21] , \sa_count[14].r.part0[20] , 
	\sa_count[14].r.part0[19] , \sa_count[14].r.part0[18] , 
	\sa_count[14].r.part0[17] , \sa_count[14].r.part0[16] , 
	\sa_count[14].r.part0[15] , \sa_count[14].r.part0[14] , 
	\sa_count[14].r.part0[13] , \sa_count[14].r.part0[12] , 
	\sa_count[14].r.part0[11] , \sa_count[14].r.part0[10] , 
	\sa_count[14].r.part0[9] , \sa_count[14].r.part0[8] , 
	\sa_count[14].r.part0[7] , \sa_count[14].r.part0[6] , 
	\sa_count[14].r.part0[5] , \sa_count[14].r.part0[4] , 
	\sa_count[14].r.part0[3] , \sa_count[14].r.part0[2] , 
	\sa_count[14].r.part0[1] , \sa_count[14].r.part0[0] , 
	\sa_count[13].r.part1[31] , \sa_count[13].r.part1[30] , 
	\sa_count[13].r.part1[29] , \sa_count[13].r.part1[28] , 
	\sa_count[13].r.part1[27] , \sa_count[13].r.part1[26] , 
	\sa_count[13].r.part1[25] , \sa_count[13].r.part1[24] , 
	\sa_count[13].r.part1[23] , \sa_count[13].r.part1[22] , 
	\sa_count[13].r.part1[21] , \sa_count[13].r.part1[20] , 
	\sa_count[13].r.part1[19] , \sa_count[13].r.part1[18] , 
	\sa_count[13].r.part1[17] , \sa_count[13].r.part1[16] , 
	\sa_count[13].r.part1[15] , \sa_count[13].r.part1[14] , 
	\sa_count[13].r.part1[13] , \sa_count[13].r.part1[12] , 
	\sa_count[13].r.part1[11] , \sa_count[13].r.part1[10] , 
	\sa_count[13].r.part1[9] , \sa_count[13].r.part1[8] , 
	\sa_count[13].r.part1[7] , \sa_count[13].r.part1[6] , 
	\sa_count[13].r.part1[5] , \sa_count[13].r.part1[4] , 
	\sa_count[13].r.part1[3] , \sa_count[13].r.part1[2] , 
	\sa_count[13].r.part1[1] , \sa_count[13].r.part1[0] , 
	\sa_count[13].r.part0[31] , \sa_count[13].r.part0[30] , 
	\sa_count[13].r.part0[29] , \sa_count[13].r.part0[28] , 
	\sa_count[13].r.part0[27] , \sa_count[13].r.part0[26] , 
	\sa_count[13].r.part0[25] , \sa_count[13].r.part0[24] , 
	\sa_count[13].r.part0[23] , \sa_count[13].r.part0[22] , 
	\sa_count[13].r.part0[21] , \sa_count[13].r.part0[20] , 
	\sa_count[13].r.part0[19] , \sa_count[13].r.part0[18] , 
	\sa_count[13].r.part0[17] , \sa_count[13].r.part0[16] , 
	\sa_count[13].r.part0[15] , \sa_count[13].r.part0[14] , 
	\sa_count[13].r.part0[13] , \sa_count[13].r.part0[12] , 
	\sa_count[13].r.part0[11] , \sa_count[13].r.part0[10] , 
	\sa_count[13].r.part0[9] , \sa_count[13].r.part0[8] , 
	\sa_count[13].r.part0[7] , \sa_count[13].r.part0[6] , 
	\sa_count[13].r.part0[5] , \sa_count[13].r.part0[4] , 
	\sa_count[13].r.part0[3] , \sa_count[13].r.part0[2] , 
	\sa_count[13].r.part0[1] , \sa_count[13].r.part0[0] , 
	\sa_count[12].r.part1[31] , \sa_count[12].r.part1[30] , 
	\sa_count[12].r.part1[29] , \sa_count[12].r.part1[28] , 
	\sa_count[12].r.part1[27] , \sa_count[12].r.part1[26] , 
	\sa_count[12].r.part1[25] , \sa_count[12].r.part1[24] , 
	\sa_count[12].r.part1[23] , \sa_count[12].r.part1[22] , 
	\sa_count[12].r.part1[21] , \sa_count[12].r.part1[20] , 
	\sa_count[12].r.part1[19] , \sa_count[12].r.part1[18] , 
	\sa_count[12].r.part1[17] , \sa_count[12].r.part1[16] , 
	\sa_count[12].r.part1[15] , \sa_count[12].r.part1[14] , 
	\sa_count[12].r.part1[13] , \sa_count[12].r.part1[12] , 
	\sa_count[12].r.part1[11] , \sa_count[12].r.part1[10] , 
	\sa_count[12].r.part1[9] , \sa_count[12].r.part1[8] , 
	\sa_count[12].r.part1[7] , \sa_count[12].r.part1[6] , 
	\sa_count[12].r.part1[5] , \sa_count[12].r.part1[4] , 
	\sa_count[12].r.part1[3] , \sa_count[12].r.part1[2] , 
	\sa_count[12].r.part1[1] , \sa_count[12].r.part1[0] , 
	\sa_count[12].r.part0[31] , \sa_count[12].r.part0[30] , 
	\sa_count[12].r.part0[29] , \sa_count[12].r.part0[28] , 
	\sa_count[12].r.part0[27] , \sa_count[12].r.part0[26] , 
	\sa_count[12].r.part0[25] , \sa_count[12].r.part0[24] , 
	\sa_count[12].r.part0[23] , \sa_count[12].r.part0[22] , 
	\sa_count[12].r.part0[21] , \sa_count[12].r.part0[20] , 
	\sa_count[12].r.part0[19] , \sa_count[12].r.part0[18] , 
	\sa_count[12].r.part0[17] , \sa_count[12].r.part0[16] , 
	\sa_count[12].r.part0[15] , \sa_count[12].r.part0[14] , 
	\sa_count[12].r.part0[13] , \sa_count[12].r.part0[12] , 
	\sa_count[12].r.part0[11] , \sa_count[12].r.part0[10] , 
	\sa_count[12].r.part0[9] , \sa_count[12].r.part0[8] , 
	\sa_count[12].r.part0[7] , \sa_count[12].r.part0[6] , 
	\sa_count[12].r.part0[5] , \sa_count[12].r.part0[4] , 
	\sa_count[12].r.part0[3] , \sa_count[12].r.part0[2] , 
	\sa_count[12].r.part0[1] , \sa_count[12].r.part0[0] , 
	\sa_count[11].r.part1[31] , \sa_count[11].r.part1[30] , 
	\sa_count[11].r.part1[29] , \sa_count[11].r.part1[28] , 
	\sa_count[11].r.part1[27] , \sa_count[11].r.part1[26] , 
	\sa_count[11].r.part1[25] , \sa_count[11].r.part1[24] , 
	\sa_count[11].r.part1[23] , \sa_count[11].r.part1[22] , 
	\sa_count[11].r.part1[21] , \sa_count[11].r.part1[20] , 
	\sa_count[11].r.part1[19] , \sa_count[11].r.part1[18] , 
	\sa_count[11].r.part1[17] , \sa_count[11].r.part1[16] , 
	\sa_count[11].r.part1[15] , \sa_count[11].r.part1[14] , 
	\sa_count[11].r.part1[13] , \sa_count[11].r.part1[12] , 
	\sa_count[11].r.part1[11] , \sa_count[11].r.part1[10] , 
	\sa_count[11].r.part1[9] , \sa_count[11].r.part1[8] , 
	\sa_count[11].r.part1[7] , \sa_count[11].r.part1[6] , 
	\sa_count[11].r.part1[5] , \sa_count[11].r.part1[4] , 
	\sa_count[11].r.part1[3] , \sa_count[11].r.part1[2] , 
	\sa_count[11].r.part1[1] , \sa_count[11].r.part1[0] , 
	\sa_count[11].r.part0[31] , \sa_count[11].r.part0[30] , 
	\sa_count[11].r.part0[29] , \sa_count[11].r.part0[28] , 
	\sa_count[11].r.part0[27] , \sa_count[11].r.part0[26] , 
	\sa_count[11].r.part0[25] , \sa_count[11].r.part0[24] , 
	\sa_count[11].r.part0[23] , \sa_count[11].r.part0[22] , 
	\sa_count[11].r.part0[21] , \sa_count[11].r.part0[20] , 
	\sa_count[11].r.part0[19] , \sa_count[11].r.part0[18] , 
	\sa_count[11].r.part0[17] , \sa_count[11].r.part0[16] , 
	\sa_count[11].r.part0[15] , \sa_count[11].r.part0[14] , 
	\sa_count[11].r.part0[13] , \sa_count[11].r.part0[12] , 
	\sa_count[11].r.part0[11] , \sa_count[11].r.part0[10] , 
	\sa_count[11].r.part0[9] , \sa_count[11].r.part0[8] , 
	\sa_count[11].r.part0[7] , \sa_count[11].r.part0[6] , 
	\sa_count[11].r.part0[5] , \sa_count[11].r.part0[4] , 
	\sa_count[11].r.part0[3] , \sa_count[11].r.part0[2] , 
	\sa_count[11].r.part0[1] , \sa_count[11].r.part0[0] , 
	\sa_count[10].r.part1[31] , \sa_count[10].r.part1[30] , 
	\sa_count[10].r.part1[29] , \sa_count[10].r.part1[28] , 
	\sa_count[10].r.part1[27] , \sa_count[10].r.part1[26] , 
	\sa_count[10].r.part1[25] , \sa_count[10].r.part1[24] , 
	\sa_count[10].r.part1[23] , \sa_count[10].r.part1[22] , 
	\sa_count[10].r.part1[21] , \sa_count[10].r.part1[20] , 
	\sa_count[10].r.part1[19] , \sa_count[10].r.part1[18] , 
	\sa_count[10].r.part1[17] , \sa_count[10].r.part1[16] , 
	\sa_count[10].r.part1[15] , \sa_count[10].r.part1[14] , 
	\sa_count[10].r.part1[13] , \sa_count[10].r.part1[12] , 
	\sa_count[10].r.part1[11] , \sa_count[10].r.part1[10] , 
	\sa_count[10].r.part1[9] , \sa_count[10].r.part1[8] , 
	\sa_count[10].r.part1[7] , \sa_count[10].r.part1[6] , 
	\sa_count[10].r.part1[5] , \sa_count[10].r.part1[4] , 
	\sa_count[10].r.part1[3] , \sa_count[10].r.part1[2] , 
	\sa_count[10].r.part1[1] , \sa_count[10].r.part1[0] , 
	\sa_count[10].r.part0[31] , \sa_count[10].r.part0[30] , 
	\sa_count[10].r.part0[29] , \sa_count[10].r.part0[28] , 
	\sa_count[10].r.part0[27] , \sa_count[10].r.part0[26] , 
	\sa_count[10].r.part0[25] , \sa_count[10].r.part0[24] , 
	\sa_count[10].r.part0[23] , \sa_count[10].r.part0[22] , 
	\sa_count[10].r.part0[21] , \sa_count[10].r.part0[20] , 
	\sa_count[10].r.part0[19] , \sa_count[10].r.part0[18] , 
	\sa_count[10].r.part0[17] , \sa_count[10].r.part0[16] , 
	\sa_count[10].r.part0[15] , \sa_count[10].r.part0[14] , 
	\sa_count[10].r.part0[13] , \sa_count[10].r.part0[12] , 
	\sa_count[10].r.part0[11] , \sa_count[10].r.part0[10] , 
	\sa_count[10].r.part0[9] , \sa_count[10].r.part0[8] , 
	\sa_count[10].r.part0[7] , \sa_count[10].r.part0[6] , 
	\sa_count[10].r.part0[5] , \sa_count[10].r.part0[4] , 
	\sa_count[10].r.part0[3] , \sa_count[10].r.part0[2] , 
	\sa_count[10].r.part0[1] , \sa_count[10].r.part0[0] , 
	\sa_count[9].r.part1[31] , \sa_count[9].r.part1[30] , 
	\sa_count[9].r.part1[29] , \sa_count[9].r.part1[28] , 
	\sa_count[9].r.part1[27] , \sa_count[9].r.part1[26] , 
	\sa_count[9].r.part1[25] , \sa_count[9].r.part1[24] , 
	\sa_count[9].r.part1[23] , \sa_count[9].r.part1[22] , 
	\sa_count[9].r.part1[21] , \sa_count[9].r.part1[20] , 
	\sa_count[9].r.part1[19] , \sa_count[9].r.part1[18] , 
	\sa_count[9].r.part1[17] , \sa_count[9].r.part1[16] , 
	\sa_count[9].r.part1[15] , \sa_count[9].r.part1[14] , 
	\sa_count[9].r.part1[13] , \sa_count[9].r.part1[12] , 
	\sa_count[9].r.part1[11] , \sa_count[9].r.part1[10] , 
	\sa_count[9].r.part1[9] , \sa_count[9].r.part1[8] , 
	\sa_count[9].r.part1[7] , \sa_count[9].r.part1[6] , 
	\sa_count[9].r.part1[5] , \sa_count[9].r.part1[4] , 
	\sa_count[9].r.part1[3] , \sa_count[9].r.part1[2] , 
	\sa_count[9].r.part1[1] , \sa_count[9].r.part1[0] , 
	\sa_count[9].r.part0[31] , \sa_count[9].r.part0[30] , 
	\sa_count[9].r.part0[29] , \sa_count[9].r.part0[28] , 
	\sa_count[9].r.part0[27] , \sa_count[9].r.part0[26] , 
	\sa_count[9].r.part0[25] , \sa_count[9].r.part0[24] , 
	\sa_count[9].r.part0[23] , \sa_count[9].r.part0[22] , 
	\sa_count[9].r.part0[21] , \sa_count[9].r.part0[20] , 
	\sa_count[9].r.part0[19] , \sa_count[9].r.part0[18] , 
	\sa_count[9].r.part0[17] , \sa_count[9].r.part0[16] , 
	\sa_count[9].r.part0[15] , \sa_count[9].r.part0[14] , 
	\sa_count[9].r.part0[13] , \sa_count[9].r.part0[12] , 
	\sa_count[9].r.part0[11] , \sa_count[9].r.part0[10] , 
	\sa_count[9].r.part0[9] , \sa_count[9].r.part0[8] , 
	\sa_count[9].r.part0[7] , \sa_count[9].r.part0[6] , 
	\sa_count[9].r.part0[5] , \sa_count[9].r.part0[4] , 
	\sa_count[9].r.part0[3] , \sa_count[9].r.part0[2] , 
	\sa_count[9].r.part0[1] , \sa_count[9].r.part0[0] , 
	\sa_count[8].r.part1[31] , \sa_count[8].r.part1[30] , 
	\sa_count[8].r.part1[29] , \sa_count[8].r.part1[28] , 
	\sa_count[8].r.part1[27] , \sa_count[8].r.part1[26] , 
	\sa_count[8].r.part1[25] , \sa_count[8].r.part1[24] , 
	\sa_count[8].r.part1[23] , \sa_count[8].r.part1[22] , 
	\sa_count[8].r.part1[21] , \sa_count[8].r.part1[20] , 
	\sa_count[8].r.part1[19] , \sa_count[8].r.part1[18] , 
	\sa_count[8].r.part1[17] , \sa_count[8].r.part1[16] , 
	\sa_count[8].r.part1[15] , \sa_count[8].r.part1[14] , 
	\sa_count[8].r.part1[13] , \sa_count[8].r.part1[12] , 
	\sa_count[8].r.part1[11] , \sa_count[8].r.part1[10] , 
	\sa_count[8].r.part1[9] , \sa_count[8].r.part1[8] , 
	\sa_count[8].r.part1[7] , \sa_count[8].r.part1[6] , 
	\sa_count[8].r.part1[5] , \sa_count[8].r.part1[4] , 
	\sa_count[8].r.part1[3] , \sa_count[8].r.part1[2] , 
	\sa_count[8].r.part1[1] , \sa_count[8].r.part1[0] , 
	\sa_count[8].r.part0[31] , \sa_count[8].r.part0[30] , 
	\sa_count[8].r.part0[29] , \sa_count[8].r.part0[28] , 
	\sa_count[8].r.part0[27] , \sa_count[8].r.part0[26] , 
	\sa_count[8].r.part0[25] , \sa_count[8].r.part0[24] , 
	\sa_count[8].r.part0[23] , \sa_count[8].r.part0[22] , 
	\sa_count[8].r.part0[21] , \sa_count[8].r.part0[20] , 
	\sa_count[8].r.part0[19] , \sa_count[8].r.part0[18] , 
	\sa_count[8].r.part0[17] , \sa_count[8].r.part0[16] , 
	\sa_count[8].r.part0[15] , \sa_count[8].r.part0[14] , 
	\sa_count[8].r.part0[13] , \sa_count[8].r.part0[12] , 
	\sa_count[8].r.part0[11] , \sa_count[8].r.part0[10] , 
	\sa_count[8].r.part0[9] , \sa_count[8].r.part0[8] , 
	\sa_count[8].r.part0[7] , \sa_count[8].r.part0[6] , 
	\sa_count[8].r.part0[5] , \sa_count[8].r.part0[4] , 
	\sa_count[8].r.part0[3] , \sa_count[8].r.part0[2] , 
	\sa_count[8].r.part0[1] , \sa_count[8].r.part0[0] , 
	\sa_count[7].r.part1[31] , \sa_count[7].r.part1[30] , 
	\sa_count[7].r.part1[29] , \sa_count[7].r.part1[28] , 
	\sa_count[7].r.part1[27] , \sa_count[7].r.part1[26] , 
	\sa_count[7].r.part1[25] , \sa_count[7].r.part1[24] , 
	\sa_count[7].r.part1[23] , \sa_count[7].r.part1[22] , 
	\sa_count[7].r.part1[21] , \sa_count[7].r.part1[20] , 
	\sa_count[7].r.part1[19] , \sa_count[7].r.part1[18] , 
	\sa_count[7].r.part1[17] , \sa_count[7].r.part1[16] , 
	\sa_count[7].r.part1[15] , \sa_count[7].r.part1[14] , 
	\sa_count[7].r.part1[13] , \sa_count[7].r.part1[12] , 
	\sa_count[7].r.part1[11] , \sa_count[7].r.part1[10] , 
	\sa_count[7].r.part1[9] , \sa_count[7].r.part1[8] , 
	\sa_count[7].r.part1[7] , \sa_count[7].r.part1[6] , 
	\sa_count[7].r.part1[5] , \sa_count[7].r.part1[4] , 
	\sa_count[7].r.part1[3] , \sa_count[7].r.part1[2] , 
	\sa_count[7].r.part1[1] , \sa_count[7].r.part1[0] , 
	\sa_count[7].r.part0[31] , \sa_count[7].r.part0[30] , 
	\sa_count[7].r.part0[29] , \sa_count[7].r.part0[28] , 
	\sa_count[7].r.part0[27] , \sa_count[7].r.part0[26] , 
	\sa_count[7].r.part0[25] , \sa_count[7].r.part0[24] , 
	\sa_count[7].r.part0[23] , \sa_count[7].r.part0[22] , 
	\sa_count[7].r.part0[21] , \sa_count[7].r.part0[20] , 
	\sa_count[7].r.part0[19] , \sa_count[7].r.part0[18] , 
	\sa_count[7].r.part0[17] , \sa_count[7].r.part0[16] , 
	\sa_count[7].r.part0[15] , \sa_count[7].r.part0[14] , 
	\sa_count[7].r.part0[13] , \sa_count[7].r.part0[12] , 
	\sa_count[7].r.part0[11] , \sa_count[7].r.part0[10] , 
	\sa_count[7].r.part0[9] , \sa_count[7].r.part0[8] , 
	\sa_count[7].r.part0[7] , \sa_count[7].r.part0[6] , 
	\sa_count[7].r.part0[5] , \sa_count[7].r.part0[4] , 
	\sa_count[7].r.part0[3] , \sa_count[7].r.part0[2] , 
	\sa_count[7].r.part0[1] , \sa_count[7].r.part0[0] , 
	\sa_count[6].r.part1[31] , \sa_count[6].r.part1[30] , 
	\sa_count[6].r.part1[29] , \sa_count[6].r.part1[28] , 
	\sa_count[6].r.part1[27] , \sa_count[6].r.part1[26] , 
	\sa_count[6].r.part1[25] , \sa_count[6].r.part1[24] , 
	\sa_count[6].r.part1[23] , \sa_count[6].r.part1[22] , 
	\sa_count[6].r.part1[21] , \sa_count[6].r.part1[20] , 
	\sa_count[6].r.part1[19] , \sa_count[6].r.part1[18] , 
	\sa_count[6].r.part1[17] , \sa_count[6].r.part1[16] , 
	\sa_count[6].r.part1[15] , \sa_count[6].r.part1[14] , 
	\sa_count[6].r.part1[13] , \sa_count[6].r.part1[12] , 
	\sa_count[6].r.part1[11] , \sa_count[6].r.part1[10] , 
	\sa_count[6].r.part1[9] , \sa_count[6].r.part1[8] , 
	\sa_count[6].r.part1[7] , \sa_count[6].r.part1[6] , 
	\sa_count[6].r.part1[5] , \sa_count[6].r.part1[4] , 
	\sa_count[6].r.part1[3] , \sa_count[6].r.part1[2] , 
	\sa_count[6].r.part1[1] , \sa_count[6].r.part1[0] , 
	\sa_count[6].r.part0[31] , \sa_count[6].r.part0[30] , 
	\sa_count[6].r.part0[29] , \sa_count[6].r.part0[28] , 
	\sa_count[6].r.part0[27] , \sa_count[6].r.part0[26] , 
	\sa_count[6].r.part0[25] , \sa_count[6].r.part0[24] , 
	\sa_count[6].r.part0[23] , \sa_count[6].r.part0[22] , 
	\sa_count[6].r.part0[21] , \sa_count[6].r.part0[20] , 
	\sa_count[6].r.part0[19] , \sa_count[6].r.part0[18] , 
	\sa_count[6].r.part0[17] , \sa_count[6].r.part0[16] , 
	\sa_count[6].r.part0[15] , \sa_count[6].r.part0[14] , 
	\sa_count[6].r.part0[13] , \sa_count[6].r.part0[12] , 
	\sa_count[6].r.part0[11] , \sa_count[6].r.part0[10] , 
	\sa_count[6].r.part0[9] , \sa_count[6].r.part0[8] , 
	\sa_count[6].r.part0[7] , \sa_count[6].r.part0[6] , 
	\sa_count[6].r.part0[5] , \sa_count[6].r.part0[4] , 
	\sa_count[6].r.part0[3] , \sa_count[6].r.part0[2] , 
	\sa_count[6].r.part0[1] , \sa_count[6].r.part0[0] , 
	\sa_count[5].r.part1[31] , \sa_count[5].r.part1[30] , 
	\sa_count[5].r.part1[29] , \sa_count[5].r.part1[28] , 
	\sa_count[5].r.part1[27] , \sa_count[5].r.part1[26] , 
	\sa_count[5].r.part1[25] , \sa_count[5].r.part1[24] , 
	\sa_count[5].r.part1[23] , \sa_count[5].r.part1[22] , 
	\sa_count[5].r.part1[21] , \sa_count[5].r.part1[20] , 
	\sa_count[5].r.part1[19] , \sa_count[5].r.part1[18] , 
	\sa_count[5].r.part1[17] , \sa_count[5].r.part1[16] , 
	\sa_count[5].r.part1[15] , \sa_count[5].r.part1[14] , 
	\sa_count[5].r.part1[13] , \sa_count[5].r.part1[12] , 
	\sa_count[5].r.part1[11] , \sa_count[5].r.part1[10] , 
	\sa_count[5].r.part1[9] , \sa_count[5].r.part1[8] , 
	\sa_count[5].r.part1[7] , \sa_count[5].r.part1[6] , 
	\sa_count[5].r.part1[5] , \sa_count[5].r.part1[4] , 
	\sa_count[5].r.part1[3] , \sa_count[5].r.part1[2] , 
	\sa_count[5].r.part1[1] , \sa_count[5].r.part1[0] , 
	\sa_count[5].r.part0[31] , \sa_count[5].r.part0[30] , 
	\sa_count[5].r.part0[29] , \sa_count[5].r.part0[28] , 
	\sa_count[5].r.part0[27] , \sa_count[5].r.part0[26] , 
	\sa_count[5].r.part0[25] , \sa_count[5].r.part0[24] , 
	\sa_count[5].r.part0[23] , \sa_count[5].r.part0[22] , 
	\sa_count[5].r.part0[21] , \sa_count[5].r.part0[20] , 
	\sa_count[5].r.part0[19] , \sa_count[5].r.part0[18] , 
	\sa_count[5].r.part0[17] , \sa_count[5].r.part0[16] , 
	\sa_count[5].r.part0[15] , \sa_count[5].r.part0[14] , 
	\sa_count[5].r.part0[13] , \sa_count[5].r.part0[12] , 
	\sa_count[5].r.part0[11] , \sa_count[5].r.part0[10] , 
	\sa_count[5].r.part0[9] , \sa_count[5].r.part0[8] , 
	\sa_count[5].r.part0[7] , \sa_count[5].r.part0[6] , 
	\sa_count[5].r.part0[5] , \sa_count[5].r.part0[4] , 
	\sa_count[5].r.part0[3] , \sa_count[5].r.part0[2] , 
	\sa_count[5].r.part0[1] , \sa_count[5].r.part0[0] , 
	\sa_count[4].r.part1[31] , \sa_count[4].r.part1[30] , 
	\sa_count[4].r.part1[29] , \sa_count[4].r.part1[28] , 
	\sa_count[4].r.part1[27] , \sa_count[4].r.part1[26] , 
	\sa_count[4].r.part1[25] , \sa_count[4].r.part1[24] , 
	\sa_count[4].r.part1[23] , \sa_count[4].r.part1[22] , 
	\sa_count[4].r.part1[21] , \sa_count[4].r.part1[20] , 
	\sa_count[4].r.part1[19] , \sa_count[4].r.part1[18] , 
	\sa_count[4].r.part1[17] , \sa_count[4].r.part1[16] , 
	\sa_count[4].r.part1[15] , \sa_count[4].r.part1[14] , 
	\sa_count[4].r.part1[13] , \sa_count[4].r.part1[12] , 
	\sa_count[4].r.part1[11] , \sa_count[4].r.part1[10] , 
	\sa_count[4].r.part1[9] , \sa_count[4].r.part1[8] , 
	\sa_count[4].r.part1[7] , \sa_count[4].r.part1[6] , 
	\sa_count[4].r.part1[5] , \sa_count[4].r.part1[4] , 
	\sa_count[4].r.part1[3] , \sa_count[4].r.part1[2] , 
	\sa_count[4].r.part1[1] , \sa_count[4].r.part1[0] , 
	\sa_count[4].r.part0[31] , \sa_count[4].r.part0[30] , 
	\sa_count[4].r.part0[29] , \sa_count[4].r.part0[28] , 
	\sa_count[4].r.part0[27] , \sa_count[4].r.part0[26] , 
	\sa_count[4].r.part0[25] , \sa_count[4].r.part0[24] , 
	\sa_count[4].r.part0[23] , \sa_count[4].r.part0[22] , 
	\sa_count[4].r.part0[21] , \sa_count[4].r.part0[20] , 
	\sa_count[4].r.part0[19] , \sa_count[4].r.part0[18] , 
	\sa_count[4].r.part0[17] , \sa_count[4].r.part0[16] , 
	\sa_count[4].r.part0[15] , \sa_count[4].r.part0[14] , 
	\sa_count[4].r.part0[13] , \sa_count[4].r.part0[12] , 
	\sa_count[4].r.part0[11] , \sa_count[4].r.part0[10] , 
	\sa_count[4].r.part0[9] , \sa_count[4].r.part0[8] , 
	\sa_count[4].r.part0[7] , \sa_count[4].r.part0[6] , 
	\sa_count[4].r.part0[5] , \sa_count[4].r.part0[4] , 
	\sa_count[4].r.part0[3] , \sa_count[4].r.part0[2] , 
	\sa_count[4].r.part0[1] , \sa_count[4].r.part0[0] , 
	\sa_count[3].r.part1[31] , \sa_count[3].r.part1[30] , 
	\sa_count[3].r.part1[29] , \sa_count[3].r.part1[28] , 
	\sa_count[3].r.part1[27] , \sa_count[3].r.part1[26] , 
	\sa_count[3].r.part1[25] , \sa_count[3].r.part1[24] , 
	\sa_count[3].r.part1[23] , \sa_count[3].r.part1[22] , 
	\sa_count[3].r.part1[21] , \sa_count[3].r.part1[20] , 
	\sa_count[3].r.part1[19] , \sa_count[3].r.part1[18] , 
	\sa_count[3].r.part1[17] , \sa_count[3].r.part1[16] , 
	\sa_count[3].r.part1[15] , \sa_count[3].r.part1[14] , 
	\sa_count[3].r.part1[13] , \sa_count[3].r.part1[12] , 
	\sa_count[3].r.part1[11] , \sa_count[3].r.part1[10] , 
	\sa_count[3].r.part1[9] , \sa_count[3].r.part1[8] , 
	\sa_count[3].r.part1[7] , \sa_count[3].r.part1[6] , 
	\sa_count[3].r.part1[5] , \sa_count[3].r.part1[4] , 
	\sa_count[3].r.part1[3] , \sa_count[3].r.part1[2] , 
	\sa_count[3].r.part1[1] , \sa_count[3].r.part1[0] , 
	\sa_count[3].r.part0[31] , \sa_count[3].r.part0[30] , 
	\sa_count[3].r.part0[29] , \sa_count[3].r.part0[28] , 
	\sa_count[3].r.part0[27] , \sa_count[3].r.part0[26] , 
	\sa_count[3].r.part0[25] , \sa_count[3].r.part0[24] , 
	\sa_count[3].r.part0[23] , \sa_count[3].r.part0[22] , 
	\sa_count[3].r.part0[21] , \sa_count[3].r.part0[20] , 
	\sa_count[3].r.part0[19] , \sa_count[3].r.part0[18] , 
	\sa_count[3].r.part0[17] , \sa_count[3].r.part0[16] , 
	\sa_count[3].r.part0[15] , \sa_count[3].r.part0[14] , 
	\sa_count[3].r.part0[13] , \sa_count[3].r.part0[12] , 
	\sa_count[3].r.part0[11] , \sa_count[3].r.part0[10] , 
	\sa_count[3].r.part0[9] , \sa_count[3].r.part0[8] , 
	\sa_count[3].r.part0[7] , \sa_count[3].r.part0[6] , 
	\sa_count[3].r.part0[5] , \sa_count[3].r.part0[4] , 
	\sa_count[3].r.part0[3] , \sa_count[3].r.part0[2] , 
	\sa_count[3].r.part0[1] , \sa_count[3].r.part0[0] , 
	\sa_count[2].r.part1[31] , \sa_count[2].r.part1[30] , 
	\sa_count[2].r.part1[29] , \sa_count[2].r.part1[28] , 
	\sa_count[2].r.part1[27] , \sa_count[2].r.part1[26] , 
	\sa_count[2].r.part1[25] , \sa_count[2].r.part1[24] , 
	\sa_count[2].r.part1[23] , \sa_count[2].r.part1[22] , 
	\sa_count[2].r.part1[21] , \sa_count[2].r.part1[20] , 
	\sa_count[2].r.part1[19] , \sa_count[2].r.part1[18] , 
	\sa_count[2].r.part1[17] , \sa_count[2].r.part1[16] , 
	\sa_count[2].r.part1[15] , \sa_count[2].r.part1[14] , 
	\sa_count[2].r.part1[13] , \sa_count[2].r.part1[12] , 
	\sa_count[2].r.part1[11] , \sa_count[2].r.part1[10] , 
	\sa_count[2].r.part1[9] , \sa_count[2].r.part1[8] , 
	\sa_count[2].r.part1[7] , \sa_count[2].r.part1[6] , 
	\sa_count[2].r.part1[5] , \sa_count[2].r.part1[4] , 
	\sa_count[2].r.part1[3] , \sa_count[2].r.part1[2] , 
	\sa_count[2].r.part1[1] , \sa_count[2].r.part1[0] , 
	\sa_count[2].r.part0[31] , \sa_count[2].r.part0[30] , 
	\sa_count[2].r.part0[29] , \sa_count[2].r.part0[28] , 
	\sa_count[2].r.part0[27] , \sa_count[2].r.part0[26] , 
	\sa_count[2].r.part0[25] , \sa_count[2].r.part0[24] , 
	\sa_count[2].r.part0[23] , \sa_count[2].r.part0[22] , 
	\sa_count[2].r.part0[21] , \sa_count[2].r.part0[20] , 
	\sa_count[2].r.part0[19] , \sa_count[2].r.part0[18] , 
	\sa_count[2].r.part0[17] , \sa_count[2].r.part0[16] , 
	\sa_count[2].r.part0[15] , \sa_count[2].r.part0[14] , 
	\sa_count[2].r.part0[13] , \sa_count[2].r.part0[12] , 
	\sa_count[2].r.part0[11] , \sa_count[2].r.part0[10] , 
	\sa_count[2].r.part0[9] , \sa_count[2].r.part0[8] , 
	\sa_count[2].r.part0[7] , \sa_count[2].r.part0[6] , 
	\sa_count[2].r.part0[5] , \sa_count[2].r.part0[4] , 
	\sa_count[2].r.part0[3] , \sa_count[2].r.part0[2] , 
	\sa_count[2].r.part0[1] , \sa_count[2].r.part0[0] , 
	\sa_count[1].r.part1[31] , \sa_count[1].r.part1[30] , 
	\sa_count[1].r.part1[29] , \sa_count[1].r.part1[28] , 
	\sa_count[1].r.part1[27] , \sa_count[1].r.part1[26] , 
	\sa_count[1].r.part1[25] , \sa_count[1].r.part1[24] , 
	\sa_count[1].r.part1[23] , \sa_count[1].r.part1[22] , 
	\sa_count[1].r.part1[21] , \sa_count[1].r.part1[20] , 
	\sa_count[1].r.part1[19] , \sa_count[1].r.part1[18] , 
	\sa_count[1].r.part1[17] , \sa_count[1].r.part1[16] , 
	\sa_count[1].r.part1[15] , \sa_count[1].r.part1[14] , 
	\sa_count[1].r.part1[13] , \sa_count[1].r.part1[12] , 
	\sa_count[1].r.part1[11] , \sa_count[1].r.part1[10] , 
	\sa_count[1].r.part1[9] , \sa_count[1].r.part1[8] , 
	\sa_count[1].r.part1[7] , \sa_count[1].r.part1[6] , 
	\sa_count[1].r.part1[5] , \sa_count[1].r.part1[4] , 
	\sa_count[1].r.part1[3] , \sa_count[1].r.part1[2] , 
	\sa_count[1].r.part1[1] , \sa_count[1].r.part1[0] , 
	\sa_count[1].r.part0[31] , \sa_count[1].r.part0[30] , 
	\sa_count[1].r.part0[29] , \sa_count[1].r.part0[28] , 
	\sa_count[1].r.part0[27] , \sa_count[1].r.part0[26] , 
	\sa_count[1].r.part0[25] , \sa_count[1].r.part0[24] , 
	\sa_count[1].r.part0[23] , \sa_count[1].r.part0[22] , 
	\sa_count[1].r.part0[21] , \sa_count[1].r.part0[20] , 
	\sa_count[1].r.part0[19] , \sa_count[1].r.part0[18] , 
	\sa_count[1].r.part0[17] , \sa_count[1].r.part0[16] , 
	\sa_count[1].r.part0[15] , \sa_count[1].r.part0[14] , 
	\sa_count[1].r.part0[13] , \sa_count[1].r.part0[12] , 
	\sa_count[1].r.part0[11] , \sa_count[1].r.part0[10] , 
	\sa_count[1].r.part0[9] , \sa_count[1].r.part0[8] , 
	\sa_count[1].r.part0[7] , \sa_count[1].r.part0[6] , 
	\sa_count[1].r.part0[5] , \sa_count[1].r.part0[4] , 
	\sa_count[1].r.part0[3] , \sa_count[1].r.part0[2] , 
	\sa_count[1].r.part0[1] , \sa_count[1].r.part0[0] , 
	\sa_count[0].r.part1[31] , \sa_count[0].r.part1[30] , 
	\sa_count[0].r.part1[29] , \sa_count[0].r.part1[28] , 
	\sa_count[0].r.part1[27] , \sa_count[0].r.part1[26] , 
	\sa_count[0].r.part1[25] , \sa_count[0].r.part1[24] , 
	\sa_count[0].r.part1[23] , \sa_count[0].r.part1[22] , 
	\sa_count[0].r.part1[21] , \sa_count[0].r.part1[20] , 
	\sa_count[0].r.part1[19] , \sa_count[0].r.part1[18] , 
	\sa_count[0].r.part1[17] , \sa_count[0].r.part1[16] , 
	\sa_count[0].r.part1[15] , \sa_count[0].r.part1[14] , 
	\sa_count[0].r.part1[13] , \sa_count[0].r.part1[12] , 
	\sa_count[0].r.part1[11] , \sa_count[0].r.part1[10] , 
	\sa_count[0].r.part1[9] , \sa_count[0].r.part1[8] , 
	\sa_count[0].r.part1[7] , \sa_count[0].r.part1[6] , 
	\sa_count[0].r.part1[5] , \sa_count[0].r.part1[4] , 
	\sa_count[0].r.part1[3] , \sa_count[0].r.part1[2] , 
	\sa_count[0].r.part1[1] , \sa_count[0].r.part1[0] , 
	\sa_count[0].r.part0[31] , \sa_count[0].r.part0[30] , 
	\sa_count[0].r.part0[29] , \sa_count[0].r.part0[28] , 
	\sa_count[0].r.part0[27] , \sa_count[0].r.part0[26] , 
	\sa_count[0].r.part0[25] , \sa_count[0].r.part0[24] , 
	\sa_count[0].r.part0[23] , \sa_count[0].r.part0[22] , 
	\sa_count[0].r.part0[21] , \sa_count[0].r.part0[20] , 
	\sa_count[0].r.part0[19] , \sa_count[0].r.part0[18] , 
	\sa_count[0].r.part0[17] , \sa_count[0].r.part0[16] , 
	\sa_count[0].r.part0[15] , \sa_count[0].r.part0[14] , 
	\sa_count[0].r.part0[13] , \sa_count[0].r.part0[12] , 
	\sa_count[0].r.part0[11] , \sa_count[0].r.part0[10] , 
	\sa_count[0].r.part0[9] , \sa_count[0].r.part0[8] , 
	\sa_count[0].r.part0[7] , \sa_count[0].r.part0[6] , 
	\sa_count[0].r.part0[5] , \sa_count[0].r.part0[4] , 
	\sa_count[0].r.part0[3] , \sa_count[0].r.part0[2] , 
	\sa_count[0].r.part0[1] , \sa_count[0].r.part0[0] } ), 
	debug_kme_ib_tready);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output suppress_key_tlvs;
output kme_interrupt;
output [15:0] \rbus_ring_o.addr ;
output \rbus_ring_o.wr_strb ;
output [31:0] \rbus_ring_o.wr_data ;
output \rbus_ring_o.rd_strb ;
output [31:0] \rbus_ring_o.rd_data ;
output \rbus_ring_o.ack ;
output \rbus_ring_o.err_ack ;
wire [83:0] rbus_ring_o;
output \kme_cceip0_ob_out.tvalid ;
output \kme_cceip0_ob_out.tlast ;
output [0:0] \kme_cceip0_ob_out.tid ;
output [7:0] \kme_cceip0_ob_out.tstrb ;
output [7:0] \kme_cceip0_ob_out.tuser ;
output [63:0] \kme_cceip0_ob_out.tdata ;
wire [82:0] kme_cceip0_ob_out;
output \kme_cceip0_ob_in_mod.tready ;
wire [0:0] kme_cceip0_ob_in_mod;
output \kme_cceip1_ob_out.tvalid ;
output \kme_cceip1_ob_out.tlast ;
output [0:0] \kme_cceip1_ob_out.tid ;
output [7:0] \kme_cceip1_ob_out.tstrb ;
output [7:0] \kme_cceip1_ob_out.tuser ;
output [63:0] \kme_cceip1_ob_out.tdata ;
wire [82:0] kme_cceip1_ob_out;
output \kme_cceip1_ob_in_mod.tready ;
wire [0:0] kme_cceip1_ob_in_mod;
output \kme_cceip2_ob_out.tvalid ;
output \kme_cceip2_ob_out.tlast ;
output [0:0] \kme_cceip2_ob_out.tid ;
output [7:0] \kme_cceip2_ob_out.tstrb ;
output [7:0] \kme_cceip2_ob_out.tuser ;
output [63:0] \kme_cceip2_ob_out.tdata ;
wire [82:0] kme_cceip2_ob_out;
output \kme_cceip2_ob_in_mod.tready ;
wire [0:0] kme_cceip2_ob_in_mod;
output \kme_cceip3_ob_out.tvalid ;
output \kme_cceip3_ob_out.tlast ;
output [0:0] \kme_cceip3_ob_out.tid ;
output [7:0] \kme_cceip3_ob_out.tstrb ;
output [7:0] \kme_cceip3_ob_out.tuser ;
output [63:0] \kme_cceip3_ob_out.tdata ;
wire [82:0] kme_cceip3_ob_out;
output \kme_cceip3_ob_in_mod.tready ;
wire [0:0] kme_cceip3_ob_in_mod;
output \kme_cddip0_ob_out.tvalid ;
output \kme_cddip0_ob_out.tlast ;
output [0:0] \kme_cddip0_ob_out.tid ;
output [7:0] \kme_cddip0_ob_out.tstrb ;
output [7:0] \kme_cddip0_ob_out.tuser ;
output [63:0] \kme_cddip0_ob_out.tdata ;
wire [82:0] kme_cddip0_ob_out;
output \kme_cddip0_ob_in_mod.tready ;
wire [0:0] kme_cddip0_ob_in_mod;
output \kme_cddip1_ob_out.tvalid ;
output \kme_cddip1_ob_out.tlast ;
output [0:0] \kme_cddip1_ob_out.tid ;
output [7:0] \kme_cddip1_ob_out.tstrb ;
output [7:0] \kme_cddip1_ob_out.tuser ;
output [63:0] \kme_cddip1_ob_out.tdata ;
wire [82:0] kme_cddip1_ob_out;
output \kme_cddip1_ob_in_mod.tready ;
wire [0:0] kme_cddip1_ob_in_mod;
output \kme_cddip2_ob_out.tvalid ;
output \kme_cddip2_ob_out.tlast ;
output [0:0] \kme_cddip2_ob_out.tid ;
output [7:0] \kme_cddip2_ob_out.tstrb ;
output [7:0] \kme_cddip2_ob_out.tuser ;
output [63:0] \kme_cddip2_ob_out.tdata ;
wire [82:0] kme_cddip2_ob_out;
output \kme_cddip2_ob_in_mod.tready ;
wire [0:0] kme_cddip2_ob_in_mod;
output \kme_cddip3_ob_out.tvalid ;
output \kme_cddip3_ob_out.tlast ;
output [0:0] \kme_cddip3_ob_out.tid ;
output [7:0] \kme_cddip3_ob_out.tstrb ;
output [7:0] \kme_cddip3_ob_out.tuser ;
output [63:0] \kme_cddip3_ob_out.tdata ;
wire [82:0] kme_cddip3_ob_out;
output \kme_cddip3_ob_in_mod.tready ;
wire [0:0] kme_cddip3_ob_in_mod;
output [63:0] ckv_dout;
output ckv_mbe;
output [0:0] \kim_dout.valid ;
output [2:0] \kim_dout.label_index ;
output [1:0] \kim_dout.ckv_length ;
output [14:0] \kim_dout.ckv_pointer ;
output [3:0] \kim_dout.pf_num ;
output [11:0] \kim_dout.vf_num ;
output [0:0] \kim_dout.vf_valid ;
wire [37:0] kim_dout;
output kim_mbe;
output bimc_rst_n;
output cceip_encrypt_bimc_isync;
output cceip_encrypt_bimc_idat;
output cceip_validate_bimc_isync;
output cceip_validate_bimc_idat;
output cddip_decrypt_bimc_isync;
output cddip_decrypt_bimc_idat;
output axi_bimc_isync;
output axi_bimc_idat;
output \labels[7].guid_size[0] ,\labels[7].label_size[5] 
	,\labels[7].label_size[4] ,\labels[7].label_size[3] 
	,\labels[7].label_size[2] ,\labels[7].label_size[1] 
	,\labels[7].label_size[0] ,\labels[7].label[255] 
	,\labels[7].label[254] ,\labels[7].label[253] ,\labels[7].label[252] 
	,\labels[7].label[251] ,\labels[7].label[250] ,\labels[7].label[249] 
	,\labels[7].label[248] ,\labels[7].label[247] ,\labels[7].label[246] 
	,\labels[7].label[245] ,\labels[7].label[244] ,\labels[7].label[243] 
	,\labels[7].label[242] ,\labels[7].label[241] ,\labels[7].label[240] 
	,\labels[7].label[239] ,\labels[7].label[238] ,\labels[7].label[237] 
	,\labels[7].label[236] ,\labels[7].label[235] ,\labels[7].label[234] 
	,\labels[7].label[233] ,\labels[7].label[232] ,\labels[7].label[231] 
	,\labels[7].label[230] ,\labels[7].label[229] ,\labels[7].label[228] 
	,\labels[7].label[227] ,\labels[7].label[226] ,\labels[7].label[225] 
	,\labels[7].label[224] ,\labels[7].label[223] ,\labels[7].label[222] 
	,\labels[7].label[221] ,\labels[7].label[220] ,\labels[7].label[219] 
	,\labels[7].label[218] ,\labels[7].label[217] ,\labels[7].label[216] 
	,\labels[7].label[215] ,\labels[7].label[214] ,\labels[7].label[213] 
	,\labels[7].label[212] ,\labels[7].label[211] ,\labels[7].label[210] 
	,\labels[7].label[209] ,\labels[7].label[208] ,\labels[7].label[207] 
	,\labels[7].label[206] ,\labels[7].label[205] ,\labels[7].label[204] 
	,\labels[7].label[203] ,\labels[7].label[202] ,\labels[7].label[201] 
	,\labels[7].label[200] ,\labels[7].label[199] ,\labels[7].label[198] 
	,\labels[7].label[197] ,\labels[7].label[196] ,\labels[7].label[195] 
	,\labels[7].label[194] ,\labels[7].label[193] ,\labels[7].label[192] 
	,\labels[7].label[191] ,\labels[7].label[190] ,\labels[7].label[189] 
	,\labels[7].label[188] ,\labels[7].label[187] ,\labels[7].label[186] 
	,\labels[7].label[185] ,\labels[7].label[184] ,\labels[7].label[183] 
	,\labels[7].label[182] ,\labels[7].label[181] ,\labels[7].label[180] 
	,\labels[7].label[179] ,\labels[7].label[178] ,\labels[7].label[177] 
	,\labels[7].label[176] ,\labels[7].label[175] ,\labels[7].label[174] 
	,\labels[7].label[173] ,\labels[7].label[172] ,\labels[7].label[171] 
	,\labels[7].label[170] ,\labels[7].label[169] ,\labels[7].label[168] 
	,\labels[7].label[167] ,\labels[7].label[166] ,\labels[7].label[165] 
	,\labels[7].label[164] ,\labels[7].label[163] ,\labels[7].label[162] 
	,\labels[7].label[161] ,\labels[7].label[160] ,\labels[7].label[159] 
	,\labels[7].label[158] ,\labels[7].label[157] ,\labels[7].label[156] 
	,\labels[7].label[155] ,\labels[7].label[154] ,\labels[7].label[153] 
	,\labels[7].label[152] ,\labels[7].label[151] ,\labels[7].label[150] 
	,\labels[7].label[149] ,\labels[7].label[148] ,\labels[7].label[147] 
	,\labels[7].label[146] ,\labels[7].label[145] ,\labels[7].label[144] 
	,\labels[7].label[143] ,\labels[7].label[142] ,\labels[7].label[141] 
	,\labels[7].label[140] ,\labels[7].label[139] ,\labels[7].label[138] 
	,\labels[7].label[137] ,\labels[7].label[136] ,\labels[7].label[135] 
	,\labels[7].label[134] ,\labels[7].label[133] ,\labels[7].label[132] 
	,\labels[7].label[131] ,\labels[7].label[130] ,\labels[7].label[129] 
	,\labels[7].label[128] ,\labels[7].label[127] ,\labels[7].label[126] 
	,\labels[7].label[125] ,\labels[7].label[124] ,\labels[7].label[123] 
	,\labels[7].label[122] ,\labels[7].label[121] ,\labels[7].label[120] 
	,\labels[7].label[119] ,\labels[7].label[118] ,\labels[7].label[117] 
	,\labels[7].label[116] ,\labels[7].label[115] ,\labels[7].label[114] 
	,\labels[7].label[113] ,\labels[7].label[112] ,\labels[7].label[111] 
	,\labels[7].label[110] ,\labels[7].label[109] ,\labels[7].label[108] 
	,\labels[7].label[107] ,\labels[7].label[106] ,\labels[7].label[105] 
	,\labels[7].label[104] ,\labels[7].label[103] ,\labels[7].label[102] 
	,\labels[7].label[101] ,\labels[7].label[100] ,\labels[7].label[99] 
	,\labels[7].label[98] ,\labels[7].label[97] ,\labels[7].label[96] 
	,\labels[7].label[95] ,\labels[7].label[94] ,\labels[7].label[93] 
	,\labels[7].label[92] ,\labels[7].label[91] ,\labels[7].label[90] 
	,\labels[7].label[89] ,\labels[7].label[88] ,\labels[7].label[87] 
	,\labels[7].label[86] ,\labels[7].label[85] ,\labels[7].label[84] 
	,\labels[7].label[83] ,\labels[7].label[82] ,\labels[7].label[81] 
	,\labels[7].label[80] ,\labels[7].label[79] ,\labels[7].label[78] 
	,\labels[7].label[77] ,\labels[7].label[76] ,\labels[7].label[75] 
	,\labels[7].label[74] ,\labels[7].label[73] ,\labels[7].label[72] 
	,\labels[7].label[71] ,\labels[7].label[70] ,\labels[7].label[69] 
	,\labels[7].label[68] ,\labels[7].label[67] ,\labels[7].label[66] 
	,\labels[7].label[65] ,\labels[7].label[64] ,\labels[7].label[63] 
	,\labels[7].label[62] ,\labels[7].label[61] ,\labels[7].label[60] 
	,\labels[7].label[59] ,\labels[7].label[58] ,\labels[7].label[57] 
	,\labels[7].label[56] ,\labels[7].label[55] ,\labels[7].label[54] 
	,\labels[7].label[53] ,\labels[7].label[52] ,\labels[7].label[51] 
	,\labels[7].label[50] ,\labels[7].label[49] ,\labels[7].label[48] 
	,\labels[7].label[47] ,\labels[7].label[46] ,\labels[7].label[45] 
	,\labels[7].label[44] ,\labels[7].label[43] ,\labels[7].label[42] 
	,\labels[7].label[41] ,\labels[7].label[40] ,\labels[7].label[39] 
	,\labels[7].label[38] ,\labels[7].label[37] ,\labels[7].label[36] 
	,\labels[7].label[35] ,\labels[7].label[34] ,\labels[7].label[33] 
	,\labels[7].label[32] ,\labels[7].label[31] ,\labels[7].label[30] 
	,\labels[7].label[29] ,\labels[7].label[28] ,\labels[7].label[27] 
	,\labels[7].label[26] ,\labels[7].label[25] ,\labels[7].label[24] 
	,\labels[7].label[23] ,\labels[7].label[22] ,\labels[7].label[21] 
	,\labels[7].label[20] ,\labels[7].label[19] ,\labels[7].label[18] 
	,\labels[7].label[17] ,\labels[7].label[16] ,\labels[7].label[15] 
	,\labels[7].label[14] ,\labels[7].label[13] ,\labels[7].label[12] 
	,\labels[7].label[11] ,\labels[7].label[10] ,\labels[7].label[9] 
	,\labels[7].label[8] ,\labels[7].label[7] ,\labels[7].label[6] 
	,\labels[7].label[5] ,\labels[7].label[4] ,\labels[7].label[3] 
	,\labels[7].label[2] ,\labels[7].label[1] ,\labels[7].label[0] 
	,\labels[7].delimiter_valid[0] ,\labels[7].delimiter[7] 
	,\labels[7].delimiter[6] ,\labels[7].delimiter[5] 
	,\labels[7].delimiter[4] ,\labels[7].delimiter[3] 
	,\labels[7].delimiter[2] ,\labels[7].delimiter[1] 
	,\labels[7].delimiter[0] ,\labels[6].guid_size[0] 
	,\labels[6].label_size[5] ,\labels[6].label_size[4] 
	,\labels[6].label_size[3] ,\labels[6].label_size[2] 
	,\labels[6].label_size[1] ,\labels[6].label_size[0] 
	,\labels[6].label[255] ,\labels[6].label[254] ,\labels[6].label[253] 
	,\labels[6].label[252] ,\labels[6].label[251] ,\labels[6].label[250] 
	,\labels[6].label[249] ,\labels[6].label[248] ,\labels[6].label[247] 
	,\labels[6].label[246] ,\labels[6].label[245] ,\labels[6].label[244] 
	,\labels[6].label[243] ,\labels[6].label[242] ,\labels[6].label[241] 
	,\labels[6].label[240] ,\labels[6].label[239] ,\labels[6].label[238] 
	,\labels[6].label[237] ,\labels[6].label[236] ,\labels[6].label[235] 
	,\labels[6].label[234] ,\labels[6].label[233] ,\labels[6].label[232] 
	,\labels[6].label[231] ,\labels[6].label[230] ,\labels[6].label[229] 
	,\labels[6].label[228] ,\labels[6].label[227] ,\labels[6].label[226] 
	,\labels[6].label[225] ,\labels[6].label[224] ,\labels[6].label[223] 
	,\labels[6].label[222] ,\labels[6].label[221] ,\labels[6].label[220] 
	,\labels[6].label[219] ,\labels[6].label[218] ,\labels[6].label[217] 
	,\labels[6].label[216] ,\labels[6].label[215] ,\labels[6].label[214] 
	,\labels[6].label[213] ,\labels[6].label[212] ,\labels[6].label[211] 
	,\labels[6].label[210] ,\labels[6].label[209] ,\labels[6].label[208] 
	,\labels[6].label[207] ,\labels[6].label[206] ,\labels[6].label[205] 
	,\labels[6].label[204] ,\labels[6].label[203] ,\labels[6].label[202] 
	,\labels[6].label[201] ,\labels[6].label[200] ,\labels[6].label[199] 
	,\labels[6].label[198] ,\labels[6].label[197] ,\labels[6].label[196] 
	,\labels[6].label[195] ,\labels[6].label[194] ,\labels[6].label[193] 
	,\labels[6].label[192] ,\labels[6].label[191] ,\labels[6].label[190] 
	,\labels[6].label[189] ,\labels[6].label[188] ,\labels[6].label[187] 
	,\labels[6].label[186] ,\labels[6].label[185] ,\labels[6].label[184] 
	,\labels[6].label[183] ,\labels[6].label[182] ,\labels[6].label[181] 
	,\labels[6].label[180] ,\labels[6].label[179] ,\labels[6].label[178] 
	,\labels[6].label[177] ,\labels[6].label[176] ,\labels[6].label[175] 
	,\labels[6].label[174] ,\labels[6].label[173] ,\labels[6].label[172] 
	,\labels[6].label[171] ,\labels[6].label[170] ,\labels[6].label[169] 
	,\labels[6].label[168] ,\labels[6].label[167] ,\labels[6].label[166] 
	,\labels[6].label[165] ,\labels[6].label[164] ,\labels[6].label[163] 
	,\labels[6].label[162] ,\labels[6].label[161] ,\labels[6].label[160] 
	,\labels[6].label[159] ,\labels[6].label[158] ,\labels[6].label[157] 
	,\labels[6].label[156] ,\labels[6].label[155] ,\labels[6].label[154] 
	,\labels[6].label[153] ,\labels[6].label[152] ,\labels[6].label[151] 
	,\labels[6].label[150] ,\labels[6].label[149] ,\labels[6].label[148] 
	,\labels[6].label[147] ,\labels[6].label[146] ,\labels[6].label[145] 
	,\labels[6].label[144] ,\labels[6].label[143] ,\labels[6].label[142] 
	,\labels[6].label[141] ,\labels[6].label[140] ,\labels[6].label[139] 
	,\labels[6].label[138] ,\labels[6].label[137] ,\labels[6].label[136] 
	,\labels[6].label[135] ,\labels[6].label[134] ,\labels[6].label[133] 
	,\labels[6].label[132] ,\labels[6].label[131] ,\labels[6].label[130] 
	,\labels[6].label[129] ,\labels[6].label[128] ,\labels[6].label[127] 
	,\labels[6].label[126] ,\labels[6].label[125] ,\labels[6].label[124] 
	,\labels[6].label[123] ,\labels[6].label[122] ,\labels[6].label[121] 
	,\labels[6].label[120] ,\labels[6].label[119] ,\labels[6].label[118] 
	,\labels[6].label[117] ,\labels[6].label[116] ,\labels[6].label[115] 
	,\labels[6].label[114] ,\labels[6].label[113] ,\labels[6].label[112] 
	,\labels[6].label[111] ,\labels[6].label[110] ,\labels[6].label[109] 
	,\labels[6].label[108] ,\labels[6].label[107] ,\labels[6].label[106] 
	,\labels[6].label[105] ,\labels[6].label[104] ,\labels[6].label[103] 
	,\labels[6].label[102] ,\labels[6].label[101] ,\labels[6].label[100] 
	,\labels[6].label[99] ,\labels[6].label[98] ,\labels[6].label[97] 
	,\labels[6].label[96] ,\labels[6].label[95] ,\labels[6].label[94] 
	,\labels[6].label[93] ,\labels[6].label[92] ,\labels[6].label[91] 
	,\labels[6].label[90] ,\labels[6].label[89] ,\labels[6].label[88] 
	,\labels[6].label[87] ,\labels[6].label[86] ,\labels[6].label[85] 
	,\labels[6].label[84] ,\labels[6].label[83] ,\labels[6].label[82] 
	,\labels[6].label[81] ,\labels[6].label[80] ,\labels[6].label[79] 
	,\labels[6].label[78] ,\labels[6].label[77] ,\labels[6].label[76] 
	,\labels[6].label[75] ,\labels[6].label[74] ,\labels[6].label[73] 
	,\labels[6].label[72] ,\labels[6].label[71] ,\labels[6].label[70] 
	,\labels[6].label[69] ,\labels[6].label[68] ,\labels[6].label[67] 
	,\labels[6].label[66] ,\labels[6].label[65] ,\labels[6].label[64] 
	,\labels[6].label[63] ,\labels[6].label[62] ,\labels[6].label[61] 
	,\labels[6].label[60] ,\labels[6].label[59] ,\labels[6].label[58] 
	,\labels[6].label[57] ,\labels[6].label[56] ,\labels[6].label[55] 
	,\labels[6].label[54] ,\labels[6].label[53] ,\labels[6].label[52] 
	,\labels[6].label[51] ,\labels[6].label[50] ,\labels[6].label[49] 
	,\labels[6].label[48] ,\labels[6].label[47] ,\labels[6].label[46] 
	,\labels[6].label[45] ,\labels[6].label[44] ,\labels[6].label[43] 
	,\labels[6].label[42] ,\labels[6].label[41] ,\labels[6].label[40] 
	,\labels[6].label[39] ,\labels[6].label[38] ,\labels[6].label[37] 
	,\labels[6].label[36] ,\labels[6].label[35] ,\labels[6].label[34] 
	,\labels[6].label[33] ,\labels[6].label[32] ,\labels[6].label[31] 
	,\labels[6].label[30] ,\labels[6].label[29] ,\labels[6].label[28] 
	,\labels[6].label[27] ,\labels[6].label[26] ,\labels[6].label[25] 
	,\labels[6].label[24] ,\labels[6].label[23] ,\labels[6].label[22] 
	,\labels[6].label[21] ,\labels[6].label[20] ,\labels[6].label[19] 
	,\labels[6].label[18] ,\labels[6].label[17] ,\labels[6].label[16] 
	,\labels[6].label[15] ,\labels[6].label[14] ,\labels[6].label[13] 
	,\labels[6].label[12] ,\labels[6].label[11] ,\labels[6].label[10] 
	,\labels[6].label[9] ,\labels[6].label[8] ,\labels[6].label[7] 
	,\labels[6].label[6] ,\labels[6].label[5] ,\labels[6].label[4] 
	,\labels[6].label[3] ,\labels[6].label[2] ,\labels[6].label[1] 
	,\labels[6].label[0] ,\labels[6].delimiter_valid[0] 
	,\labels[6].delimiter[7] ,\labels[6].delimiter[6] 
	,\labels[6].delimiter[5] ,\labels[6].delimiter[4] 
	,\labels[6].delimiter[3] ,\labels[6].delimiter[2] 
	,\labels[6].delimiter[1] ,\labels[6].delimiter[0] 
	,\labels[5].guid_size[0] ,\labels[5].label_size[5] 
	,\labels[5].label_size[4] ,\labels[5].label_size[3] 
	,\labels[5].label_size[2] ,\labels[5].label_size[1] 
	,\labels[5].label_size[0] ,\labels[5].label[255] 
	,\labels[5].label[254] ,\labels[5].label[253] ,\labels[5].label[252] 
	,\labels[5].label[251] ,\labels[5].label[250] ,\labels[5].label[249] 
	,\labels[5].label[248] ,\labels[5].label[247] ,\labels[5].label[246] 
	,\labels[5].label[245] ,\labels[5].label[244] ,\labels[5].label[243] 
	,\labels[5].label[242] ,\labels[5].label[241] ,\labels[5].label[240] 
	,\labels[5].label[239] ,\labels[5].label[238] ,\labels[5].label[237] 
	,\labels[5].label[236] ,\labels[5].label[235] ,\labels[5].label[234] 
	,\labels[5].label[233] ,\labels[5].label[232] ,\labels[5].label[231] 
	,\labels[5].label[230] ,\labels[5].label[229] ,\labels[5].label[228] 
	,\labels[5].label[227] ,\labels[5].label[226] ,\labels[5].label[225] 
	,\labels[5].label[224] ,\labels[5].label[223] ,\labels[5].label[222] 
	,\labels[5].label[221] ,\labels[5].label[220] ,\labels[5].label[219] 
	,\labels[5].label[218] ,\labels[5].label[217] ,\labels[5].label[216] 
	,\labels[5].label[215] ,\labels[5].label[214] ,\labels[5].label[213] 
	,\labels[5].label[212] ,\labels[5].label[211] ,\labels[5].label[210] 
	,\labels[5].label[209] ,\labels[5].label[208] ,\labels[5].label[207] 
	,\labels[5].label[206] ,\labels[5].label[205] ,\labels[5].label[204] 
	,\labels[5].label[203] ,\labels[5].label[202] ,\labels[5].label[201] 
	,\labels[5].label[200] ,\labels[5].label[199] ,\labels[5].label[198] 
	,\labels[5].label[197] ,\labels[5].label[196] ,\labels[5].label[195] 
	,\labels[5].label[194] ,\labels[5].label[193] ,\labels[5].label[192] 
	,\labels[5].label[191] ,\labels[5].label[190] ,\labels[5].label[189] 
	,\labels[5].label[188] ,\labels[5].label[187] ,\labels[5].label[186] 
	,\labels[5].label[185] ,\labels[5].label[184] ,\labels[5].label[183] 
	,\labels[5].label[182] ,\labels[5].label[181] ,\labels[5].label[180] 
	,\labels[5].label[179] ,\labels[5].label[178] ,\labels[5].label[177] 
	,\labels[5].label[176] ,\labels[5].label[175] ,\labels[5].label[174] 
	,\labels[5].label[173] ,\labels[5].label[172] ,\labels[5].label[171] 
	,\labels[5].label[170] ,\labels[5].label[169] ,\labels[5].label[168] 
	,\labels[5].label[167] ,\labels[5].label[166] ,\labels[5].label[165] 
	,\labels[5].label[164] ,\labels[5].label[163] ,\labels[5].label[162] 
	,\labels[5].label[161] ,\labels[5].label[160] ,\labels[5].label[159] 
	,\labels[5].label[158] ,\labels[5].label[157] ,\labels[5].label[156] 
	,\labels[5].label[155] ,\labels[5].label[154] ,\labels[5].label[153] 
	,\labels[5].label[152] ,\labels[5].label[151] ,\labels[5].label[150] 
	,\labels[5].label[149] ,\labels[5].label[148] ,\labels[5].label[147] 
	,\labels[5].label[146] ,\labels[5].label[145] ,\labels[5].label[144] 
	,\labels[5].label[143] ,\labels[5].label[142] ,\labels[5].label[141] 
	,\labels[5].label[140] ,\labels[5].label[139] ,\labels[5].label[138] 
	,\labels[5].label[137] ,\labels[5].label[136] ,\labels[5].label[135] 
	,\labels[5].label[134] ,\labels[5].label[133] ,\labels[5].label[132] 
	,\labels[5].label[131] ,\labels[5].label[130] ,\labels[5].label[129] 
	,\labels[5].label[128] ,\labels[5].label[127] ,\labels[5].label[126] 
	,\labels[5].label[125] ,\labels[5].label[124] ,\labels[5].label[123] 
	,\labels[5].label[122] ,\labels[5].label[121] ,\labels[5].label[120] 
	,\labels[5].label[119] ,\labels[5].label[118] ,\labels[5].label[117] 
	,\labels[5].label[116] ,\labels[5].label[115] ,\labels[5].label[114] 
	,\labels[5].label[113] ,\labels[5].label[112] ,\labels[5].label[111] 
	,\labels[5].label[110] ,\labels[5].label[109] ,\labels[5].label[108] 
	,\labels[5].label[107] ,\labels[5].label[106] ,\labels[5].label[105] 
	,\labels[5].label[104] ,\labels[5].label[103] ,\labels[5].label[102] 
	,\labels[5].label[101] ,\labels[5].label[100] ,\labels[5].label[99] 
	,\labels[5].label[98] ,\labels[5].label[97] ,\labels[5].label[96] 
	,\labels[5].label[95] ,\labels[5].label[94] ,\labels[5].label[93] 
	,\labels[5].label[92] ,\labels[5].label[91] ,\labels[5].label[90] 
	,\labels[5].label[89] ,\labels[5].label[88] ,\labels[5].label[87] 
	,\labels[5].label[86] ,\labels[5].label[85] ,\labels[5].label[84] 
	,\labels[5].label[83] ,\labels[5].label[82] ,\labels[5].label[81] 
	,\labels[5].label[80] ,\labels[5].label[79] ,\labels[5].label[78] 
	,\labels[5].label[77] ,\labels[5].label[76] ,\labels[5].label[75] 
	,\labels[5].label[74] ,\labels[5].label[73] ,\labels[5].label[72] 
	,\labels[5].label[71] ,\labels[5].label[70] ,\labels[5].label[69] 
	,\labels[5].label[68] ,\labels[5].label[67] ,\labels[5].label[66] 
	,\labels[5].label[65] ,\labels[5].label[64] ,\labels[5].label[63] 
	,\labels[5].label[62] ,\labels[5].label[61] ,\labels[5].label[60] 
	,\labels[5].label[59] ,\labels[5].label[58] ,\labels[5].label[57] 
	,\labels[5].label[56] ,\labels[5].label[55] ,\labels[5].label[54] 
	,\labels[5].label[53] ,\labels[5].label[52] ,\labels[5].label[51] 
	,\labels[5].label[50] ,\labels[5].label[49] ,\labels[5].label[48] 
	,\labels[5].label[47] ,\labels[5].label[46] ,\labels[5].label[45] 
	,\labels[5].label[44] ,\labels[5].label[43] ,\labels[5].label[42] 
	,\labels[5].label[41] ,\labels[5].label[40] ,\labels[5].label[39] 
	,\labels[5].label[38] ,\labels[5].label[37] ,\labels[5].label[36] 
	,\labels[5].label[35] ,\labels[5].label[34] ,\labels[5].label[33] 
	,\labels[5].label[32] ,\labels[5].label[31] ,\labels[5].label[30] 
	,\labels[5].label[29] ,\labels[5].label[28] ,\labels[5].label[27] 
	,\labels[5].label[26] ,\labels[5].label[25] ,\labels[5].label[24] 
	,\labels[5].label[23] ,\labels[5].label[22] ,\labels[5].label[21] 
	,\labels[5].label[20] ,\labels[5].label[19] ,\labels[5].label[18] 
	,\labels[5].label[17] ,\labels[5].label[16] ,\labels[5].label[15] 
	,\labels[5].label[14] ,\labels[5].label[13] ,\labels[5].label[12] 
	,\labels[5].label[11] ,\labels[5].label[10] ,\labels[5].label[9] 
	,\labels[5].label[8] ,\labels[5].label[7] ,\labels[5].label[6] 
	,\labels[5].label[5] ,\labels[5].label[4] ,\labels[5].label[3] 
	,\labels[5].label[2] ,\labels[5].label[1] ,\labels[5].label[0] 
	,\labels[5].delimiter_valid[0] ,\labels[5].delimiter[7] 
	,\labels[5].delimiter[6] ,\labels[5].delimiter[5] 
	,\labels[5].delimiter[4] ,\labels[5].delimiter[3] 
	,\labels[5].delimiter[2] ,\labels[5].delimiter[1] 
	,\labels[5].delimiter[0] ,\labels[4].guid_size[0] 
	,\labels[4].label_size[5] ,\labels[4].label_size[4] 
	,\labels[4].label_size[3] ,\labels[4].label_size[2] 
	,\labels[4].label_size[1] ,\labels[4].label_size[0] 
	,\labels[4].label[255] ,\labels[4].label[254] ,\labels[4].label[253] 
	,\labels[4].label[252] ,\labels[4].label[251] ,\labels[4].label[250] 
	,\labels[4].label[249] ,\labels[4].label[248] ,\labels[4].label[247] 
	,\labels[4].label[246] ,\labels[4].label[245] ,\labels[4].label[244] 
	,\labels[4].label[243] ,\labels[4].label[242] ,\labels[4].label[241] 
	,\labels[4].label[240] ,\labels[4].label[239] ,\labels[4].label[238] 
	,\labels[4].label[237] ,\labels[4].label[236] ,\labels[4].label[235] 
	,\labels[4].label[234] ,\labels[4].label[233] ,\labels[4].label[232] 
	,\labels[4].label[231] ,\labels[4].label[230] ,\labels[4].label[229] 
	,\labels[4].label[228] ,\labels[4].label[227] ,\labels[4].label[226] 
	,\labels[4].label[225] ,\labels[4].label[224] ,\labels[4].label[223] 
	,\labels[4].label[222] ,\labels[4].label[221] ,\labels[4].label[220] 
	,\labels[4].label[219] ,\labels[4].label[218] ,\labels[4].label[217] 
	,\labels[4].label[216] ,\labels[4].label[215] ,\labels[4].label[214] 
	,\labels[4].label[213] ,\labels[4].label[212] ,\labels[4].label[211] 
	,\labels[4].label[210] ,\labels[4].label[209] ,\labels[4].label[208] 
	,\labels[4].label[207] ,\labels[4].label[206] ,\labels[4].label[205] 
	,\labels[4].label[204] ,\labels[4].label[203] ,\labels[4].label[202] 
	,\labels[4].label[201] ,\labels[4].label[200] ,\labels[4].label[199] 
	,\labels[4].label[198] ,\labels[4].label[197] ,\labels[4].label[196] 
	,\labels[4].label[195] ,\labels[4].label[194] ,\labels[4].label[193] 
	,\labels[4].label[192] ,\labels[4].label[191] ,\labels[4].label[190] 
	,\labels[4].label[189] ,\labels[4].label[188] ,\labels[4].label[187] 
	,\labels[4].label[186] ,\labels[4].label[185] ,\labels[4].label[184] 
	,\labels[4].label[183] ,\labels[4].label[182] ,\labels[4].label[181] 
	,\labels[4].label[180] ,\labels[4].label[179] ,\labels[4].label[178] 
	,\labels[4].label[177] ,\labels[4].label[176] ,\labels[4].label[175] 
	,\labels[4].label[174] ,\labels[4].label[173] ,\labels[4].label[172] 
	,\labels[4].label[171] ,\labels[4].label[170] ,\labels[4].label[169] 
	,\labels[4].label[168] ,\labels[4].label[167] ,\labels[4].label[166] 
	,\labels[4].label[165] ,\labels[4].label[164] ,\labels[4].label[163] 
	,\labels[4].label[162] ,\labels[4].label[161] ,\labels[4].label[160] 
	,\labels[4].label[159] ,\labels[4].label[158] ,\labels[4].label[157] 
	,\labels[4].label[156] ,\labels[4].label[155] ,\labels[4].label[154] 
	,\labels[4].label[153] ,\labels[4].label[152] ,\labels[4].label[151] 
	,\labels[4].label[150] ,\labels[4].label[149] ,\labels[4].label[148] 
	,\labels[4].label[147] ,\labels[4].label[146] ,\labels[4].label[145] 
	,\labels[4].label[144] ,\labels[4].label[143] ,\labels[4].label[142] 
	,\labels[4].label[141] ,\labels[4].label[140] ,\labels[4].label[139] 
	,\labels[4].label[138] ,\labels[4].label[137] ,\labels[4].label[136] 
	,\labels[4].label[135] ,\labels[4].label[134] ,\labels[4].label[133] 
	,\labels[4].label[132] ,\labels[4].label[131] ,\labels[4].label[130] 
	,\labels[4].label[129] ,\labels[4].label[128] ,\labels[4].label[127] 
	,\labels[4].label[126] ,\labels[4].label[125] ,\labels[4].label[124] 
	,\labels[4].label[123] ,\labels[4].label[122] ,\labels[4].label[121] 
	,\labels[4].label[120] ,\labels[4].label[119] ,\labels[4].label[118] 
	,\labels[4].label[117] ,\labels[4].label[116] ,\labels[4].label[115] 
	,\labels[4].label[114] ,\labels[4].label[113] ,\labels[4].label[112] 
	,\labels[4].label[111] ,\labels[4].label[110] ,\labels[4].label[109] 
	,\labels[4].label[108] ,\labels[4].label[107] ,\labels[4].label[106] 
	,\labels[4].label[105] ,\labels[4].label[104] ,\labels[4].label[103] 
	,\labels[4].label[102] ,\labels[4].label[101] ,\labels[4].label[100] 
	,\labels[4].label[99] ,\labels[4].label[98] ,\labels[4].label[97] 
	,\labels[4].label[96] ,\labels[4].label[95] ,\labels[4].label[94] 
	,\labels[4].label[93] ,\labels[4].label[92] ,\labels[4].label[91] 
	,\labels[4].label[90] ,\labels[4].label[89] ,\labels[4].label[88] 
	,\labels[4].label[87] ,\labels[4].label[86] ,\labels[4].label[85] 
	,\labels[4].label[84] ,\labels[4].label[83] ,\labels[4].label[82] 
	,\labels[4].label[81] ,\labels[4].label[80] ,\labels[4].label[79] 
	,\labels[4].label[78] ,\labels[4].label[77] ,\labels[4].label[76] 
	,\labels[4].label[75] ,\labels[4].label[74] ,\labels[4].label[73] 
	,\labels[4].label[72] ,\labels[4].label[71] ,\labels[4].label[70] 
	,\labels[4].label[69] ,\labels[4].label[68] ,\labels[4].label[67] 
	,\labels[4].label[66] ,\labels[4].label[65] ,\labels[4].label[64] 
	,\labels[4].label[63] ,\labels[4].label[62] ,\labels[4].label[61] 
	,\labels[4].label[60] ,\labels[4].label[59] ,\labels[4].label[58] 
	,\labels[4].label[57] ,\labels[4].label[56] ,\labels[4].label[55] 
	,\labels[4].label[54] ,\labels[4].label[53] ,\labels[4].label[52] 
	,\labels[4].label[51] ,\labels[4].label[50] ,\labels[4].label[49] 
	,\labels[4].label[48] ,\labels[4].label[47] ,\labels[4].label[46] 
	,\labels[4].label[45] ,\labels[4].label[44] ,\labels[4].label[43] 
	,\labels[4].label[42] ,\labels[4].label[41] ,\labels[4].label[40] 
	,\labels[4].label[39] ,\labels[4].label[38] ,\labels[4].label[37] 
	,\labels[4].label[36] ,\labels[4].label[35] ,\labels[4].label[34] 
	,\labels[4].label[33] ,\labels[4].label[32] ,\labels[4].label[31] 
	,\labels[4].label[30] ,\labels[4].label[29] ,\labels[4].label[28] 
	,\labels[4].label[27] ,\labels[4].label[26] ,\labels[4].label[25] 
	,\labels[4].label[24] ,\labels[4].label[23] ,\labels[4].label[22] 
	,\labels[4].label[21] ,\labels[4].label[20] ,\labels[4].label[19] 
	,\labels[4].label[18] ,\labels[4].label[17] ,\labels[4].label[16] 
	,\labels[4].label[15] ,\labels[4].label[14] ,\labels[4].label[13] 
	,\labels[4].label[12] ,\labels[4].label[11] ,\labels[4].label[10] 
	,\labels[4].label[9] ,\labels[4].label[8] ,\labels[4].label[7] 
	,\labels[4].label[6] ,\labels[4].label[5] ,\labels[4].label[4] 
	,\labels[4].label[3] ,\labels[4].label[2] ,\labels[4].label[1] 
	,\labels[4].label[0] ,\labels[4].delimiter_valid[0] 
	,\labels[4].delimiter[7] ,\labels[4].delimiter[6] 
	,\labels[4].delimiter[5] ,\labels[4].delimiter[4] 
	,\labels[4].delimiter[3] ,\labels[4].delimiter[2] 
	,\labels[4].delimiter[1] ,\labels[4].delimiter[0] 
	,\labels[3].guid_size[0] ,\labels[3].label_size[5] 
	,\labels[3].label_size[4] ,\labels[3].label_size[3] 
	,\labels[3].label_size[2] ,\labels[3].label_size[1] 
	,\labels[3].label_size[0] ,\labels[3].label[255] 
	,\labels[3].label[254] ,\labels[3].label[253] ,\labels[3].label[252] 
	,\labels[3].label[251] ,\labels[3].label[250] ,\labels[3].label[249] 
	,\labels[3].label[248] ,\labels[3].label[247] ,\labels[3].label[246] 
	,\labels[3].label[245] ,\labels[3].label[244] ,\labels[3].label[243] 
	,\labels[3].label[242] ,\labels[3].label[241] ,\labels[3].label[240] 
	,\labels[3].label[239] ,\labels[3].label[238] ,\labels[3].label[237] 
	,\labels[3].label[236] ,\labels[3].label[235] ,\labels[3].label[234] 
	,\labels[3].label[233] ,\labels[3].label[232] ,\labels[3].label[231] 
	,\labels[3].label[230] ,\labels[3].label[229] ,\labels[3].label[228] 
	,\labels[3].label[227] ,\labels[3].label[226] ,\labels[3].label[225] 
	,\labels[3].label[224] ,\labels[3].label[223] ,\labels[3].label[222] 
	,\labels[3].label[221] ,\labels[3].label[220] ,\labels[3].label[219] 
	,\labels[3].label[218] ,\labels[3].label[217] ,\labels[3].label[216] 
	,\labels[3].label[215] ,\labels[3].label[214] ,\labels[3].label[213] 
	,\labels[3].label[212] ,\labels[3].label[211] ,\labels[3].label[210] 
	,\labels[3].label[209] ,\labels[3].label[208] ,\labels[3].label[207] 
	,\labels[3].label[206] ,\labels[3].label[205] ,\labels[3].label[204] 
	,\labels[3].label[203] ,\labels[3].label[202] ,\labels[3].label[201] 
	,\labels[3].label[200] ,\labels[3].label[199] ,\labels[3].label[198] 
	,\labels[3].label[197] ,\labels[3].label[196] ,\labels[3].label[195] 
	,\labels[3].label[194] ,\labels[3].label[193] ,\labels[3].label[192] 
	,\labels[3].label[191] ,\labels[3].label[190] ,\labels[3].label[189] 
	,\labels[3].label[188] ,\labels[3].label[187] ,\labels[3].label[186] 
	,\labels[3].label[185] ,\labels[3].label[184] ,\labels[3].label[183] 
	,\labels[3].label[182] ,\labels[3].label[181] ,\labels[3].label[180] 
	,\labels[3].label[179] ,\labels[3].label[178] ,\labels[3].label[177] 
	,\labels[3].label[176] ,\labels[3].label[175] ,\labels[3].label[174] 
	,\labels[3].label[173] ,\labels[3].label[172] ,\labels[3].label[171] 
	,\labels[3].label[170] ,\labels[3].label[169] ,\labels[3].label[168] 
	,\labels[3].label[167] ,\labels[3].label[166] ,\labels[3].label[165] 
	,\labels[3].label[164] ,\labels[3].label[163] ,\labels[3].label[162] 
	,\labels[3].label[161] ,\labels[3].label[160] ,\labels[3].label[159] 
	,\labels[3].label[158] ,\labels[3].label[157] ,\labels[3].label[156] 
	,\labels[3].label[155] ,\labels[3].label[154] ,\labels[3].label[153] 
	,\labels[3].label[152] ,\labels[3].label[151] ,\labels[3].label[150] 
	,\labels[3].label[149] ,\labels[3].label[148] ,\labels[3].label[147] 
	,\labels[3].label[146] ,\labels[3].label[145] ,\labels[3].label[144] 
	,\labels[3].label[143] ,\labels[3].label[142] ,\labels[3].label[141] 
	,\labels[3].label[140] ,\labels[3].label[139] ,\labels[3].label[138] 
	,\labels[3].label[137] ,\labels[3].label[136] ,\labels[3].label[135] 
	,\labels[3].label[134] ,\labels[3].label[133] ,\labels[3].label[132] 
	,\labels[3].label[131] ,\labels[3].label[130] ,\labels[3].label[129] 
	,\labels[3].label[128] ,\labels[3].label[127] ,\labels[3].label[126] 
	,\labels[3].label[125] ,\labels[3].label[124] ,\labels[3].label[123] 
	,\labels[3].label[122] ,\labels[3].label[121] ,\labels[3].label[120] 
	,\labels[3].label[119] ,\labels[3].label[118] ,\labels[3].label[117] 
	,\labels[3].label[116] ,\labels[3].label[115] ,\labels[3].label[114] 
	,\labels[3].label[113] ,\labels[3].label[112] ,\labels[3].label[111] 
	,\labels[3].label[110] ,\labels[3].label[109] ,\labels[3].label[108] 
	,\labels[3].label[107] ,\labels[3].label[106] ,\labels[3].label[105] 
	,\labels[3].label[104] ,\labels[3].label[103] ,\labels[3].label[102] 
	,\labels[3].label[101] ,\labels[3].label[100] ,\labels[3].label[99] 
	,\labels[3].label[98] ,\labels[3].label[97] ,\labels[3].label[96] 
	,\labels[3].label[95] ,\labels[3].label[94] ,\labels[3].label[93] 
	,\labels[3].label[92] ,\labels[3].label[91] ,\labels[3].label[90] 
	,\labels[3].label[89] ,\labels[3].label[88] ,\labels[3].label[87] 
	,\labels[3].label[86] ,\labels[3].label[85] ,\labels[3].label[84] 
	,\labels[3].label[83] ,\labels[3].label[82] ,\labels[3].label[81] 
	,\labels[3].label[80] ,\labels[3].label[79] ,\labels[3].label[78] 
	,\labels[3].label[77] ,\labels[3].label[76] ,\labels[3].label[75] 
	,\labels[3].label[74] ,\labels[3].label[73] ,\labels[3].label[72] 
	,\labels[3].label[71] ,\labels[3].label[70] ,\labels[3].label[69] 
	,\labels[3].label[68] ,\labels[3].label[67] ,\labels[3].label[66] 
	,\labels[3].label[65] ,\labels[3].label[64] ,\labels[3].label[63] 
	,\labels[3].label[62] ,\labels[3].label[61] ,\labels[3].label[60] 
	,\labels[3].label[59] ,\labels[3].label[58] ,\labels[3].label[57] 
	,\labels[3].label[56] ,\labels[3].label[55] ,\labels[3].label[54] 
	,\labels[3].label[53] ,\labels[3].label[52] ,\labels[3].label[51] 
	,\labels[3].label[50] ,\labels[3].label[49] ,\labels[3].label[48] 
	,\labels[3].label[47] ,\labels[3].label[46] ,\labels[3].label[45] 
	,\labels[3].label[44] ,\labels[3].label[43] ,\labels[3].label[42] 
	,\labels[3].label[41] ,\labels[3].label[40] ,\labels[3].label[39] 
	,\labels[3].label[38] ,\labels[3].label[37] ,\labels[3].label[36] 
	,\labels[3].label[35] ,\labels[3].label[34] ,\labels[3].label[33] 
	,\labels[3].label[32] ,\labels[3].label[31] ,\labels[3].label[30] 
	,\labels[3].label[29] ,\labels[3].label[28] ,\labels[3].label[27] 
	,\labels[3].label[26] ,\labels[3].label[25] ,\labels[3].label[24] 
	,\labels[3].label[23] ,\labels[3].label[22] ,\labels[3].label[21] 
	,\labels[3].label[20] ,\labels[3].label[19] ,\labels[3].label[18] 
	,\labels[3].label[17] ,\labels[3].label[16] ,\labels[3].label[15] 
	,\labels[3].label[14] ,\labels[3].label[13] ,\labels[3].label[12] 
	,\labels[3].label[11] ,\labels[3].label[10] ,\labels[3].label[9] 
	,\labels[3].label[8] ,\labels[3].label[7] ,\labels[3].label[6] 
	,\labels[3].label[5] ,\labels[3].label[4] ,\labels[3].label[3] 
	,\labels[3].label[2] ,\labels[3].label[1] ,\labels[3].label[0] 
	,\labels[3].delimiter_valid[0] ,\labels[3].delimiter[7] 
	,\labels[3].delimiter[6] ,\labels[3].delimiter[5] 
	,\labels[3].delimiter[4] ,\labels[3].delimiter[3] 
	,\labels[3].delimiter[2] ,\labels[3].delimiter[1] 
	,\labels[3].delimiter[0] ,\labels[2].guid_size[0] 
	,\labels[2].label_size[5] ,\labels[2].label_size[4] 
	,\labels[2].label_size[3] ,\labels[2].label_size[2] 
	,\labels[2].label_size[1] ,\labels[2].label_size[0] 
	,\labels[2].label[255] ,\labels[2].label[254] ,\labels[2].label[253] 
	,\labels[2].label[252] ,\labels[2].label[251] ,\labels[2].label[250] 
	,\labels[2].label[249] ,\labels[2].label[248] ,\labels[2].label[247] 
	,\labels[2].label[246] ,\labels[2].label[245] ,\labels[2].label[244] 
	,\labels[2].label[243] ,\labels[2].label[242] ,\labels[2].label[241] 
	,\labels[2].label[240] ,\labels[2].label[239] ,\labels[2].label[238] 
	,\labels[2].label[237] ,\labels[2].label[236] ,\labels[2].label[235] 
	,\labels[2].label[234] ,\labels[2].label[233] ,\labels[2].label[232] 
	,\labels[2].label[231] ,\labels[2].label[230] ,\labels[2].label[229] 
	,\labels[2].label[228] ,\labels[2].label[227] ,\labels[2].label[226] 
	,\labels[2].label[225] ,\labels[2].label[224] ,\labels[2].label[223] 
	,\labels[2].label[222] ,\labels[2].label[221] ,\labels[2].label[220] 
	,\labels[2].label[219] ,\labels[2].label[218] ,\labels[2].label[217] 
	,\labels[2].label[216] ,\labels[2].label[215] ,\labels[2].label[214] 
	,\labels[2].label[213] ,\labels[2].label[212] ,\labels[2].label[211] 
	,\labels[2].label[210] ,\labels[2].label[209] ,\labels[2].label[208] 
	,\labels[2].label[207] ,\labels[2].label[206] ,\labels[2].label[205] 
	,\labels[2].label[204] ,\labels[2].label[203] ,\labels[2].label[202] 
	,\labels[2].label[201] ,\labels[2].label[200] ,\labels[2].label[199] 
	,\labels[2].label[198] ,\labels[2].label[197] ,\labels[2].label[196] 
	,\labels[2].label[195] ,\labels[2].label[194] ,\labels[2].label[193] 
	,\labels[2].label[192] ,\labels[2].label[191] ,\labels[2].label[190] 
	,\labels[2].label[189] ,\labels[2].label[188] ,\labels[2].label[187] 
	,\labels[2].label[186] ,\labels[2].label[185] ,\labels[2].label[184] 
	,\labels[2].label[183] ,\labels[2].label[182] ,\labels[2].label[181] 
	,\labels[2].label[180] ,\labels[2].label[179] ,\labels[2].label[178] 
	,\labels[2].label[177] ,\labels[2].label[176] ,\labels[2].label[175] 
	,\labels[2].label[174] ,\labels[2].label[173] ,\labels[2].label[172] 
	,\labels[2].label[171] ,\labels[2].label[170] ,\labels[2].label[169] 
	,\labels[2].label[168] ,\labels[2].label[167] ,\labels[2].label[166] 
	,\labels[2].label[165] ,\labels[2].label[164] ,\labels[2].label[163] 
	,\labels[2].label[162] ,\labels[2].label[161] ,\labels[2].label[160] 
	,\labels[2].label[159] ,\labels[2].label[158] ,\labels[2].label[157] 
	,\labels[2].label[156] ,\labels[2].label[155] ,\labels[2].label[154] 
	,\labels[2].label[153] ,\labels[2].label[152] ,\labels[2].label[151] 
	,\labels[2].label[150] ,\labels[2].label[149] ,\labels[2].label[148] 
	,\labels[2].label[147] ,\labels[2].label[146] ,\labels[2].label[145] 
	,\labels[2].label[144] ,\labels[2].label[143] ,\labels[2].label[142] 
	,\labels[2].label[141] ,\labels[2].label[140] ,\labels[2].label[139] 
	,\labels[2].label[138] ,\labels[2].label[137] ,\labels[2].label[136] 
	,\labels[2].label[135] ,\labels[2].label[134] ,\labels[2].label[133] 
	,\labels[2].label[132] ,\labels[2].label[131] ,\labels[2].label[130] 
	,\labels[2].label[129] ,\labels[2].label[128] ,\labels[2].label[127] 
	,\labels[2].label[126] ,\labels[2].label[125] ,\labels[2].label[124] 
	,\labels[2].label[123] ,\labels[2].label[122] ,\labels[2].label[121] 
	,\labels[2].label[120] ,\labels[2].label[119] ,\labels[2].label[118] 
	,\labels[2].label[117] ,\labels[2].label[116] ,\labels[2].label[115] 
	,\labels[2].label[114] ,\labels[2].label[113] ,\labels[2].label[112] 
	,\labels[2].label[111] ,\labels[2].label[110] ,\labels[2].label[109] 
	,\labels[2].label[108] ,\labels[2].label[107] ,\labels[2].label[106] 
	,\labels[2].label[105] ,\labels[2].label[104] ,\labels[2].label[103] 
	,\labels[2].label[102] ,\labels[2].label[101] ,\labels[2].label[100] 
	,\labels[2].label[99] ,\labels[2].label[98] ,\labels[2].label[97] 
	,\labels[2].label[96] ,\labels[2].label[95] ,\labels[2].label[94] 
	,\labels[2].label[93] ,\labels[2].label[92] ,\labels[2].label[91] 
	,\labels[2].label[90] ,\labels[2].label[89] ,\labels[2].label[88] 
	,\labels[2].label[87] ,\labels[2].label[86] ,\labels[2].label[85] 
	,\labels[2].label[84] ,\labels[2].label[83] ,\labels[2].label[82] 
	,\labels[2].label[81] ,\labels[2].label[80] ,\labels[2].label[79] 
	,\labels[2].label[78] ,\labels[2].label[77] ,\labels[2].label[76] 
	,\labels[2].label[75] ,\labels[2].label[74] ,\labels[2].label[73] 
	,\labels[2].label[72] ,\labels[2].label[71] ,\labels[2].label[70] 
	,\labels[2].label[69] ,\labels[2].label[68] ,\labels[2].label[67] 
	,\labels[2].label[66] ,\labels[2].label[65] ,\labels[2].label[64] 
	,\labels[2].label[63] ,\labels[2].label[62] ,\labels[2].label[61] 
	,\labels[2].label[60] ,\labels[2].label[59] ,\labels[2].label[58] 
	,\labels[2].label[57] ,\labels[2].label[56] ,\labels[2].label[55] 
	,\labels[2].label[54] ,\labels[2].label[53] ,\labels[2].label[52] 
	,\labels[2].label[51] ,\labels[2].label[50] ,\labels[2].label[49] 
	,\labels[2].label[48] ,\labels[2].label[47] ,\labels[2].label[46] 
	,\labels[2].label[45] ,\labels[2].label[44] ,\labels[2].label[43] 
	,\labels[2].label[42] ,\labels[2].label[41] ,\labels[2].label[40] 
	,\labels[2].label[39] ,\labels[2].label[38] ,\labels[2].label[37] 
	,\labels[2].label[36] ,\labels[2].label[35] ,\labels[2].label[34] 
	,\labels[2].label[33] ,\labels[2].label[32] ,\labels[2].label[31] 
	,\labels[2].label[30] ,\labels[2].label[29] ,\labels[2].label[28] 
	,\labels[2].label[27] ,\labels[2].label[26] ,\labels[2].label[25] 
	,\labels[2].label[24] ,\labels[2].label[23] ,\labels[2].label[22] 
	,\labels[2].label[21] ,\labels[2].label[20] ,\labels[2].label[19] 
	,\labels[2].label[18] ,\labels[2].label[17] ,\labels[2].label[16] 
	,\labels[2].label[15] ,\labels[2].label[14] ,\labels[2].label[13] 
	,\labels[2].label[12] ,\labels[2].label[11] ,\labels[2].label[10] 
	,\labels[2].label[9] ,\labels[2].label[8] ,\labels[2].label[7] 
	,\labels[2].label[6] ,\labels[2].label[5] ,\labels[2].label[4] 
	,\labels[2].label[3] ,\labels[2].label[2] ,\labels[2].label[1] 
	,\labels[2].label[0] ,\labels[2].delimiter_valid[0] 
	,\labels[2].delimiter[7] ,\labels[2].delimiter[6] 
	,\labels[2].delimiter[5] ,\labels[2].delimiter[4] 
	,\labels[2].delimiter[3] ,\labels[2].delimiter[2] 
	,\labels[2].delimiter[1] ,\labels[2].delimiter[0] 
	,\labels[1].guid_size[0] ,\labels[1].label_size[5] 
	,\labels[1].label_size[4] ,\labels[1].label_size[3] 
	,\labels[1].label_size[2] ,\labels[1].label_size[1] 
	,\labels[1].label_size[0] ,\labels[1].label[255] 
	,\labels[1].label[254] ,\labels[1].label[253] ,\labels[1].label[252] 
	,\labels[1].label[251] ,\labels[1].label[250] ,\labels[1].label[249] 
	,\labels[1].label[248] ,\labels[1].label[247] ,\labels[1].label[246] 
	,\labels[1].label[245] ,\labels[1].label[244] ,\labels[1].label[243] 
	,\labels[1].label[242] ,\labels[1].label[241] ,\labels[1].label[240] 
	,\labels[1].label[239] ,\labels[1].label[238] ,\labels[1].label[237] 
	,\labels[1].label[236] ,\labels[1].label[235] ,\labels[1].label[234] 
	,\labels[1].label[233] ,\labels[1].label[232] ,\labels[1].label[231] 
	,\labels[1].label[230] ,\labels[1].label[229] ,\labels[1].label[228] 
	,\labels[1].label[227] ,\labels[1].label[226] ,\labels[1].label[225] 
	,\labels[1].label[224] ,\labels[1].label[223] ,\labels[1].label[222] 
	,\labels[1].label[221] ,\labels[1].label[220] ,\labels[1].label[219] 
	,\labels[1].label[218] ,\labels[1].label[217] ,\labels[1].label[216] 
	,\labels[1].label[215] ,\labels[1].label[214] ,\labels[1].label[213] 
	,\labels[1].label[212] ,\labels[1].label[211] ,\labels[1].label[210] 
	,\labels[1].label[209] ,\labels[1].label[208] ,\labels[1].label[207] 
	,\labels[1].label[206] ,\labels[1].label[205] ,\labels[1].label[204] 
	,\labels[1].label[203] ,\labels[1].label[202] ,\labels[1].label[201] 
	,\labels[1].label[200] ,\labels[1].label[199] ,\labels[1].label[198] 
	,\labels[1].label[197] ,\labels[1].label[196] ,\labels[1].label[195] 
	,\labels[1].label[194] ,\labels[1].label[193] ,\labels[1].label[192] 
	,\labels[1].label[191] ,\labels[1].label[190] ,\labels[1].label[189] 
	,\labels[1].label[188] ,\labels[1].label[187] ,\labels[1].label[186] 
	,\labels[1].label[185] ,\labels[1].label[184] ,\labels[1].label[183] 
	,\labels[1].label[182] ,\labels[1].label[181] ,\labels[1].label[180] 
	,\labels[1].label[179] ,\labels[1].label[178] ,\labels[1].label[177] 
	,\labels[1].label[176] ,\labels[1].label[175] ,\labels[1].label[174] 
	,\labels[1].label[173] ,\labels[1].label[172] ,\labels[1].label[171] 
	,\labels[1].label[170] ,\labels[1].label[169] ,\labels[1].label[168] 
	,\labels[1].label[167] ,\labels[1].label[166] ,\labels[1].label[165] 
	,\labels[1].label[164] ,\labels[1].label[163] ,\labels[1].label[162] 
	,\labels[1].label[161] ,\labels[1].label[160] ,\labels[1].label[159] 
	,\labels[1].label[158] ,\labels[1].label[157] ,\labels[1].label[156] 
	,\labels[1].label[155] ,\labels[1].label[154] ,\labels[1].label[153] 
	,\labels[1].label[152] ,\labels[1].label[151] ,\labels[1].label[150] 
	,\labels[1].label[149] ,\labels[1].label[148] ,\labels[1].label[147] 
	,\labels[1].label[146] ,\labels[1].label[145] ,\labels[1].label[144] 
	,\labels[1].label[143] ,\labels[1].label[142] ,\labels[1].label[141] 
	,\labels[1].label[140] ,\labels[1].label[139] ,\labels[1].label[138] 
	,\labels[1].label[137] ,\labels[1].label[136] ,\labels[1].label[135] 
	,\labels[1].label[134] ,\labels[1].label[133] ,\labels[1].label[132] 
	,\labels[1].label[131] ,\labels[1].label[130] ,\labels[1].label[129] 
	,\labels[1].label[128] ,\labels[1].label[127] ,\labels[1].label[126] 
	,\labels[1].label[125] ,\labels[1].label[124] ,\labels[1].label[123] 
	,\labels[1].label[122] ,\labels[1].label[121] ,\labels[1].label[120] 
	,\labels[1].label[119] ,\labels[1].label[118] ,\labels[1].label[117] 
	,\labels[1].label[116] ,\labels[1].label[115] ,\labels[1].label[114] 
	,\labels[1].label[113] ,\labels[1].label[112] ,\labels[1].label[111] 
	,\labels[1].label[110] ,\labels[1].label[109] ,\labels[1].label[108] 
	,\labels[1].label[107] ,\labels[1].label[106] ,\labels[1].label[105] 
	,\labels[1].label[104] ,\labels[1].label[103] ,\labels[1].label[102] 
	,\labels[1].label[101] ,\labels[1].label[100] ,\labels[1].label[99] 
	,\labels[1].label[98] ,\labels[1].label[97] ,\labels[1].label[96] 
	,\labels[1].label[95] ,\labels[1].label[94] ,\labels[1].label[93] 
	,\labels[1].label[92] ,\labels[1].label[91] ,\labels[1].label[90] 
	,\labels[1].label[89] ,\labels[1].label[88] ,\labels[1].label[87] 
	,\labels[1].label[86] ,\labels[1].label[85] ,\labels[1].label[84] 
	,\labels[1].label[83] ,\labels[1].label[82] ,\labels[1].label[81] 
	,\labels[1].label[80] ,\labels[1].label[79] ,\labels[1].label[78] 
	,\labels[1].label[77] ,\labels[1].label[76] ,\labels[1].label[75] 
	,\labels[1].label[74] ,\labels[1].label[73] ,\labels[1].label[72] 
	,\labels[1].label[71] ,\labels[1].label[70] ,\labels[1].label[69] 
	,\labels[1].label[68] ,\labels[1].label[67] ,\labels[1].label[66] 
	,\labels[1].label[65] ,\labels[1].label[64] ,\labels[1].label[63] 
	,\labels[1].label[62] ,\labels[1].label[61] ,\labels[1].label[60] 
	,\labels[1].label[59] ,\labels[1].label[58] ,\labels[1].label[57] 
	,\labels[1].label[56] ,\labels[1].label[55] ,\labels[1].label[54] 
	,\labels[1].label[53] ,\labels[1].label[52] ,\labels[1].label[51] 
	,\labels[1].label[50] ,\labels[1].label[49] ,\labels[1].label[48] 
	,\labels[1].label[47] ,\labels[1].label[46] ,\labels[1].label[45] 
	,\labels[1].label[44] ,\labels[1].label[43] ,\labels[1].label[42] 
	,\labels[1].label[41] ,\labels[1].label[40] ,\labels[1].label[39] 
	,\labels[1].label[38] ,\labels[1].label[37] ,\labels[1].label[36] 
	,\labels[1].label[35] ,\labels[1].label[34] ,\labels[1].label[33] 
	,\labels[1].label[32] ,\labels[1].label[31] ,\labels[1].label[30] 
	,\labels[1].label[29] ,\labels[1].label[28] ,\labels[1].label[27] 
	,\labels[1].label[26] ,\labels[1].label[25] ,\labels[1].label[24] 
	,\labels[1].label[23] ,\labels[1].label[22] ,\labels[1].label[21] 
	,\labels[1].label[20] ,\labels[1].label[19] ,\labels[1].label[18] 
	,\labels[1].label[17] ,\labels[1].label[16] ,\labels[1].label[15] 
	,\labels[1].label[14] ,\labels[1].label[13] ,\labels[1].label[12] 
	,\labels[1].label[11] ,\labels[1].label[10] ,\labels[1].label[9] 
	,\labels[1].label[8] ,\labels[1].label[7] ,\labels[1].label[6] 
	,\labels[1].label[5] ,\labels[1].label[4] ,\labels[1].label[3] 
	,\labels[1].label[2] ,\labels[1].label[1] ,\labels[1].label[0] 
	,\labels[1].delimiter_valid[0] ,\labels[1].delimiter[7] 
	,\labels[1].delimiter[6] ,\labels[1].delimiter[5] 
	,\labels[1].delimiter[4] ,\labels[1].delimiter[3] 
	,\labels[1].delimiter[2] ,\labels[1].delimiter[1] 
	,\labels[1].delimiter[0] ,\labels[0].guid_size[0] 
	,\labels[0].label_size[5] ,\labels[0].label_size[4] 
	,\labels[0].label_size[3] ,\labels[0].label_size[2] 
	,\labels[0].label_size[1] ,\labels[0].label_size[0] 
	,\labels[0].label[255] ,\labels[0].label[254] ,\labels[0].label[253] 
	,\labels[0].label[252] ,\labels[0].label[251] ,\labels[0].label[250] 
	,\labels[0].label[249] ,\labels[0].label[248] ,\labels[0].label[247] 
	,\labels[0].label[246] ,\labels[0].label[245] ,\labels[0].label[244] 
	,\labels[0].label[243] ,\labels[0].label[242] ,\labels[0].label[241] 
	,\labels[0].label[240] ,\labels[0].label[239] ,\labels[0].label[238] 
	,\labels[0].label[237] ,\labels[0].label[236] ,\labels[0].label[235] 
	,\labels[0].label[234] ,\labels[0].label[233] ,\labels[0].label[232] 
	,\labels[0].label[231] ,\labels[0].label[230] ,\labels[0].label[229] 
	,\labels[0].label[228] ,\labels[0].label[227] ,\labels[0].label[226] 
	,\labels[0].label[225] ,\labels[0].label[224] ,\labels[0].label[223] 
	,\labels[0].label[222] ,\labels[0].label[221] ,\labels[0].label[220] 
	,\labels[0].label[219] ,\labels[0].label[218] ,\labels[0].label[217] 
	,\labels[0].label[216] ,\labels[0].label[215] ,\labels[0].label[214] 
	,\labels[0].label[213] ,\labels[0].label[212] ,\labels[0].label[211] 
	,\labels[0].label[210] ,\labels[0].label[209] ,\labels[0].label[208] 
	,\labels[0].label[207] ,\labels[0].label[206] ,\labels[0].label[205] 
	,\labels[0].label[204] ,\labels[0].label[203] ,\labels[0].label[202] 
	,\labels[0].label[201] ,\labels[0].label[200] ,\labels[0].label[199] 
	,\labels[0].label[198] ,\labels[0].label[197] ,\labels[0].label[196] 
	,\labels[0].label[195] ,\labels[0].label[194] ,\labels[0].label[193] 
	,\labels[0].label[192] ,\labels[0].label[191] ,\labels[0].label[190] 
	,\labels[0].label[189] ,\labels[0].label[188] ,\labels[0].label[187] 
	,\labels[0].label[186] ,\labels[0].label[185] ,\labels[0].label[184] 
	,\labels[0].label[183] ,\labels[0].label[182] ,\labels[0].label[181] 
	,\labels[0].label[180] ,\labels[0].label[179] ,\labels[0].label[178] 
	,\labels[0].label[177] ,\labels[0].label[176] ,\labels[0].label[175] 
	,\labels[0].label[174] ,\labels[0].label[173] ,\labels[0].label[172] 
	,\labels[0].label[171] ,\labels[0].label[170] ,\labels[0].label[169] 
	,\labels[0].label[168] ,\labels[0].label[167] ,\labels[0].label[166] 
	,\labels[0].label[165] ,\labels[0].label[164] ,\labels[0].label[163] 
	,\labels[0].label[162] ,\labels[0].label[161] ,\labels[0].label[160] 
	,\labels[0].label[159] ,\labels[0].label[158] ,\labels[0].label[157] 
	,\labels[0].label[156] ,\labels[0].label[155] ,\labels[0].label[154] 
	,\labels[0].label[153] ,\labels[0].label[152] ,\labels[0].label[151] 
	,\labels[0].label[150] ,\labels[0].label[149] ,\labels[0].label[148] 
	,\labels[0].label[147] ,\labels[0].label[146] ,\labels[0].label[145] 
	,\labels[0].label[144] ,\labels[0].label[143] ,\labels[0].label[142] 
	,\labels[0].label[141] ,\labels[0].label[140] ,\labels[0].label[139] 
	,\labels[0].label[138] ,\labels[0].label[137] ,\labels[0].label[136] 
	,\labels[0].label[135] ,\labels[0].label[134] ,\labels[0].label[133] 
	,\labels[0].label[132] ,\labels[0].label[131] ,\labels[0].label[130] 
	,\labels[0].label[129] ,\labels[0].label[128] ,\labels[0].label[127] 
	,\labels[0].label[126] ,\labels[0].label[125] ,\labels[0].label[124] 
	,\labels[0].label[123] ,\labels[0].label[122] ,\labels[0].label[121] 
	,\labels[0].label[120] ,\labels[0].label[119] ,\labels[0].label[118] 
	,\labels[0].label[117] ,\labels[0].label[116] ,\labels[0].label[115] 
	,\labels[0].label[114] ,\labels[0].label[113] ,\labels[0].label[112] 
	,\labels[0].label[111] ,\labels[0].label[110] ,\labels[0].label[109] 
	,\labels[0].label[108] ,\labels[0].label[107] ,\labels[0].label[106] 
	,\labels[0].label[105] ,\labels[0].label[104] ,\labels[0].label[103] 
	,\labels[0].label[102] ,\labels[0].label[101] ,\labels[0].label[100] 
	,\labels[0].label[99] ,\labels[0].label[98] ,\labels[0].label[97] 
	,\labels[0].label[96] ,\labels[0].label[95] ,\labels[0].label[94] 
	,\labels[0].label[93] ,\labels[0].label[92] ,\labels[0].label[91] 
	,\labels[0].label[90] ,\labels[0].label[89] ,\labels[0].label[88] 
	,\labels[0].label[87] ,\labels[0].label[86] ,\labels[0].label[85] 
	,\labels[0].label[84] ,\labels[0].label[83] ,\labels[0].label[82] 
	,\labels[0].label[81] ,\labels[0].label[80] ,\labels[0].label[79] 
	,\labels[0].label[78] ,\labels[0].label[77] ,\labels[0].label[76] 
	,\labels[0].label[75] ,\labels[0].label[74] ,\labels[0].label[73] 
	,\labels[0].label[72] ,\labels[0].label[71] ,\labels[0].label[70] 
	,\labels[0].label[69] ,\labels[0].label[68] ,\labels[0].label[67] 
	,\labels[0].label[66] ,\labels[0].label[65] ,\labels[0].label[64] 
	,\labels[0].label[63] ,\labels[0].label[62] ,\labels[0].label[61] 
	,\labels[0].label[60] ,\labels[0].label[59] ,\labels[0].label[58] 
	,\labels[0].label[57] ,\labels[0].label[56] ,\labels[0].label[55] 
	,\labels[0].label[54] ,\labels[0].label[53] ,\labels[0].label[52] 
	,\labels[0].label[51] ,\labels[0].label[50] ,\labels[0].label[49] 
	,\labels[0].label[48] ,\labels[0].label[47] ,\labels[0].label[46] 
	,\labels[0].label[45] ,\labels[0].label[44] ,\labels[0].label[43] 
	,\labels[0].label[42] ,\labels[0].label[41] ,\labels[0].label[40] 
	,\labels[0].label[39] ,\labels[0].label[38] ,\labels[0].label[37] 
	,\labels[0].label[36] ,\labels[0].label[35] ,\labels[0].label[34] 
	,\labels[0].label[33] ,\labels[0].label[32] ,\labels[0].label[31] 
	,\labels[0].label[30] ,\labels[0].label[29] ,\labels[0].label[28] 
	,\labels[0].label[27] ,\labels[0].label[26] ,\labels[0].label[25] 
	,\labels[0].label[24] ,\labels[0].label[23] ,\labels[0].label[22] 
	,\labels[0].label[21] ,\labels[0].label[20] ,\labels[0].label[19] 
	,\labels[0].label[18] ,\labels[0].label[17] ,\labels[0].label[16] 
	,\labels[0].label[15] ,\labels[0].label[14] ,\labels[0].label[13] 
	,\labels[0].label[12] ,\labels[0].label[11] ,\labels[0].label[10] 
	,\labels[0].label[9] ,\labels[0].label[8] ,\labels[0].label[7] 
	,\labels[0].label[6] ,\labels[0].label[5] ,\labels[0].label[4] 
	,\labels[0].label[3] ,\labels[0].label[2] ,\labels[0].label[1] 
	,\labels[0].label[0] ,\labels[0].delimiter_valid[0] 
	,\labels[0].delimiter[7] ,\labels[0].delimiter[6] 
	,\labels[0].delimiter[5] ,\labels[0].delimiter[4] 
	,\labels[0].delimiter[3] ,\labels[0].delimiter[2] 
	,\labels[0].delimiter[1] ,\labels[0].delimiter[0] ;
output seed0_valid;
output [255:0] seed0_internal_state_key;
output [127:0] seed0_internal_state_value;
output [47:0] seed0_reseed_interval;
output seed1_valid;
output [255:0] seed1_internal_state_key;
output [127:0] seed1_internal_state_value;
output [47:0] seed1_reseed_interval;
output [8:0] \tready_override.r.part0 ;
wire \tready_override.f.txc_tready_override ;
wire \tready_override.f.engine_7_tready_override ;
wire \tready_override.f.engine_6_tready_override ;
wire \tready_override.f.engine_5_tready_override ;
wire \tready_override.f.engine_4_tready_override ;
wire \tready_override.f.engine_3_tready_override ;
wire \tready_override.f.engine_2_tready_override ;
wire \tready_override.f.engine_1_tready_override ;
wire \tready_override.f.engine_0_tready_override ;
wire [8:0] tready_override;
output [6:0] \cceip_encrypt_kop_fifo_override.r.part0 ;
wire \cceip_encrypt_kop_fifo_override.f.gcm_status_data_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.tlv_sb_data_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.kdf_cmd_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.kdfstream_cmd_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.keyfilter_cmd_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.gcm_tag_data_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.gcm_cmd_fifo ;
wire [6:0] cceip_encrypt_kop_fifo_override;
output [6:0] \cceip_validate_kop_fifo_override.r.part0 ;
wire \cceip_validate_kop_fifo_override.f.gcm_status_data_fifo ;
wire \cceip_validate_kop_fifo_override.f.tlv_sb_data_fifo ;
wire \cceip_validate_kop_fifo_override.f.kdf_cmd_fifo ;
wire \cceip_validate_kop_fifo_override.f.kdfstream_cmd_fifo ;
wire \cceip_validate_kop_fifo_override.f.keyfilter_cmd_fifo ;
wire \cceip_validate_kop_fifo_override.f.gcm_tag_data_fifo ;
wire \cceip_validate_kop_fifo_override.f.gcm_cmd_fifo ;
wire [6:0] cceip_validate_kop_fifo_override;
output [6:0] \cddip_decrypt_kop_fifo_override.r.part0 ;
wire \cddip_decrypt_kop_fifo_override.f.gcm_status_data_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.tlv_sb_data_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.kdf_cmd_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.kdfstream_cmd_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.keyfilter_cmd_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.gcm_tag_data_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.gcm_cmd_fifo ;
wire [6:0] cddip_decrypt_kop_fifo_override;
output manual_txc;
output always_validate_kim_ref;
output kdf_test_mode_en;
output [31:0] kdf_test_key_size;
output [31:0] \sa_global_ctrl.r.part0 ;
wire [29:0] \sa_global_ctrl.f.spare ;
wire \sa_global_ctrl.f.sa_snap ;
wire \sa_global_ctrl.f.sa_clear_live ;
wire [31:0] sa_global_ctrl;
output \sa_ctrl[31].r.part0[31] ,\sa_ctrl[31].r.part0[30] 
	,\sa_ctrl[31].r.part0[29] ,\sa_ctrl[31].r.part0[28] 
	,\sa_ctrl[31].r.part0[27] ,\sa_ctrl[31].r.part0[26] 
	,\sa_ctrl[31].r.part0[25] ,\sa_ctrl[31].r.part0[24] 
	,\sa_ctrl[31].r.part0[23] ,\sa_ctrl[31].r.part0[22] 
	,\sa_ctrl[31].r.part0[21] ,\sa_ctrl[31].r.part0[20] 
	,\sa_ctrl[31].r.part0[19] ,\sa_ctrl[31].r.part0[18] 
	,\sa_ctrl[31].r.part0[17] ,\sa_ctrl[31].r.part0[16] 
	,\sa_ctrl[31].r.part0[15] ,\sa_ctrl[31].r.part0[14] 
	,\sa_ctrl[31].r.part0[13] ,\sa_ctrl[31].r.part0[12] 
	,\sa_ctrl[31].r.part0[11] ,\sa_ctrl[31].r.part0[10] 
	,\sa_ctrl[31].r.part0[9] ,\sa_ctrl[31].r.part0[8] 
	,\sa_ctrl[31].r.part0[7] ,\sa_ctrl[31].r.part0[6] 
	,\sa_ctrl[31].r.part0[5] ,\sa_ctrl[31].r.part0[4] 
	,\sa_ctrl[31].r.part0[3] ,\sa_ctrl[31].r.part0[2] 
	,\sa_ctrl[31].r.part0[1] ,\sa_ctrl[31].r.part0[0] 
	,\sa_ctrl[30].r.part0[31] ,\sa_ctrl[30].r.part0[30] 
	,\sa_ctrl[30].r.part0[29] ,\sa_ctrl[30].r.part0[28] 
	,\sa_ctrl[30].r.part0[27] ,\sa_ctrl[30].r.part0[26] 
	,\sa_ctrl[30].r.part0[25] ,\sa_ctrl[30].r.part0[24] 
	,\sa_ctrl[30].r.part0[23] ,\sa_ctrl[30].r.part0[22] 
	,\sa_ctrl[30].r.part0[21] ,\sa_ctrl[30].r.part0[20] 
	,\sa_ctrl[30].r.part0[19] ,\sa_ctrl[30].r.part0[18] 
	,\sa_ctrl[30].r.part0[17] ,\sa_ctrl[30].r.part0[16] 
	,\sa_ctrl[30].r.part0[15] ,\sa_ctrl[30].r.part0[14] 
	,\sa_ctrl[30].r.part0[13] ,\sa_ctrl[30].r.part0[12] 
	,\sa_ctrl[30].r.part0[11] ,\sa_ctrl[30].r.part0[10] 
	,\sa_ctrl[30].r.part0[9] ,\sa_ctrl[30].r.part0[8] 
	,\sa_ctrl[30].r.part0[7] ,\sa_ctrl[30].r.part0[6] 
	,\sa_ctrl[30].r.part0[5] ,\sa_ctrl[30].r.part0[4] 
	,\sa_ctrl[30].r.part0[3] ,\sa_ctrl[30].r.part0[2] 
	,\sa_ctrl[30].r.part0[1] ,\sa_ctrl[30].r.part0[0] 
	,\sa_ctrl[29].r.part0[31] ,\sa_ctrl[29].r.part0[30] 
	,\sa_ctrl[29].r.part0[29] ,\sa_ctrl[29].r.part0[28] 
	,\sa_ctrl[29].r.part0[27] ,\sa_ctrl[29].r.part0[26] 
	,\sa_ctrl[29].r.part0[25] ,\sa_ctrl[29].r.part0[24] 
	,\sa_ctrl[29].r.part0[23] ,\sa_ctrl[29].r.part0[22] 
	,\sa_ctrl[29].r.part0[21] ,\sa_ctrl[29].r.part0[20] 
	,\sa_ctrl[29].r.part0[19] ,\sa_ctrl[29].r.part0[18] 
	,\sa_ctrl[29].r.part0[17] ,\sa_ctrl[29].r.part0[16] 
	,\sa_ctrl[29].r.part0[15] ,\sa_ctrl[29].r.part0[14] 
	,\sa_ctrl[29].r.part0[13] ,\sa_ctrl[29].r.part0[12] 
	,\sa_ctrl[29].r.part0[11] ,\sa_ctrl[29].r.part0[10] 
	,\sa_ctrl[29].r.part0[9] ,\sa_ctrl[29].r.part0[8] 
	,\sa_ctrl[29].r.part0[7] ,\sa_ctrl[29].r.part0[6] 
	,\sa_ctrl[29].r.part0[5] ,\sa_ctrl[29].r.part0[4] 
	,\sa_ctrl[29].r.part0[3] ,\sa_ctrl[29].r.part0[2] 
	,\sa_ctrl[29].r.part0[1] ,\sa_ctrl[29].r.part0[0] 
	,\sa_ctrl[28].r.part0[31] ,\sa_ctrl[28].r.part0[30] 
	,\sa_ctrl[28].r.part0[29] ,\sa_ctrl[28].r.part0[28] 
	,\sa_ctrl[28].r.part0[27] ,\sa_ctrl[28].r.part0[26] 
	,\sa_ctrl[28].r.part0[25] ,\sa_ctrl[28].r.part0[24] 
	,\sa_ctrl[28].r.part0[23] ,\sa_ctrl[28].r.part0[22] 
	,\sa_ctrl[28].r.part0[21] ,\sa_ctrl[28].r.part0[20] 
	,\sa_ctrl[28].r.part0[19] ,\sa_ctrl[28].r.part0[18] 
	,\sa_ctrl[28].r.part0[17] ,\sa_ctrl[28].r.part0[16] 
	,\sa_ctrl[28].r.part0[15] ,\sa_ctrl[28].r.part0[14] 
	,\sa_ctrl[28].r.part0[13] ,\sa_ctrl[28].r.part0[12] 
	,\sa_ctrl[28].r.part0[11] ,\sa_ctrl[28].r.part0[10] 
	,\sa_ctrl[28].r.part0[9] ,\sa_ctrl[28].r.part0[8] 
	,\sa_ctrl[28].r.part0[7] ,\sa_ctrl[28].r.part0[6] 
	,\sa_ctrl[28].r.part0[5] ,\sa_ctrl[28].r.part0[4] 
	,\sa_ctrl[28].r.part0[3] ,\sa_ctrl[28].r.part0[2] 
	,\sa_ctrl[28].r.part0[1] ,\sa_ctrl[28].r.part0[0] 
	,\sa_ctrl[27].r.part0[31] ,\sa_ctrl[27].r.part0[30] 
	,\sa_ctrl[27].r.part0[29] ,\sa_ctrl[27].r.part0[28] 
	,\sa_ctrl[27].r.part0[27] ,\sa_ctrl[27].r.part0[26] 
	,\sa_ctrl[27].r.part0[25] ,\sa_ctrl[27].r.part0[24] 
	,\sa_ctrl[27].r.part0[23] ,\sa_ctrl[27].r.part0[22] 
	,\sa_ctrl[27].r.part0[21] ,\sa_ctrl[27].r.part0[20] 
	,\sa_ctrl[27].r.part0[19] ,\sa_ctrl[27].r.part0[18] 
	,\sa_ctrl[27].r.part0[17] ,\sa_ctrl[27].r.part0[16] 
	,\sa_ctrl[27].r.part0[15] ,\sa_ctrl[27].r.part0[14] 
	,\sa_ctrl[27].r.part0[13] ,\sa_ctrl[27].r.part0[12] 
	,\sa_ctrl[27].r.part0[11] ,\sa_ctrl[27].r.part0[10] 
	,\sa_ctrl[27].r.part0[9] ,\sa_ctrl[27].r.part0[8] 
	,\sa_ctrl[27].r.part0[7] ,\sa_ctrl[27].r.part0[6] 
	,\sa_ctrl[27].r.part0[5] ,\sa_ctrl[27].r.part0[4] 
	,\sa_ctrl[27].r.part0[3] ,\sa_ctrl[27].r.part0[2] 
	,\sa_ctrl[27].r.part0[1] ,\sa_ctrl[27].r.part0[0] 
	,\sa_ctrl[26].r.part0[31] ,\sa_ctrl[26].r.part0[30] 
	,\sa_ctrl[26].r.part0[29] ,\sa_ctrl[26].r.part0[28] 
	,\sa_ctrl[26].r.part0[27] ,\sa_ctrl[26].r.part0[26] 
	,\sa_ctrl[26].r.part0[25] ,\sa_ctrl[26].r.part0[24] 
	,\sa_ctrl[26].r.part0[23] ,\sa_ctrl[26].r.part0[22] 
	,\sa_ctrl[26].r.part0[21] ,\sa_ctrl[26].r.part0[20] 
	,\sa_ctrl[26].r.part0[19] ,\sa_ctrl[26].r.part0[18] 
	,\sa_ctrl[26].r.part0[17] ,\sa_ctrl[26].r.part0[16] 
	,\sa_ctrl[26].r.part0[15] ,\sa_ctrl[26].r.part0[14] 
	,\sa_ctrl[26].r.part0[13] ,\sa_ctrl[26].r.part0[12] 
	,\sa_ctrl[26].r.part0[11] ,\sa_ctrl[26].r.part0[10] 
	,\sa_ctrl[26].r.part0[9] ,\sa_ctrl[26].r.part0[8] 
	,\sa_ctrl[26].r.part0[7] ,\sa_ctrl[26].r.part0[6] 
	,\sa_ctrl[26].r.part0[5] ,\sa_ctrl[26].r.part0[4] 
	,\sa_ctrl[26].r.part0[3] ,\sa_ctrl[26].r.part0[2] 
	,\sa_ctrl[26].r.part0[1] ,\sa_ctrl[26].r.part0[0] 
	,\sa_ctrl[25].r.part0[31] ,\sa_ctrl[25].r.part0[30] 
	,\sa_ctrl[25].r.part0[29] ,\sa_ctrl[25].r.part0[28] 
	,\sa_ctrl[25].r.part0[27] ,\sa_ctrl[25].r.part0[26] 
	,\sa_ctrl[25].r.part0[25] ,\sa_ctrl[25].r.part0[24] 
	,\sa_ctrl[25].r.part0[23] ,\sa_ctrl[25].r.part0[22] 
	,\sa_ctrl[25].r.part0[21] ,\sa_ctrl[25].r.part0[20] 
	,\sa_ctrl[25].r.part0[19] ,\sa_ctrl[25].r.part0[18] 
	,\sa_ctrl[25].r.part0[17] ,\sa_ctrl[25].r.part0[16] 
	,\sa_ctrl[25].r.part0[15] ,\sa_ctrl[25].r.part0[14] 
	,\sa_ctrl[25].r.part0[13] ,\sa_ctrl[25].r.part0[12] 
	,\sa_ctrl[25].r.part0[11] ,\sa_ctrl[25].r.part0[10] 
	,\sa_ctrl[25].r.part0[9] ,\sa_ctrl[25].r.part0[8] 
	,\sa_ctrl[25].r.part0[7] ,\sa_ctrl[25].r.part0[6] 
	,\sa_ctrl[25].r.part0[5] ,\sa_ctrl[25].r.part0[4] 
	,\sa_ctrl[25].r.part0[3] ,\sa_ctrl[25].r.part0[2] 
	,\sa_ctrl[25].r.part0[1] ,\sa_ctrl[25].r.part0[0] 
	,\sa_ctrl[24].r.part0[31] ,\sa_ctrl[24].r.part0[30] 
	,\sa_ctrl[24].r.part0[29] ,\sa_ctrl[24].r.part0[28] 
	,\sa_ctrl[24].r.part0[27] ,\sa_ctrl[24].r.part0[26] 
	,\sa_ctrl[24].r.part0[25] ,\sa_ctrl[24].r.part0[24] 
	,\sa_ctrl[24].r.part0[23] ,\sa_ctrl[24].r.part0[22] 
	,\sa_ctrl[24].r.part0[21] ,\sa_ctrl[24].r.part0[20] 
	,\sa_ctrl[24].r.part0[19] ,\sa_ctrl[24].r.part0[18] 
	,\sa_ctrl[24].r.part0[17] ,\sa_ctrl[24].r.part0[16] 
	,\sa_ctrl[24].r.part0[15] ,\sa_ctrl[24].r.part0[14] 
	,\sa_ctrl[24].r.part0[13] ,\sa_ctrl[24].r.part0[12] 
	,\sa_ctrl[24].r.part0[11] ,\sa_ctrl[24].r.part0[10] 
	,\sa_ctrl[24].r.part0[9] ,\sa_ctrl[24].r.part0[8] 
	,\sa_ctrl[24].r.part0[7] ,\sa_ctrl[24].r.part0[6] 
	,\sa_ctrl[24].r.part0[5] ,\sa_ctrl[24].r.part0[4] 
	,\sa_ctrl[24].r.part0[3] ,\sa_ctrl[24].r.part0[2] 
	,\sa_ctrl[24].r.part0[1] ,\sa_ctrl[24].r.part0[0] 
	,\sa_ctrl[23].r.part0[31] ,\sa_ctrl[23].r.part0[30] 
	,\sa_ctrl[23].r.part0[29] ,\sa_ctrl[23].r.part0[28] 
	,\sa_ctrl[23].r.part0[27] ,\sa_ctrl[23].r.part0[26] 
	,\sa_ctrl[23].r.part0[25] ,\sa_ctrl[23].r.part0[24] 
	,\sa_ctrl[23].r.part0[23] ,\sa_ctrl[23].r.part0[22] 
	,\sa_ctrl[23].r.part0[21] ,\sa_ctrl[23].r.part0[20] 
	,\sa_ctrl[23].r.part0[19] ,\sa_ctrl[23].r.part0[18] 
	,\sa_ctrl[23].r.part0[17] ,\sa_ctrl[23].r.part0[16] 
	,\sa_ctrl[23].r.part0[15] ,\sa_ctrl[23].r.part0[14] 
	,\sa_ctrl[23].r.part0[13] ,\sa_ctrl[23].r.part0[12] 
	,\sa_ctrl[23].r.part0[11] ,\sa_ctrl[23].r.part0[10] 
	,\sa_ctrl[23].r.part0[9] ,\sa_ctrl[23].r.part0[8] 
	,\sa_ctrl[23].r.part0[7] ,\sa_ctrl[23].r.part0[6] 
	,\sa_ctrl[23].r.part0[5] ,\sa_ctrl[23].r.part0[4] 
	,\sa_ctrl[23].r.part0[3] ,\sa_ctrl[23].r.part0[2] 
	,\sa_ctrl[23].r.part0[1] ,\sa_ctrl[23].r.part0[0] 
	,\sa_ctrl[22].r.part0[31] ,\sa_ctrl[22].r.part0[30] 
	,\sa_ctrl[22].r.part0[29] ,\sa_ctrl[22].r.part0[28] 
	,\sa_ctrl[22].r.part0[27] ,\sa_ctrl[22].r.part0[26] 
	,\sa_ctrl[22].r.part0[25] ,\sa_ctrl[22].r.part0[24] 
	,\sa_ctrl[22].r.part0[23] ,\sa_ctrl[22].r.part0[22] 
	,\sa_ctrl[22].r.part0[21] ,\sa_ctrl[22].r.part0[20] 
	,\sa_ctrl[22].r.part0[19] ,\sa_ctrl[22].r.part0[18] 
	,\sa_ctrl[22].r.part0[17] ,\sa_ctrl[22].r.part0[16] 
	,\sa_ctrl[22].r.part0[15] ,\sa_ctrl[22].r.part0[14] 
	,\sa_ctrl[22].r.part0[13] ,\sa_ctrl[22].r.part0[12] 
	,\sa_ctrl[22].r.part0[11] ,\sa_ctrl[22].r.part0[10] 
	,\sa_ctrl[22].r.part0[9] ,\sa_ctrl[22].r.part0[8] 
	,\sa_ctrl[22].r.part0[7] ,\sa_ctrl[22].r.part0[6] 
	,\sa_ctrl[22].r.part0[5] ,\sa_ctrl[22].r.part0[4] 
	,\sa_ctrl[22].r.part0[3] ,\sa_ctrl[22].r.part0[2] 
	,\sa_ctrl[22].r.part0[1] ,\sa_ctrl[22].r.part0[0] 
	,\sa_ctrl[21].r.part0[31] ,\sa_ctrl[21].r.part0[30] 
	,\sa_ctrl[21].r.part0[29] ,\sa_ctrl[21].r.part0[28] 
	,\sa_ctrl[21].r.part0[27] ,\sa_ctrl[21].r.part0[26] 
	,\sa_ctrl[21].r.part0[25] ,\sa_ctrl[21].r.part0[24] 
	,\sa_ctrl[21].r.part0[23] ,\sa_ctrl[21].r.part0[22] 
	,\sa_ctrl[21].r.part0[21] ,\sa_ctrl[21].r.part0[20] 
	,\sa_ctrl[21].r.part0[19] ,\sa_ctrl[21].r.part0[18] 
	,\sa_ctrl[21].r.part0[17] ,\sa_ctrl[21].r.part0[16] 
	,\sa_ctrl[21].r.part0[15] ,\sa_ctrl[21].r.part0[14] 
	,\sa_ctrl[21].r.part0[13] ,\sa_ctrl[21].r.part0[12] 
	,\sa_ctrl[21].r.part0[11] ,\sa_ctrl[21].r.part0[10] 
	,\sa_ctrl[21].r.part0[9] ,\sa_ctrl[21].r.part0[8] 
	,\sa_ctrl[21].r.part0[7] ,\sa_ctrl[21].r.part0[6] 
	,\sa_ctrl[21].r.part0[5] ,\sa_ctrl[21].r.part0[4] 
	,\sa_ctrl[21].r.part0[3] ,\sa_ctrl[21].r.part0[2] 
	,\sa_ctrl[21].r.part0[1] ,\sa_ctrl[21].r.part0[0] 
	,\sa_ctrl[20].r.part0[31] ,\sa_ctrl[20].r.part0[30] 
	,\sa_ctrl[20].r.part0[29] ,\sa_ctrl[20].r.part0[28] 
	,\sa_ctrl[20].r.part0[27] ,\sa_ctrl[20].r.part0[26] 
	,\sa_ctrl[20].r.part0[25] ,\sa_ctrl[20].r.part0[24] 
	,\sa_ctrl[20].r.part0[23] ,\sa_ctrl[20].r.part0[22] 
	,\sa_ctrl[20].r.part0[21] ,\sa_ctrl[20].r.part0[20] 
	,\sa_ctrl[20].r.part0[19] ,\sa_ctrl[20].r.part0[18] 
	,\sa_ctrl[20].r.part0[17] ,\sa_ctrl[20].r.part0[16] 
	,\sa_ctrl[20].r.part0[15] ,\sa_ctrl[20].r.part0[14] 
	,\sa_ctrl[20].r.part0[13] ,\sa_ctrl[20].r.part0[12] 
	,\sa_ctrl[20].r.part0[11] ,\sa_ctrl[20].r.part0[10] 
	,\sa_ctrl[20].r.part0[9] ,\sa_ctrl[20].r.part0[8] 
	,\sa_ctrl[20].r.part0[7] ,\sa_ctrl[20].r.part0[6] 
	,\sa_ctrl[20].r.part0[5] ,\sa_ctrl[20].r.part0[4] 
	,\sa_ctrl[20].r.part0[3] ,\sa_ctrl[20].r.part0[2] 
	,\sa_ctrl[20].r.part0[1] ,\sa_ctrl[20].r.part0[0] 
	,\sa_ctrl[19].r.part0[31] ,\sa_ctrl[19].r.part0[30] 
	,\sa_ctrl[19].r.part0[29] ,\sa_ctrl[19].r.part0[28] 
	,\sa_ctrl[19].r.part0[27] ,\sa_ctrl[19].r.part0[26] 
	,\sa_ctrl[19].r.part0[25] ,\sa_ctrl[19].r.part0[24] 
	,\sa_ctrl[19].r.part0[23] ,\sa_ctrl[19].r.part0[22] 
	,\sa_ctrl[19].r.part0[21] ,\sa_ctrl[19].r.part0[20] 
	,\sa_ctrl[19].r.part0[19] ,\sa_ctrl[19].r.part0[18] 
	,\sa_ctrl[19].r.part0[17] ,\sa_ctrl[19].r.part0[16] 
	,\sa_ctrl[19].r.part0[15] ,\sa_ctrl[19].r.part0[14] 
	,\sa_ctrl[19].r.part0[13] ,\sa_ctrl[19].r.part0[12] 
	,\sa_ctrl[19].r.part0[11] ,\sa_ctrl[19].r.part0[10] 
	,\sa_ctrl[19].r.part0[9] ,\sa_ctrl[19].r.part0[8] 
	,\sa_ctrl[19].r.part0[7] ,\sa_ctrl[19].r.part0[6] 
	,\sa_ctrl[19].r.part0[5] ,\sa_ctrl[19].r.part0[4] 
	,\sa_ctrl[19].r.part0[3] ,\sa_ctrl[19].r.part0[2] 
	,\sa_ctrl[19].r.part0[1] ,\sa_ctrl[19].r.part0[0] 
	,\sa_ctrl[18].r.part0[31] ,\sa_ctrl[18].r.part0[30] 
	,\sa_ctrl[18].r.part0[29] ,\sa_ctrl[18].r.part0[28] 
	,\sa_ctrl[18].r.part0[27] ,\sa_ctrl[18].r.part0[26] 
	,\sa_ctrl[18].r.part0[25] ,\sa_ctrl[18].r.part0[24] 
	,\sa_ctrl[18].r.part0[23] ,\sa_ctrl[18].r.part0[22] 
	,\sa_ctrl[18].r.part0[21] ,\sa_ctrl[18].r.part0[20] 
	,\sa_ctrl[18].r.part0[19] ,\sa_ctrl[18].r.part0[18] 
	,\sa_ctrl[18].r.part0[17] ,\sa_ctrl[18].r.part0[16] 
	,\sa_ctrl[18].r.part0[15] ,\sa_ctrl[18].r.part0[14] 
	,\sa_ctrl[18].r.part0[13] ,\sa_ctrl[18].r.part0[12] 
	,\sa_ctrl[18].r.part0[11] ,\sa_ctrl[18].r.part0[10] 
	,\sa_ctrl[18].r.part0[9] ,\sa_ctrl[18].r.part0[8] 
	,\sa_ctrl[18].r.part0[7] ,\sa_ctrl[18].r.part0[6] 
	,\sa_ctrl[18].r.part0[5] ,\sa_ctrl[18].r.part0[4] 
	,\sa_ctrl[18].r.part0[3] ,\sa_ctrl[18].r.part0[2] 
	,\sa_ctrl[18].r.part0[1] ,\sa_ctrl[18].r.part0[0] 
	,\sa_ctrl[17].r.part0[31] ,\sa_ctrl[17].r.part0[30] 
	,\sa_ctrl[17].r.part0[29] ,\sa_ctrl[17].r.part0[28] 
	,\sa_ctrl[17].r.part0[27] ,\sa_ctrl[17].r.part0[26] 
	,\sa_ctrl[17].r.part0[25] ,\sa_ctrl[17].r.part0[24] 
	,\sa_ctrl[17].r.part0[23] ,\sa_ctrl[17].r.part0[22] 
	,\sa_ctrl[17].r.part0[21] ,\sa_ctrl[17].r.part0[20] 
	,\sa_ctrl[17].r.part0[19] ,\sa_ctrl[17].r.part0[18] 
	,\sa_ctrl[17].r.part0[17] ,\sa_ctrl[17].r.part0[16] 
	,\sa_ctrl[17].r.part0[15] ,\sa_ctrl[17].r.part0[14] 
	,\sa_ctrl[17].r.part0[13] ,\sa_ctrl[17].r.part0[12] 
	,\sa_ctrl[17].r.part0[11] ,\sa_ctrl[17].r.part0[10] 
	,\sa_ctrl[17].r.part0[9] ,\sa_ctrl[17].r.part0[8] 
	,\sa_ctrl[17].r.part0[7] ,\sa_ctrl[17].r.part0[6] 
	,\sa_ctrl[17].r.part0[5] ,\sa_ctrl[17].r.part0[4] 
	,\sa_ctrl[17].r.part0[3] ,\sa_ctrl[17].r.part0[2] 
	,\sa_ctrl[17].r.part0[1] ,\sa_ctrl[17].r.part0[0] 
	,\sa_ctrl[16].r.part0[31] ,\sa_ctrl[16].r.part0[30] 
	,\sa_ctrl[16].r.part0[29] ,\sa_ctrl[16].r.part0[28] 
	,\sa_ctrl[16].r.part0[27] ,\sa_ctrl[16].r.part0[26] 
	,\sa_ctrl[16].r.part0[25] ,\sa_ctrl[16].r.part0[24] 
	,\sa_ctrl[16].r.part0[23] ,\sa_ctrl[16].r.part0[22] 
	,\sa_ctrl[16].r.part0[21] ,\sa_ctrl[16].r.part0[20] 
	,\sa_ctrl[16].r.part0[19] ,\sa_ctrl[16].r.part0[18] 
	,\sa_ctrl[16].r.part0[17] ,\sa_ctrl[16].r.part0[16] 
	,\sa_ctrl[16].r.part0[15] ,\sa_ctrl[16].r.part0[14] 
	,\sa_ctrl[16].r.part0[13] ,\sa_ctrl[16].r.part0[12] 
	,\sa_ctrl[16].r.part0[11] ,\sa_ctrl[16].r.part0[10] 
	,\sa_ctrl[16].r.part0[9] ,\sa_ctrl[16].r.part0[8] 
	,\sa_ctrl[16].r.part0[7] ,\sa_ctrl[16].r.part0[6] 
	,\sa_ctrl[16].r.part0[5] ,\sa_ctrl[16].r.part0[4] 
	,\sa_ctrl[16].r.part0[3] ,\sa_ctrl[16].r.part0[2] 
	,\sa_ctrl[16].r.part0[1] ,\sa_ctrl[16].r.part0[0] 
	,\sa_ctrl[15].r.part0[31] ,\sa_ctrl[15].r.part0[30] 
	,\sa_ctrl[15].r.part0[29] ,\sa_ctrl[15].r.part0[28] 
	,\sa_ctrl[15].r.part0[27] ,\sa_ctrl[15].r.part0[26] 
	,\sa_ctrl[15].r.part0[25] ,\sa_ctrl[15].r.part0[24] 
	,\sa_ctrl[15].r.part0[23] ,\sa_ctrl[15].r.part0[22] 
	,\sa_ctrl[15].r.part0[21] ,\sa_ctrl[15].r.part0[20] 
	,\sa_ctrl[15].r.part0[19] ,\sa_ctrl[15].r.part0[18] 
	,\sa_ctrl[15].r.part0[17] ,\sa_ctrl[15].r.part0[16] 
	,\sa_ctrl[15].r.part0[15] ,\sa_ctrl[15].r.part0[14] 
	,\sa_ctrl[15].r.part0[13] ,\sa_ctrl[15].r.part0[12] 
	,\sa_ctrl[15].r.part0[11] ,\sa_ctrl[15].r.part0[10] 
	,\sa_ctrl[15].r.part0[9] ,\sa_ctrl[15].r.part0[8] 
	,\sa_ctrl[15].r.part0[7] ,\sa_ctrl[15].r.part0[6] 
	,\sa_ctrl[15].r.part0[5] ,\sa_ctrl[15].r.part0[4] 
	,\sa_ctrl[15].r.part0[3] ,\sa_ctrl[15].r.part0[2] 
	,\sa_ctrl[15].r.part0[1] ,\sa_ctrl[15].r.part0[0] 
	,\sa_ctrl[14].r.part0[31] ,\sa_ctrl[14].r.part0[30] 
	,\sa_ctrl[14].r.part0[29] ,\sa_ctrl[14].r.part0[28] 
	,\sa_ctrl[14].r.part0[27] ,\sa_ctrl[14].r.part0[26] 
	,\sa_ctrl[14].r.part0[25] ,\sa_ctrl[14].r.part0[24] 
	,\sa_ctrl[14].r.part0[23] ,\sa_ctrl[14].r.part0[22] 
	,\sa_ctrl[14].r.part0[21] ,\sa_ctrl[14].r.part0[20] 
	,\sa_ctrl[14].r.part0[19] ,\sa_ctrl[14].r.part0[18] 
	,\sa_ctrl[14].r.part0[17] ,\sa_ctrl[14].r.part0[16] 
	,\sa_ctrl[14].r.part0[15] ,\sa_ctrl[14].r.part0[14] 
	,\sa_ctrl[14].r.part0[13] ,\sa_ctrl[14].r.part0[12] 
	,\sa_ctrl[14].r.part0[11] ,\sa_ctrl[14].r.part0[10] 
	,\sa_ctrl[14].r.part0[9] ,\sa_ctrl[14].r.part0[8] 
	,\sa_ctrl[14].r.part0[7] ,\sa_ctrl[14].r.part0[6] 
	,\sa_ctrl[14].r.part0[5] ,\sa_ctrl[14].r.part0[4] 
	,\sa_ctrl[14].r.part0[3] ,\sa_ctrl[14].r.part0[2] 
	,\sa_ctrl[14].r.part0[1] ,\sa_ctrl[14].r.part0[0] 
	,\sa_ctrl[13].r.part0[31] ,\sa_ctrl[13].r.part0[30] 
	,\sa_ctrl[13].r.part0[29] ,\sa_ctrl[13].r.part0[28] 
	,\sa_ctrl[13].r.part0[27] ,\sa_ctrl[13].r.part0[26] 
	,\sa_ctrl[13].r.part0[25] ,\sa_ctrl[13].r.part0[24] 
	,\sa_ctrl[13].r.part0[23] ,\sa_ctrl[13].r.part0[22] 
	,\sa_ctrl[13].r.part0[21] ,\sa_ctrl[13].r.part0[20] 
	,\sa_ctrl[13].r.part0[19] ,\sa_ctrl[13].r.part0[18] 
	,\sa_ctrl[13].r.part0[17] ,\sa_ctrl[13].r.part0[16] 
	,\sa_ctrl[13].r.part0[15] ,\sa_ctrl[13].r.part0[14] 
	,\sa_ctrl[13].r.part0[13] ,\sa_ctrl[13].r.part0[12] 
	,\sa_ctrl[13].r.part0[11] ,\sa_ctrl[13].r.part0[10] 
	,\sa_ctrl[13].r.part0[9] ,\sa_ctrl[13].r.part0[8] 
	,\sa_ctrl[13].r.part0[7] ,\sa_ctrl[13].r.part0[6] 
	,\sa_ctrl[13].r.part0[5] ,\sa_ctrl[13].r.part0[4] 
	,\sa_ctrl[13].r.part0[3] ,\sa_ctrl[13].r.part0[2] 
	,\sa_ctrl[13].r.part0[1] ,\sa_ctrl[13].r.part0[0] 
	,\sa_ctrl[12].r.part0[31] ,\sa_ctrl[12].r.part0[30] 
	,\sa_ctrl[12].r.part0[29] ,\sa_ctrl[12].r.part0[28] 
	,\sa_ctrl[12].r.part0[27] ,\sa_ctrl[12].r.part0[26] 
	,\sa_ctrl[12].r.part0[25] ,\sa_ctrl[12].r.part0[24] 
	,\sa_ctrl[12].r.part0[23] ,\sa_ctrl[12].r.part0[22] 
	,\sa_ctrl[12].r.part0[21] ,\sa_ctrl[12].r.part0[20] 
	,\sa_ctrl[12].r.part0[19] ,\sa_ctrl[12].r.part0[18] 
	,\sa_ctrl[12].r.part0[17] ,\sa_ctrl[12].r.part0[16] 
	,\sa_ctrl[12].r.part0[15] ,\sa_ctrl[12].r.part0[14] 
	,\sa_ctrl[12].r.part0[13] ,\sa_ctrl[12].r.part0[12] 
	,\sa_ctrl[12].r.part0[11] ,\sa_ctrl[12].r.part0[10] 
	,\sa_ctrl[12].r.part0[9] ,\sa_ctrl[12].r.part0[8] 
	,\sa_ctrl[12].r.part0[7] ,\sa_ctrl[12].r.part0[6] 
	,\sa_ctrl[12].r.part0[5] ,\sa_ctrl[12].r.part0[4] 
	,\sa_ctrl[12].r.part0[3] ,\sa_ctrl[12].r.part0[2] 
	,\sa_ctrl[12].r.part0[1] ,\sa_ctrl[12].r.part0[0] 
	,\sa_ctrl[11].r.part0[31] ,\sa_ctrl[11].r.part0[30] 
	,\sa_ctrl[11].r.part0[29] ,\sa_ctrl[11].r.part0[28] 
	,\sa_ctrl[11].r.part0[27] ,\sa_ctrl[11].r.part0[26] 
	,\sa_ctrl[11].r.part0[25] ,\sa_ctrl[11].r.part0[24] 
	,\sa_ctrl[11].r.part0[23] ,\sa_ctrl[11].r.part0[22] 
	,\sa_ctrl[11].r.part0[21] ,\sa_ctrl[11].r.part0[20] 
	,\sa_ctrl[11].r.part0[19] ,\sa_ctrl[11].r.part0[18] 
	,\sa_ctrl[11].r.part0[17] ,\sa_ctrl[11].r.part0[16] 
	,\sa_ctrl[11].r.part0[15] ,\sa_ctrl[11].r.part0[14] 
	,\sa_ctrl[11].r.part0[13] ,\sa_ctrl[11].r.part0[12] 
	,\sa_ctrl[11].r.part0[11] ,\sa_ctrl[11].r.part0[10] 
	,\sa_ctrl[11].r.part0[9] ,\sa_ctrl[11].r.part0[8] 
	,\sa_ctrl[11].r.part0[7] ,\sa_ctrl[11].r.part0[6] 
	,\sa_ctrl[11].r.part0[5] ,\sa_ctrl[11].r.part0[4] 
	,\sa_ctrl[11].r.part0[3] ,\sa_ctrl[11].r.part0[2] 
	,\sa_ctrl[11].r.part0[1] ,\sa_ctrl[11].r.part0[0] 
	,\sa_ctrl[10].r.part0[31] ,\sa_ctrl[10].r.part0[30] 
	,\sa_ctrl[10].r.part0[29] ,\sa_ctrl[10].r.part0[28] 
	,\sa_ctrl[10].r.part0[27] ,\sa_ctrl[10].r.part0[26] 
	,\sa_ctrl[10].r.part0[25] ,\sa_ctrl[10].r.part0[24] 
	,\sa_ctrl[10].r.part0[23] ,\sa_ctrl[10].r.part0[22] 
	,\sa_ctrl[10].r.part0[21] ,\sa_ctrl[10].r.part0[20] 
	,\sa_ctrl[10].r.part0[19] ,\sa_ctrl[10].r.part0[18] 
	,\sa_ctrl[10].r.part0[17] ,\sa_ctrl[10].r.part0[16] 
	,\sa_ctrl[10].r.part0[15] ,\sa_ctrl[10].r.part0[14] 
	,\sa_ctrl[10].r.part0[13] ,\sa_ctrl[10].r.part0[12] 
	,\sa_ctrl[10].r.part0[11] ,\sa_ctrl[10].r.part0[10] 
	,\sa_ctrl[10].r.part0[9] ,\sa_ctrl[10].r.part0[8] 
	,\sa_ctrl[10].r.part0[7] ,\sa_ctrl[10].r.part0[6] 
	,\sa_ctrl[10].r.part0[5] ,\sa_ctrl[10].r.part0[4] 
	,\sa_ctrl[10].r.part0[3] ,\sa_ctrl[10].r.part0[2] 
	,\sa_ctrl[10].r.part0[1] ,\sa_ctrl[10].r.part0[0] 
	,\sa_ctrl[9].r.part0[31] ,\sa_ctrl[9].r.part0[30] 
	,\sa_ctrl[9].r.part0[29] ,\sa_ctrl[9].r.part0[28] 
	,\sa_ctrl[9].r.part0[27] ,\sa_ctrl[9].r.part0[26] 
	,\sa_ctrl[9].r.part0[25] ,\sa_ctrl[9].r.part0[24] 
	,\sa_ctrl[9].r.part0[23] ,\sa_ctrl[9].r.part0[22] 
	,\sa_ctrl[9].r.part0[21] ,\sa_ctrl[9].r.part0[20] 
	,\sa_ctrl[9].r.part0[19] ,\sa_ctrl[9].r.part0[18] 
	,\sa_ctrl[9].r.part0[17] ,\sa_ctrl[9].r.part0[16] 
	,\sa_ctrl[9].r.part0[15] ,\sa_ctrl[9].r.part0[14] 
	,\sa_ctrl[9].r.part0[13] ,\sa_ctrl[9].r.part0[12] 
	,\sa_ctrl[9].r.part0[11] ,\sa_ctrl[9].r.part0[10] 
	,\sa_ctrl[9].r.part0[9] ,\sa_ctrl[9].r.part0[8] 
	,\sa_ctrl[9].r.part0[7] ,\sa_ctrl[9].r.part0[6] 
	,\sa_ctrl[9].r.part0[5] ,\sa_ctrl[9].r.part0[4] 
	,\sa_ctrl[9].r.part0[3] ,\sa_ctrl[9].r.part0[2] 
	,\sa_ctrl[9].r.part0[1] ,\sa_ctrl[9].r.part0[0] 
	,\sa_ctrl[8].r.part0[31] ,\sa_ctrl[8].r.part0[30] 
	,\sa_ctrl[8].r.part0[29] ,\sa_ctrl[8].r.part0[28] 
	,\sa_ctrl[8].r.part0[27] ,\sa_ctrl[8].r.part0[26] 
	,\sa_ctrl[8].r.part0[25] ,\sa_ctrl[8].r.part0[24] 
	,\sa_ctrl[8].r.part0[23] ,\sa_ctrl[8].r.part0[22] 
	,\sa_ctrl[8].r.part0[21] ,\sa_ctrl[8].r.part0[20] 
	,\sa_ctrl[8].r.part0[19] ,\sa_ctrl[8].r.part0[18] 
	,\sa_ctrl[8].r.part0[17] ,\sa_ctrl[8].r.part0[16] 
	,\sa_ctrl[8].r.part0[15] ,\sa_ctrl[8].r.part0[14] 
	,\sa_ctrl[8].r.part0[13] ,\sa_ctrl[8].r.part0[12] 
	,\sa_ctrl[8].r.part0[11] ,\sa_ctrl[8].r.part0[10] 
	,\sa_ctrl[8].r.part0[9] ,\sa_ctrl[8].r.part0[8] 
	,\sa_ctrl[8].r.part0[7] ,\sa_ctrl[8].r.part0[6] 
	,\sa_ctrl[8].r.part0[5] ,\sa_ctrl[8].r.part0[4] 
	,\sa_ctrl[8].r.part0[3] ,\sa_ctrl[8].r.part0[2] 
	,\sa_ctrl[8].r.part0[1] ,\sa_ctrl[8].r.part0[0] 
	,\sa_ctrl[7].r.part0[31] ,\sa_ctrl[7].r.part0[30] 
	,\sa_ctrl[7].r.part0[29] ,\sa_ctrl[7].r.part0[28] 
	,\sa_ctrl[7].r.part0[27] ,\sa_ctrl[7].r.part0[26] 
	,\sa_ctrl[7].r.part0[25] ,\sa_ctrl[7].r.part0[24] 
	,\sa_ctrl[7].r.part0[23] ,\sa_ctrl[7].r.part0[22] 
	,\sa_ctrl[7].r.part0[21] ,\sa_ctrl[7].r.part0[20] 
	,\sa_ctrl[7].r.part0[19] ,\sa_ctrl[7].r.part0[18] 
	,\sa_ctrl[7].r.part0[17] ,\sa_ctrl[7].r.part0[16] 
	,\sa_ctrl[7].r.part0[15] ,\sa_ctrl[7].r.part0[14] 
	,\sa_ctrl[7].r.part0[13] ,\sa_ctrl[7].r.part0[12] 
	,\sa_ctrl[7].r.part0[11] ,\sa_ctrl[7].r.part0[10] 
	,\sa_ctrl[7].r.part0[9] ,\sa_ctrl[7].r.part0[8] 
	,\sa_ctrl[7].r.part0[7] ,\sa_ctrl[7].r.part0[6] 
	,\sa_ctrl[7].r.part0[5] ,\sa_ctrl[7].r.part0[4] 
	,\sa_ctrl[7].r.part0[3] ,\sa_ctrl[7].r.part0[2] 
	,\sa_ctrl[7].r.part0[1] ,\sa_ctrl[7].r.part0[0] 
	,\sa_ctrl[6].r.part0[31] ,\sa_ctrl[6].r.part0[30] 
	,\sa_ctrl[6].r.part0[29] ,\sa_ctrl[6].r.part0[28] 
	,\sa_ctrl[6].r.part0[27] ,\sa_ctrl[6].r.part0[26] 
	,\sa_ctrl[6].r.part0[25] ,\sa_ctrl[6].r.part0[24] 
	,\sa_ctrl[6].r.part0[23] ,\sa_ctrl[6].r.part0[22] 
	,\sa_ctrl[6].r.part0[21] ,\sa_ctrl[6].r.part0[20] 
	,\sa_ctrl[6].r.part0[19] ,\sa_ctrl[6].r.part0[18] 
	,\sa_ctrl[6].r.part0[17] ,\sa_ctrl[6].r.part0[16] 
	,\sa_ctrl[6].r.part0[15] ,\sa_ctrl[6].r.part0[14] 
	,\sa_ctrl[6].r.part0[13] ,\sa_ctrl[6].r.part0[12] 
	,\sa_ctrl[6].r.part0[11] ,\sa_ctrl[6].r.part0[10] 
	,\sa_ctrl[6].r.part0[9] ,\sa_ctrl[6].r.part0[8] 
	,\sa_ctrl[6].r.part0[7] ,\sa_ctrl[6].r.part0[6] 
	,\sa_ctrl[6].r.part0[5] ,\sa_ctrl[6].r.part0[4] 
	,\sa_ctrl[6].r.part0[3] ,\sa_ctrl[6].r.part0[2] 
	,\sa_ctrl[6].r.part0[1] ,\sa_ctrl[6].r.part0[0] 
	,\sa_ctrl[5].r.part0[31] ,\sa_ctrl[5].r.part0[30] 
	,\sa_ctrl[5].r.part0[29] ,\sa_ctrl[5].r.part0[28] 
	,\sa_ctrl[5].r.part0[27] ,\sa_ctrl[5].r.part0[26] 
	,\sa_ctrl[5].r.part0[25] ,\sa_ctrl[5].r.part0[24] 
	,\sa_ctrl[5].r.part0[23] ,\sa_ctrl[5].r.part0[22] 
	,\sa_ctrl[5].r.part0[21] ,\sa_ctrl[5].r.part0[20] 
	,\sa_ctrl[5].r.part0[19] ,\sa_ctrl[5].r.part0[18] 
	,\sa_ctrl[5].r.part0[17] ,\sa_ctrl[5].r.part0[16] 
	,\sa_ctrl[5].r.part0[15] ,\sa_ctrl[5].r.part0[14] 
	,\sa_ctrl[5].r.part0[13] ,\sa_ctrl[5].r.part0[12] 
	,\sa_ctrl[5].r.part0[11] ,\sa_ctrl[5].r.part0[10] 
	,\sa_ctrl[5].r.part0[9] ,\sa_ctrl[5].r.part0[8] 
	,\sa_ctrl[5].r.part0[7] ,\sa_ctrl[5].r.part0[6] 
	,\sa_ctrl[5].r.part0[5] ,\sa_ctrl[5].r.part0[4] 
	,\sa_ctrl[5].r.part0[3] ,\sa_ctrl[5].r.part0[2] 
	,\sa_ctrl[5].r.part0[1] ,\sa_ctrl[5].r.part0[0] 
	,\sa_ctrl[4].r.part0[31] ,\sa_ctrl[4].r.part0[30] 
	,\sa_ctrl[4].r.part0[29] ,\sa_ctrl[4].r.part0[28] 
	,\sa_ctrl[4].r.part0[27] ,\sa_ctrl[4].r.part0[26] 
	,\sa_ctrl[4].r.part0[25] ,\sa_ctrl[4].r.part0[24] 
	,\sa_ctrl[4].r.part0[23] ,\sa_ctrl[4].r.part0[22] 
	,\sa_ctrl[4].r.part0[21] ,\sa_ctrl[4].r.part0[20] 
	,\sa_ctrl[4].r.part0[19] ,\sa_ctrl[4].r.part0[18] 
	,\sa_ctrl[4].r.part0[17] ,\sa_ctrl[4].r.part0[16] 
	,\sa_ctrl[4].r.part0[15] ,\sa_ctrl[4].r.part0[14] 
	,\sa_ctrl[4].r.part0[13] ,\sa_ctrl[4].r.part0[12] 
	,\sa_ctrl[4].r.part0[11] ,\sa_ctrl[4].r.part0[10] 
	,\sa_ctrl[4].r.part0[9] ,\sa_ctrl[4].r.part0[8] 
	,\sa_ctrl[4].r.part0[7] ,\sa_ctrl[4].r.part0[6] 
	,\sa_ctrl[4].r.part0[5] ,\sa_ctrl[4].r.part0[4] 
	,\sa_ctrl[4].r.part0[3] ,\sa_ctrl[4].r.part0[2] 
	,\sa_ctrl[4].r.part0[1] ,\sa_ctrl[4].r.part0[0] 
	,\sa_ctrl[3].r.part0[31] ,\sa_ctrl[3].r.part0[30] 
	,\sa_ctrl[3].r.part0[29] ,\sa_ctrl[3].r.part0[28] 
	,\sa_ctrl[3].r.part0[27] ,\sa_ctrl[3].r.part0[26] 
	,\sa_ctrl[3].r.part0[25] ,\sa_ctrl[3].r.part0[24] 
	,\sa_ctrl[3].r.part0[23] ,\sa_ctrl[3].r.part0[22] 
	,\sa_ctrl[3].r.part0[21] ,\sa_ctrl[3].r.part0[20] 
	,\sa_ctrl[3].r.part0[19] ,\sa_ctrl[3].r.part0[18] 
	,\sa_ctrl[3].r.part0[17] ,\sa_ctrl[3].r.part0[16] 
	,\sa_ctrl[3].r.part0[15] ,\sa_ctrl[3].r.part0[14] 
	,\sa_ctrl[3].r.part0[13] ,\sa_ctrl[3].r.part0[12] 
	,\sa_ctrl[3].r.part0[11] ,\sa_ctrl[3].r.part0[10] 
	,\sa_ctrl[3].r.part0[9] ,\sa_ctrl[3].r.part0[8] 
	,\sa_ctrl[3].r.part0[7] ,\sa_ctrl[3].r.part0[6] 
	,\sa_ctrl[3].r.part0[5] ,\sa_ctrl[3].r.part0[4] 
	,\sa_ctrl[3].r.part0[3] ,\sa_ctrl[3].r.part0[2] 
	,\sa_ctrl[3].r.part0[1] ,\sa_ctrl[3].r.part0[0] 
	,\sa_ctrl[2].r.part0[31] ,\sa_ctrl[2].r.part0[30] 
	,\sa_ctrl[2].r.part0[29] ,\sa_ctrl[2].r.part0[28] 
	,\sa_ctrl[2].r.part0[27] ,\sa_ctrl[2].r.part0[26] 
	,\sa_ctrl[2].r.part0[25] ,\sa_ctrl[2].r.part0[24] 
	,\sa_ctrl[2].r.part0[23] ,\sa_ctrl[2].r.part0[22] 
	,\sa_ctrl[2].r.part0[21] ,\sa_ctrl[2].r.part0[20] 
	,\sa_ctrl[2].r.part0[19] ,\sa_ctrl[2].r.part0[18] 
	,\sa_ctrl[2].r.part0[17] ,\sa_ctrl[2].r.part0[16] 
	,\sa_ctrl[2].r.part0[15] ,\sa_ctrl[2].r.part0[14] 
	,\sa_ctrl[2].r.part0[13] ,\sa_ctrl[2].r.part0[12] 
	,\sa_ctrl[2].r.part0[11] ,\sa_ctrl[2].r.part0[10] 
	,\sa_ctrl[2].r.part0[9] ,\sa_ctrl[2].r.part0[8] 
	,\sa_ctrl[2].r.part0[7] ,\sa_ctrl[2].r.part0[6] 
	,\sa_ctrl[2].r.part0[5] ,\sa_ctrl[2].r.part0[4] 
	,\sa_ctrl[2].r.part0[3] ,\sa_ctrl[2].r.part0[2] 
	,\sa_ctrl[2].r.part0[1] ,\sa_ctrl[2].r.part0[0] 
	,\sa_ctrl[1].r.part0[31] ,\sa_ctrl[1].r.part0[30] 
	,\sa_ctrl[1].r.part0[29] ,\sa_ctrl[1].r.part0[28] 
	,\sa_ctrl[1].r.part0[27] ,\sa_ctrl[1].r.part0[26] 
	,\sa_ctrl[1].r.part0[25] ,\sa_ctrl[1].r.part0[24] 
	,\sa_ctrl[1].r.part0[23] ,\sa_ctrl[1].r.part0[22] 
	,\sa_ctrl[1].r.part0[21] ,\sa_ctrl[1].r.part0[20] 
	,\sa_ctrl[1].r.part0[19] ,\sa_ctrl[1].r.part0[18] 
	,\sa_ctrl[1].r.part0[17] ,\sa_ctrl[1].r.part0[16] 
	,\sa_ctrl[1].r.part0[15] ,\sa_ctrl[1].r.part0[14] 
	,\sa_ctrl[1].r.part0[13] ,\sa_ctrl[1].r.part0[12] 
	,\sa_ctrl[1].r.part0[11] ,\sa_ctrl[1].r.part0[10] 
	,\sa_ctrl[1].r.part0[9] ,\sa_ctrl[1].r.part0[8] 
	,\sa_ctrl[1].r.part0[7] ,\sa_ctrl[1].r.part0[6] 
	,\sa_ctrl[1].r.part0[5] ,\sa_ctrl[1].r.part0[4] 
	,\sa_ctrl[1].r.part0[3] ,\sa_ctrl[1].r.part0[2] 
	,\sa_ctrl[1].r.part0[1] ,\sa_ctrl[1].r.part0[0] 
	,\sa_ctrl[0].r.part0[31] ,\sa_ctrl[0].r.part0[30] 
	,\sa_ctrl[0].r.part0[29] ,\sa_ctrl[0].r.part0[28] 
	,\sa_ctrl[0].r.part0[27] ,\sa_ctrl[0].r.part0[26] 
	,\sa_ctrl[0].r.part0[25] ,\sa_ctrl[0].r.part0[24] 
	,\sa_ctrl[0].r.part0[23] ,\sa_ctrl[0].r.part0[22] 
	,\sa_ctrl[0].r.part0[21] ,\sa_ctrl[0].r.part0[20] 
	,\sa_ctrl[0].r.part0[19] ,\sa_ctrl[0].r.part0[18] 
	,\sa_ctrl[0].r.part0[17] ,\sa_ctrl[0].r.part0[16] 
	,\sa_ctrl[0].r.part0[15] ,\sa_ctrl[0].r.part0[14] 
	,\sa_ctrl[0].r.part0[13] ,\sa_ctrl[0].r.part0[12] 
	,\sa_ctrl[0].r.part0[11] ,\sa_ctrl[0].r.part0[10] 
	,\sa_ctrl[0].r.part0[9] ,\sa_ctrl[0].r.part0[8] 
	,\sa_ctrl[0].r.part0[7] ,\sa_ctrl[0].r.part0[6] 
	,\sa_ctrl[0].r.part0[5] ,\sa_ctrl[0].r.part0[4] 
	,\sa_ctrl[0].r.part0[3] ,\sa_ctrl[0].r.part0[2] 
	,\sa_ctrl[0].r.part0[1] ,\sa_ctrl[0].r.part0[0] ;
output debug_kme_ib_tvalid;
output debug_kme_ib_tlast;
output [0:0] debug_kme_ib_tid;
output [7:0] debug_kme_ib_tstrb;
output [7:0] debug_kme_ib_tuser;
output [63:0] debug_kme_ib_tdata;
input clk;
input rst_n;
input ovstb;
input lvm;
input mlvm;
input [15:0] \rbus_ring_i.addr ;
input \rbus_ring_i.wr_strb ;
input [31:0] \rbus_ring_i.wr_data ;
input \rbus_ring_i.rd_strb ;
input [31:0] \rbus_ring_i.rd_data ;
input \rbus_ring_i.ack ;
input \rbus_ring_i.err_ack ;
wire [83:0] rbus_ring_i;
input [15:0] cfg_start_addr;
input [15:0] cfg_end_addr;
input \kme_cceip0_ob_out_pre.tvalid ;
input \kme_cceip0_ob_out_pre.tlast ;
input [0:0] \kme_cceip0_ob_out_pre.tid ;
input [7:0] \kme_cceip0_ob_out_pre.tstrb ;
input [7:0] \kme_cceip0_ob_out_pre.tuser ;
input [63:0] \kme_cceip0_ob_out_pre.tdata ;
wire [82:0] kme_cceip0_ob_out_pre;
input \kme_cceip0_ob_in.tready ;
wire [0:0] kme_cceip0_ob_in;
input \kme_cceip1_ob_out_pre.tvalid ;
input \kme_cceip1_ob_out_pre.tlast ;
input [0:0] \kme_cceip1_ob_out_pre.tid ;
input [7:0] \kme_cceip1_ob_out_pre.tstrb ;
input [7:0] \kme_cceip1_ob_out_pre.tuser ;
input [63:0] \kme_cceip1_ob_out_pre.tdata ;
wire [82:0] kme_cceip1_ob_out_pre;
input \kme_cceip1_ob_in.tready ;
wire [0:0] kme_cceip1_ob_in;
input \kme_cceip2_ob_out_pre.tvalid ;
input \kme_cceip2_ob_out_pre.tlast ;
input [0:0] \kme_cceip2_ob_out_pre.tid ;
input [7:0] \kme_cceip2_ob_out_pre.tstrb ;
input [7:0] \kme_cceip2_ob_out_pre.tuser ;
input [63:0] \kme_cceip2_ob_out_pre.tdata ;
wire [82:0] kme_cceip2_ob_out_pre;
input \kme_cceip2_ob_in.tready ;
wire [0:0] kme_cceip2_ob_in;
input \kme_cceip3_ob_out_pre.tvalid ;
input \kme_cceip3_ob_out_pre.tlast ;
input [0:0] \kme_cceip3_ob_out_pre.tid ;
input [7:0] \kme_cceip3_ob_out_pre.tstrb ;
input [7:0] \kme_cceip3_ob_out_pre.tuser ;
input [63:0] \kme_cceip3_ob_out_pre.tdata ;
wire [82:0] kme_cceip3_ob_out_pre;
input \kme_cceip3_ob_in.tready ;
wire [0:0] kme_cceip3_ob_in;
input \kme_cddip0_ob_out_pre.tvalid ;
input \kme_cddip0_ob_out_pre.tlast ;
input [0:0] \kme_cddip0_ob_out_pre.tid ;
input [7:0] \kme_cddip0_ob_out_pre.tstrb ;
input [7:0] \kme_cddip0_ob_out_pre.tuser ;
input [63:0] \kme_cddip0_ob_out_pre.tdata ;
wire [82:0] kme_cddip0_ob_out_pre;
input \kme_cddip0_ob_in.tready ;
wire [0:0] kme_cddip0_ob_in;
input \kme_cddip1_ob_out_pre.tvalid ;
input \kme_cddip1_ob_out_pre.tlast ;
input [0:0] \kme_cddip1_ob_out_pre.tid ;
input [7:0] \kme_cddip1_ob_out_pre.tstrb ;
input [7:0] \kme_cddip1_ob_out_pre.tuser ;
input [63:0] \kme_cddip1_ob_out_pre.tdata ;
wire [82:0] kme_cddip1_ob_out_pre;
input \kme_cddip1_ob_in.tready ;
wire [0:0] kme_cddip1_ob_in;
input \kme_cddip2_ob_out_pre.tvalid ;
input \kme_cddip2_ob_out_pre.tlast ;
input [0:0] \kme_cddip2_ob_out_pre.tid ;
input [7:0] \kme_cddip2_ob_out_pre.tstrb ;
input [7:0] \kme_cddip2_ob_out_pre.tuser ;
input [63:0] \kme_cddip2_ob_out_pre.tdata ;
wire [82:0] kme_cddip2_ob_out_pre;
input \kme_cddip2_ob_in.tready ;
wire [0:0] kme_cddip2_ob_in;
input \kme_cddip3_ob_out_pre.tvalid ;
input \kme_cddip3_ob_out_pre.tlast ;
input [0:0] \kme_cddip3_ob_out_pre.tid ;
input [7:0] \kme_cddip3_ob_out_pre.tstrb ;
input [7:0] \kme_cddip3_ob_out_pre.tuser ;
input [63:0] \kme_cddip3_ob_out_pre.tdata ;
wire [82:0] kme_cddip3_ob_out_pre;
input \kme_cddip3_ob_in.tready ;
wire [0:0] kme_cddip3_ob_in;
input ckv_rd;
input [14:0] ckv_addr;
input kim_rd;
input [13:0] kim_addr;
input cceip_encrypt_bimc_osync;
input cceip_encrypt_bimc_odat;
input cceip_encrypt_mbe;
input cceip_validate_bimc_osync;
input cceip_validate_bimc_odat;
input cceip_validate_mbe;
input cddip_decrypt_bimc_osync;
input cddip_decrypt_bimc_odat;
input cddip_decrypt_mbe;
input axi_bimc_osync;
input axi_bimc_odat;
input axi_mbe;
input seed0_invalidate;
input seed1_invalidate;
input set_txc_bp_int;
input set_gcm_tag_fail_int;
input set_key_tlv_miscmp_int;
input set_tlv_bip2_error_int;
input [7:0] set_rsm_is_backpressuring;
input [31:0] \idle_components.r.part0 ;
wire [19:0] \idle_components.f.num_key_tlvs_in_flight ;
wire \idle_components.f.cddip0_key_tlv_rsm_idle ;
wire \idle_components.f.cddip1_key_tlv_rsm_idle ;
wire \idle_components.f.cddip2_key_tlv_rsm_idle ;
wire \idle_components.f.cddip3_key_tlv_rsm_idle ;
wire \idle_components.f.cceip0_key_tlv_rsm_idle ;
wire \idle_components.f.cceip1_key_tlv_rsm_idle ;
wire \idle_components.f.cceip2_key_tlv_rsm_idle ;
wire \idle_components.f.cceip3_key_tlv_rsm_idle ;
wire \idle_components.f.no_key_tlv_in_flight ;
wire \idle_components.f.tlv_parser_idle ;
wire \idle_components.f.drng_idle ;
wire \idle_components.f.kme_slv_empty ;
wire [31:0] idle_components;
input \sa_snapshot[31].r.part1[31] ,\sa_snapshot[31].r.part1[30] 
	,\sa_snapshot[31].r.part1[29] ,\sa_snapshot[31].r.part1[28] 
	,\sa_snapshot[31].r.part1[27] ,\sa_snapshot[31].r.part1[26] 
	,\sa_snapshot[31].r.part1[25] ,\sa_snapshot[31].r.part1[24] 
	,\sa_snapshot[31].r.part1[23] ,\sa_snapshot[31].r.part1[22] 
	,\sa_snapshot[31].r.part1[21] ,\sa_snapshot[31].r.part1[20] 
	,\sa_snapshot[31].r.part1[19] ,\sa_snapshot[31].r.part1[18] 
	,\sa_snapshot[31].r.part1[17] ,\sa_snapshot[31].r.part1[16] 
	,\sa_snapshot[31].r.part1[15] ,\sa_snapshot[31].r.part1[14] 
	,\sa_snapshot[31].r.part1[13] ,\sa_snapshot[31].r.part1[12] 
	,\sa_snapshot[31].r.part1[11] ,\sa_snapshot[31].r.part1[10] 
	,\sa_snapshot[31].r.part1[9] ,\sa_snapshot[31].r.part1[8] 
	,\sa_snapshot[31].r.part1[7] ,\sa_snapshot[31].r.part1[6] 
	,\sa_snapshot[31].r.part1[5] ,\sa_snapshot[31].r.part1[4] 
	,\sa_snapshot[31].r.part1[3] ,\sa_snapshot[31].r.part1[2] 
	,\sa_snapshot[31].r.part1[1] ,\sa_snapshot[31].r.part1[0] 
	,\sa_snapshot[31].r.part0[31] ,\sa_snapshot[31].r.part0[30] 
	,\sa_snapshot[31].r.part0[29] ,\sa_snapshot[31].r.part0[28] 
	,\sa_snapshot[31].r.part0[27] ,\sa_snapshot[31].r.part0[26] 
	,\sa_snapshot[31].r.part0[25] ,\sa_snapshot[31].r.part0[24] 
	,\sa_snapshot[31].r.part0[23] ,\sa_snapshot[31].r.part0[22] 
	,\sa_snapshot[31].r.part0[21] ,\sa_snapshot[31].r.part0[20] 
	,\sa_snapshot[31].r.part0[19] ,\sa_snapshot[31].r.part0[18] 
	,\sa_snapshot[31].r.part0[17] ,\sa_snapshot[31].r.part0[16] 
	,\sa_snapshot[31].r.part0[15] ,\sa_snapshot[31].r.part0[14] 
	,\sa_snapshot[31].r.part0[13] ,\sa_snapshot[31].r.part0[12] 
	,\sa_snapshot[31].r.part0[11] ,\sa_snapshot[31].r.part0[10] 
	,\sa_snapshot[31].r.part0[9] ,\sa_snapshot[31].r.part0[8] 
	,\sa_snapshot[31].r.part0[7] ,\sa_snapshot[31].r.part0[6] 
	,\sa_snapshot[31].r.part0[5] ,\sa_snapshot[31].r.part0[4] 
	,\sa_snapshot[31].r.part0[3] ,\sa_snapshot[31].r.part0[2] 
	,\sa_snapshot[31].r.part0[1] ,\sa_snapshot[31].r.part0[0] 
	,\sa_snapshot[30].r.part1[31] ,\sa_snapshot[30].r.part1[30] 
	,\sa_snapshot[30].r.part1[29] ,\sa_snapshot[30].r.part1[28] 
	,\sa_snapshot[30].r.part1[27] ,\sa_snapshot[30].r.part1[26] 
	,\sa_snapshot[30].r.part1[25] ,\sa_snapshot[30].r.part1[24] 
	,\sa_snapshot[30].r.part1[23] ,\sa_snapshot[30].r.part1[22] 
	,\sa_snapshot[30].r.part1[21] ,\sa_snapshot[30].r.part1[20] 
	,\sa_snapshot[30].r.part1[19] ,\sa_snapshot[30].r.part1[18] 
	,\sa_snapshot[30].r.part1[17] ,\sa_snapshot[30].r.part1[16] 
	,\sa_snapshot[30].r.part1[15] ,\sa_snapshot[30].r.part1[14] 
	,\sa_snapshot[30].r.part1[13] ,\sa_snapshot[30].r.part1[12] 
	,\sa_snapshot[30].r.part1[11] ,\sa_snapshot[30].r.part1[10] 
	,\sa_snapshot[30].r.part1[9] ,\sa_snapshot[30].r.part1[8] 
	,\sa_snapshot[30].r.part1[7] ,\sa_snapshot[30].r.part1[6] 
	,\sa_snapshot[30].r.part1[5] ,\sa_snapshot[30].r.part1[4] 
	,\sa_snapshot[30].r.part1[3] ,\sa_snapshot[30].r.part1[2] 
	,\sa_snapshot[30].r.part1[1] ,\sa_snapshot[30].r.part1[0] 
	,\sa_snapshot[30].r.part0[31] ,\sa_snapshot[30].r.part0[30] 
	,\sa_snapshot[30].r.part0[29] ,\sa_snapshot[30].r.part0[28] 
	,\sa_snapshot[30].r.part0[27] ,\sa_snapshot[30].r.part0[26] 
	,\sa_snapshot[30].r.part0[25] ,\sa_snapshot[30].r.part0[24] 
	,\sa_snapshot[30].r.part0[23] ,\sa_snapshot[30].r.part0[22] 
	,\sa_snapshot[30].r.part0[21] ,\sa_snapshot[30].r.part0[20] 
	,\sa_snapshot[30].r.part0[19] ,\sa_snapshot[30].r.part0[18] 
	,\sa_snapshot[30].r.part0[17] ,\sa_snapshot[30].r.part0[16] 
	,\sa_snapshot[30].r.part0[15] ,\sa_snapshot[30].r.part0[14] 
	,\sa_snapshot[30].r.part0[13] ,\sa_snapshot[30].r.part0[12] 
	,\sa_snapshot[30].r.part0[11] ,\sa_snapshot[30].r.part0[10] 
	,\sa_snapshot[30].r.part0[9] ,\sa_snapshot[30].r.part0[8] 
	,\sa_snapshot[30].r.part0[7] ,\sa_snapshot[30].r.part0[6] 
	,\sa_snapshot[30].r.part0[5] ,\sa_snapshot[30].r.part0[4] 
	,\sa_snapshot[30].r.part0[3] ,\sa_snapshot[30].r.part0[2] 
	,\sa_snapshot[30].r.part0[1] ,\sa_snapshot[30].r.part0[0] 
	,\sa_snapshot[29].r.part1[31] ,\sa_snapshot[29].r.part1[30] 
	,\sa_snapshot[29].r.part1[29] ,\sa_snapshot[29].r.part1[28] 
	,\sa_snapshot[29].r.part1[27] ,\sa_snapshot[29].r.part1[26] 
	,\sa_snapshot[29].r.part1[25] ,\sa_snapshot[29].r.part1[24] 
	,\sa_snapshot[29].r.part1[23] ,\sa_snapshot[29].r.part1[22] 
	,\sa_snapshot[29].r.part1[21] ,\sa_snapshot[29].r.part1[20] 
	,\sa_snapshot[29].r.part1[19] ,\sa_snapshot[29].r.part1[18] 
	,\sa_snapshot[29].r.part1[17] ,\sa_snapshot[29].r.part1[16] 
	,\sa_snapshot[29].r.part1[15] ,\sa_snapshot[29].r.part1[14] 
	,\sa_snapshot[29].r.part1[13] ,\sa_snapshot[29].r.part1[12] 
	,\sa_snapshot[29].r.part1[11] ,\sa_snapshot[29].r.part1[10] 
	,\sa_snapshot[29].r.part1[9] ,\sa_snapshot[29].r.part1[8] 
	,\sa_snapshot[29].r.part1[7] ,\sa_snapshot[29].r.part1[6] 
	,\sa_snapshot[29].r.part1[5] ,\sa_snapshot[29].r.part1[4] 
	,\sa_snapshot[29].r.part1[3] ,\sa_snapshot[29].r.part1[2] 
	,\sa_snapshot[29].r.part1[1] ,\sa_snapshot[29].r.part1[0] 
	,\sa_snapshot[29].r.part0[31] ,\sa_snapshot[29].r.part0[30] 
	,\sa_snapshot[29].r.part0[29] ,\sa_snapshot[29].r.part0[28] 
	,\sa_snapshot[29].r.part0[27] ,\sa_snapshot[29].r.part0[26] 
	,\sa_snapshot[29].r.part0[25] ,\sa_snapshot[29].r.part0[24] 
	,\sa_snapshot[29].r.part0[23] ,\sa_snapshot[29].r.part0[22] 
	,\sa_snapshot[29].r.part0[21] ,\sa_snapshot[29].r.part0[20] 
	,\sa_snapshot[29].r.part0[19] ,\sa_snapshot[29].r.part0[18] 
	,\sa_snapshot[29].r.part0[17] ,\sa_snapshot[29].r.part0[16] 
	,\sa_snapshot[29].r.part0[15] ,\sa_snapshot[29].r.part0[14] 
	,\sa_snapshot[29].r.part0[13] ,\sa_snapshot[29].r.part0[12] 
	,\sa_snapshot[29].r.part0[11] ,\sa_snapshot[29].r.part0[10] 
	,\sa_snapshot[29].r.part0[9] ,\sa_snapshot[29].r.part0[8] 
	,\sa_snapshot[29].r.part0[7] ,\sa_snapshot[29].r.part0[6] 
	,\sa_snapshot[29].r.part0[5] ,\sa_snapshot[29].r.part0[4] 
	,\sa_snapshot[29].r.part0[3] ,\sa_snapshot[29].r.part0[2] 
	,\sa_snapshot[29].r.part0[1] ,\sa_snapshot[29].r.part0[0] 
	,\sa_snapshot[28].r.part1[31] ,\sa_snapshot[28].r.part1[30] 
	,\sa_snapshot[28].r.part1[29] ,\sa_snapshot[28].r.part1[28] 
	,\sa_snapshot[28].r.part1[27] ,\sa_snapshot[28].r.part1[26] 
	,\sa_snapshot[28].r.part1[25] ,\sa_snapshot[28].r.part1[24] 
	,\sa_snapshot[28].r.part1[23] ,\sa_snapshot[28].r.part1[22] 
	,\sa_snapshot[28].r.part1[21] ,\sa_snapshot[28].r.part1[20] 
	,\sa_snapshot[28].r.part1[19] ,\sa_snapshot[28].r.part1[18] 
	,\sa_snapshot[28].r.part1[17] ,\sa_snapshot[28].r.part1[16] 
	,\sa_snapshot[28].r.part1[15] ,\sa_snapshot[28].r.part1[14] 
	,\sa_snapshot[28].r.part1[13] ,\sa_snapshot[28].r.part1[12] 
	,\sa_snapshot[28].r.part1[11] ,\sa_snapshot[28].r.part1[10] 
	,\sa_snapshot[28].r.part1[9] ,\sa_snapshot[28].r.part1[8] 
	,\sa_snapshot[28].r.part1[7] ,\sa_snapshot[28].r.part1[6] 
	,\sa_snapshot[28].r.part1[5] ,\sa_snapshot[28].r.part1[4] 
	,\sa_snapshot[28].r.part1[3] ,\sa_snapshot[28].r.part1[2] 
	,\sa_snapshot[28].r.part1[1] ,\sa_snapshot[28].r.part1[0] 
	,\sa_snapshot[28].r.part0[31] ,\sa_snapshot[28].r.part0[30] 
	,\sa_snapshot[28].r.part0[29] ,\sa_snapshot[28].r.part0[28] 
	,\sa_snapshot[28].r.part0[27] ,\sa_snapshot[28].r.part0[26] 
	,\sa_snapshot[28].r.part0[25] ,\sa_snapshot[28].r.part0[24] 
	,\sa_snapshot[28].r.part0[23] ,\sa_snapshot[28].r.part0[22] 
	,\sa_snapshot[28].r.part0[21] ,\sa_snapshot[28].r.part0[20] 
	,\sa_snapshot[28].r.part0[19] ,\sa_snapshot[28].r.part0[18] 
	,\sa_snapshot[28].r.part0[17] ,\sa_snapshot[28].r.part0[16] 
	,\sa_snapshot[28].r.part0[15] ,\sa_snapshot[28].r.part0[14] 
	,\sa_snapshot[28].r.part0[13] ,\sa_snapshot[28].r.part0[12] 
	,\sa_snapshot[28].r.part0[11] ,\sa_snapshot[28].r.part0[10] 
	,\sa_snapshot[28].r.part0[9] ,\sa_snapshot[28].r.part0[8] 
	,\sa_snapshot[28].r.part0[7] ,\sa_snapshot[28].r.part0[6] 
	,\sa_snapshot[28].r.part0[5] ,\sa_snapshot[28].r.part0[4] 
	,\sa_snapshot[28].r.part0[3] ,\sa_snapshot[28].r.part0[2] 
	,\sa_snapshot[28].r.part0[1] ,\sa_snapshot[28].r.part0[0] 
	,\sa_snapshot[27].r.part1[31] ,\sa_snapshot[27].r.part1[30] 
	,\sa_snapshot[27].r.part1[29] ,\sa_snapshot[27].r.part1[28] 
	,\sa_snapshot[27].r.part1[27] ,\sa_snapshot[27].r.part1[26] 
	,\sa_snapshot[27].r.part1[25] ,\sa_snapshot[27].r.part1[24] 
	,\sa_snapshot[27].r.part1[23] ,\sa_snapshot[27].r.part1[22] 
	,\sa_snapshot[27].r.part1[21] ,\sa_snapshot[27].r.part1[20] 
	,\sa_snapshot[27].r.part1[19] ,\sa_snapshot[27].r.part1[18] 
	,\sa_snapshot[27].r.part1[17] ,\sa_snapshot[27].r.part1[16] 
	,\sa_snapshot[27].r.part1[15] ,\sa_snapshot[27].r.part1[14] 
	,\sa_snapshot[27].r.part1[13] ,\sa_snapshot[27].r.part1[12] 
	,\sa_snapshot[27].r.part1[11] ,\sa_snapshot[27].r.part1[10] 
	,\sa_snapshot[27].r.part1[9] ,\sa_snapshot[27].r.part1[8] 
	,\sa_snapshot[27].r.part1[7] ,\sa_snapshot[27].r.part1[6] 
	,\sa_snapshot[27].r.part1[5] ,\sa_snapshot[27].r.part1[4] 
	,\sa_snapshot[27].r.part1[3] ,\sa_snapshot[27].r.part1[2] 
	,\sa_snapshot[27].r.part1[1] ,\sa_snapshot[27].r.part1[0] 
	,\sa_snapshot[27].r.part0[31] ,\sa_snapshot[27].r.part0[30] 
	,\sa_snapshot[27].r.part0[29] ,\sa_snapshot[27].r.part0[28] 
	,\sa_snapshot[27].r.part0[27] ,\sa_snapshot[27].r.part0[26] 
	,\sa_snapshot[27].r.part0[25] ,\sa_snapshot[27].r.part0[24] 
	,\sa_snapshot[27].r.part0[23] ,\sa_snapshot[27].r.part0[22] 
	,\sa_snapshot[27].r.part0[21] ,\sa_snapshot[27].r.part0[20] 
	,\sa_snapshot[27].r.part0[19] ,\sa_snapshot[27].r.part0[18] 
	,\sa_snapshot[27].r.part0[17] ,\sa_snapshot[27].r.part0[16] 
	,\sa_snapshot[27].r.part0[15] ,\sa_snapshot[27].r.part0[14] 
	,\sa_snapshot[27].r.part0[13] ,\sa_snapshot[27].r.part0[12] 
	,\sa_snapshot[27].r.part0[11] ,\sa_snapshot[27].r.part0[10] 
	,\sa_snapshot[27].r.part0[9] ,\sa_snapshot[27].r.part0[8] 
	,\sa_snapshot[27].r.part0[7] ,\sa_snapshot[27].r.part0[6] 
	,\sa_snapshot[27].r.part0[5] ,\sa_snapshot[27].r.part0[4] 
	,\sa_snapshot[27].r.part0[3] ,\sa_snapshot[27].r.part0[2] 
	,\sa_snapshot[27].r.part0[1] ,\sa_snapshot[27].r.part0[0] 
	,\sa_snapshot[26].r.part1[31] ,\sa_snapshot[26].r.part1[30] 
	,\sa_snapshot[26].r.part1[29] ,\sa_snapshot[26].r.part1[28] 
	,\sa_snapshot[26].r.part1[27] ,\sa_snapshot[26].r.part1[26] 
	,\sa_snapshot[26].r.part1[25] ,\sa_snapshot[26].r.part1[24] 
	,\sa_snapshot[26].r.part1[23] ,\sa_snapshot[26].r.part1[22] 
	,\sa_snapshot[26].r.part1[21] ,\sa_snapshot[26].r.part1[20] 
	,\sa_snapshot[26].r.part1[19] ,\sa_snapshot[26].r.part1[18] 
	,\sa_snapshot[26].r.part1[17] ,\sa_snapshot[26].r.part1[16] 
	,\sa_snapshot[26].r.part1[15] ,\sa_snapshot[26].r.part1[14] 
	,\sa_snapshot[26].r.part1[13] ,\sa_snapshot[26].r.part1[12] 
	,\sa_snapshot[26].r.part1[11] ,\sa_snapshot[26].r.part1[10] 
	,\sa_snapshot[26].r.part1[9] ,\sa_snapshot[26].r.part1[8] 
	,\sa_snapshot[26].r.part1[7] ,\sa_snapshot[26].r.part1[6] 
	,\sa_snapshot[26].r.part1[5] ,\sa_snapshot[26].r.part1[4] 
	,\sa_snapshot[26].r.part1[3] ,\sa_snapshot[26].r.part1[2] 
	,\sa_snapshot[26].r.part1[1] ,\sa_snapshot[26].r.part1[0] 
	,\sa_snapshot[26].r.part0[31] ,\sa_snapshot[26].r.part0[30] 
	,\sa_snapshot[26].r.part0[29] ,\sa_snapshot[26].r.part0[28] 
	,\sa_snapshot[26].r.part0[27] ,\sa_snapshot[26].r.part0[26] 
	,\sa_snapshot[26].r.part0[25] ,\sa_snapshot[26].r.part0[24] 
	,\sa_snapshot[26].r.part0[23] ,\sa_snapshot[26].r.part0[22] 
	,\sa_snapshot[26].r.part0[21] ,\sa_snapshot[26].r.part0[20] 
	,\sa_snapshot[26].r.part0[19] ,\sa_snapshot[26].r.part0[18] 
	,\sa_snapshot[26].r.part0[17] ,\sa_snapshot[26].r.part0[16] 
	,\sa_snapshot[26].r.part0[15] ,\sa_snapshot[26].r.part0[14] 
	,\sa_snapshot[26].r.part0[13] ,\sa_snapshot[26].r.part0[12] 
	,\sa_snapshot[26].r.part0[11] ,\sa_snapshot[26].r.part0[10] 
	,\sa_snapshot[26].r.part0[9] ,\sa_snapshot[26].r.part0[8] 
	,\sa_snapshot[26].r.part0[7] ,\sa_snapshot[26].r.part0[6] 
	,\sa_snapshot[26].r.part0[5] ,\sa_snapshot[26].r.part0[4] 
	,\sa_snapshot[26].r.part0[3] ,\sa_snapshot[26].r.part0[2] 
	,\sa_snapshot[26].r.part0[1] ,\sa_snapshot[26].r.part0[0] 
	,\sa_snapshot[25].r.part1[31] ,\sa_snapshot[25].r.part1[30] 
	,\sa_snapshot[25].r.part1[29] ,\sa_snapshot[25].r.part1[28] 
	,\sa_snapshot[25].r.part1[27] ,\sa_snapshot[25].r.part1[26] 
	,\sa_snapshot[25].r.part1[25] ,\sa_snapshot[25].r.part1[24] 
	,\sa_snapshot[25].r.part1[23] ,\sa_snapshot[25].r.part1[22] 
	,\sa_snapshot[25].r.part1[21] ,\sa_snapshot[25].r.part1[20] 
	,\sa_snapshot[25].r.part1[19] ,\sa_snapshot[25].r.part1[18] 
	,\sa_snapshot[25].r.part1[17] ,\sa_snapshot[25].r.part1[16] 
	,\sa_snapshot[25].r.part1[15] ,\sa_snapshot[25].r.part1[14] 
	,\sa_snapshot[25].r.part1[13] ,\sa_snapshot[25].r.part1[12] 
	,\sa_snapshot[25].r.part1[11] ,\sa_snapshot[25].r.part1[10] 
	,\sa_snapshot[25].r.part1[9] ,\sa_snapshot[25].r.part1[8] 
	,\sa_snapshot[25].r.part1[7] ,\sa_snapshot[25].r.part1[6] 
	,\sa_snapshot[25].r.part1[5] ,\sa_snapshot[25].r.part1[4] 
	,\sa_snapshot[25].r.part1[3] ,\sa_snapshot[25].r.part1[2] 
	,\sa_snapshot[25].r.part1[1] ,\sa_snapshot[25].r.part1[0] 
	,\sa_snapshot[25].r.part0[31] ,\sa_snapshot[25].r.part0[30] 
	,\sa_snapshot[25].r.part0[29] ,\sa_snapshot[25].r.part0[28] 
	,\sa_snapshot[25].r.part0[27] ,\sa_snapshot[25].r.part0[26] 
	,\sa_snapshot[25].r.part0[25] ,\sa_snapshot[25].r.part0[24] 
	,\sa_snapshot[25].r.part0[23] ,\sa_snapshot[25].r.part0[22] 
	,\sa_snapshot[25].r.part0[21] ,\sa_snapshot[25].r.part0[20] 
	,\sa_snapshot[25].r.part0[19] ,\sa_snapshot[25].r.part0[18] 
	,\sa_snapshot[25].r.part0[17] ,\sa_snapshot[25].r.part0[16] 
	,\sa_snapshot[25].r.part0[15] ,\sa_snapshot[25].r.part0[14] 
	,\sa_snapshot[25].r.part0[13] ,\sa_snapshot[25].r.part0[12] 
	,\sa_snapshot[25].r.part0[11] ,\sa_snapshot[25].r.part0[10] 
	,\sa_snapshot[25].r.part0[9] ,\sa_snapshot[25].r.part0[8] 
	,\sa_snapshot[25].r.part0[7] ,\sa_snapshot[25].r.part0[6] 
	,\sa_snapshot[25].r.part0[5] ,\sa_snapshot[25].r.part0[4] 
	,\sa_snapshot[25].r.part0[3] ,\sa_snapshot[25].r.part0[2] 
	,\sa_snapshot[25].r.part0[1] ,\sa_snapshot[25].r.part0[0] 
	,\sa_snapshot[24].r.part1[31] ,\sa_snapshot[24].r.part1[30] 
	,\sa_snapshot[24].r.part1[29] ,\sa_snapshot[24].r.part1[28] 
	,\sa_snapshot[24].r.part1[27] ,\sa_snapshot[24].r.part1[26] 
	,\sa_snapshot[24].r.part1[25] ,\sa_snapshot[24].r.part1[24] 
	,\sa_snapshot[24].r.part1[23] ,\sa_snapshot[24].r.part1[22] 
	,\sa_snapshot[24].r.part1[21] ,\sa_snapshot[24].r.part1[20] 
	,\sa_snapshot[24].r.part1[19] ,\sa_snapshot[24].r.part1[18] 
	,\sa_snapshot[24].r.part1[17] ,\sa_snapshot[24].r.part1[16] 
	,\sa_snapshot[24].r.part1[15] ,\sa_snapshot[24].r.part1[14] 
	,\sa_snapshot[24].r.part1[13] ,\sa_snapshot[24].r.part1[12] 
	,\sa_snapshot[24].r.part1[11] ,\sa_snapshot[24].r.part1[10] 
	,\sa_snapshot[24].r.part1[9] ,\sa_snapshot[24].r.part1[8] 
	,\sa_snapshot[24].r.part1[7] ,\sa_snapshot[24].r.part1[6] 
	,\sa_snapshot[24].r.part1[5] ,\sa_snapshot[24].r.part1[4] 
	,\sa_snapshot[24].r.part1[3] ,\sa_snapshot[24].r.part1[2] 
	,\sa_snapshot[24].r.part1[1] ,\sa_snapshot[24].r.part1[0] 
	,\sa_snapshot[24].r.part0[31] ,\sa_snapshot[24].r.part0[30] 
	,\sa_snapshot[24].r.part0[29] ,\sa_snapshot[24].r.part0[28] 
	,\sa_snapshot[24].r.part0[27] ,\sa_snapshot[24].r.part0[26] 
	,\sa_snapshot[24].r.part0[25] ,\sa_snapshot[24].r.part0[24] 
	,\sa_snapshot[24].r.part0[23] ,\sa_snapshot[24].r.part0[22] 
	,\sa_snapshot[24].r.part0[21] ,\sa_snapshot[24].r.part0[20] 
	,\sa_snapshot[24].r.part0[19] ,\sa_snapshot[24].r.part0[18] 
	,\sa_snapshot[24].r.part0[17] ,\sa_snapshot[24].r.part0[16] 
	,\sa_snapshot[24].r.part0[15] ,\sa_snapshot[24].r.part0[14] 
	,\sa_snapshot[24].r.part0[13] ,\sa_snapshot[24].r.part0[12] 
	,\sa_snapshot[24].r.part0[11] ,\sa_snapshot[24].r.part0[10] 
	,\sa_snapshot[24].r.part0[9] ,\sa_snapshot[24].r.part0[8] 
	,\sa_snapshot[24].r.part0[7] ,\sa_snapshot[24].r.part0[6] 
	,\sa_snapshot[24].r.part0[5] ,\sa_snapshot[24].r.part0[4] 
	,\sa_snapshot[24].r.part0[3] ,\sa_snapshot[24].r.part0[2] 
	,\sa_snapshot[24].r.part0[1] ,\sa_snapshot[24].r.part0[0] 
	,\sa_snapshot[23].r.part1[31] ,\sa_snapshot[23].r.part1[30] 
	,\sa_snapshot[23].r.part1[29] ,\sa_snapshot[23].r.part1[28] 
	,\sa_snapshot[23].r.part1[27] ,\sa_snapshot[23].r.part1[26] 
	,\sa_snapshot[23].r.part1[25] ,\sa_snapshot[23].r.part1[24] 
	,\sa_snapshot[23].r.part1[23] ,\sa_snapshot[23].r.part1[22] 
	,\sa_snapshot[23].r.part1[21] ,\sa_snapshot[23].r.part1[20] 
	,\sa_snapshot[23].r.part1[19] ,\sa_snapshot[23].r.part1[18] 
	,\sa_snapshot[23].r.part1[17] ,\sa_snapshot[23].r.part1[16] 
	,\sa_snapshot[23].r.part1[15] ,\sa_snapshot[23].r.part1[14] 
	,\sa_snapshot[23].r.part1[13] ,\sa_snapshot[23].r.part1[12] 
	,\sa_snapshot[23].r.part1[11] ,\sa_snapshot[23].r.part1[10] 
	,\sa_snapshot[23].r.part1[9] ,\sa_snapshot[23].r.part1[8] 
	,\sa_snapshot[23].r.part1[7] ,\sa_snapshot[23].r.part1[6] 
	,\sa_snapshot[23].r.part1[5] ,\sa_snapshot[23].r.part1[4] 
	,\sa_snapshot[23].r.part1[3] ,\sa_snapshot[23].r.part1[2] 
	,\sa_snapshot[23].r.part1[1] ,\sa_snapshot[23].r.part1[0] 
	,\sa_snapshot[23].r.part0[31] ,\sa_snapshot[23].r.part0[30] 
	,\sa_snapshot[23].r.part0[29] ,\sa_snapshot[23].r.part0[28] 
	,\sa_snapshot[23].r.part0[27] ,\sa_snapshot[23].r.part0[26] 
	,\sa_snapshot[23].r.part0[25] ,\sa_snapshot[23].r.part0[24] 
	,\sa_snapshot[23].r.part0[23] ,\sa_snapshot[23].r.part0[22] 
	,\sa_snapshot[23].r.part0[21] ,\sa_snapshot[23].r.part0[20] 
	,\sa_snapshot[23].r.part0[19] ,\sa_snapshot[23].r.part0[18] 
	,\sa_snapshot[23].r.part0[17] ,\sa_snapshot[23].r.part0[16] 
	,\sa_snapshot[23].r.part0[15] ,\sa_snapshot[23].r.part0[14] 
	,\sa_snapshot[23].r.part0[13] ,\sa_snapshot[23].r.part0[12] 
	,\sa_snapshot[23].r.part0[11] ,\sa_snapshot[23].r.part0[10] 
	,\sa_snapshot[23].r.part0[9] ,\sa_snapshot[23].r.part0[8] 
	,\sa_snapshot[23].r.part0[7] ,\sa_snapshot[23].r.part0[6] 
	,\sa_snapshot[23].r.part0[5] ,\sa_snapshot[23].r.part0[4] 
	,\sa_snapshot[23].r.part0[3] ,\sa_snapshot[23].r.part0[2] 
	,\sa_snapshot[23].r.part0[1] ,\sa_snapshot[23].r.part0[0] 
	,\sa_snapshot[22].r.part1[31] ,\sa_snapshot[22].r.part1[30] 
	,\sa_snapshot[22].r.part1[29] ,\sa_snapshot[22].r.part1[28] 
	,\sa_snapshot[22].r.part1[27] ,\sa_snapshot[22].r.part1[26] 
	,\sa_snapshot[22].r.part1[25] ,\sa_snapshot[22].r.part1[24] 
	,\sa_snapshot[22].r.part1[23] ,\sa_snapshot[22].r.part1[22] 
	,\sa_snapshot[22].r.part1[21] ,\sa_snapshot[22].r.part1[20] 
	,\sa_snapshot[22].r.part1[19] ,\sa_snapshot[22].r.part1[18] 
	,\sa_snapshot[22].r.part1[17] ,\sa_snapshot[22].r.part1[16] 
	,\sa_snapshot[22].r.part1[15] ,\sa_snapshot[22].r.part1[14] 
	,\sa_snapshot[22].r.part1[13] ,\sa_snapshot[22].r.part1[12] 
	,\sa_snapshot[22].r.part1[11] ,\sa_snapshot[22].r.part1[10] 
	,\sa_snapshot[22].r.part1[9] ,\sa_snapshot[22].r.part1[8] 
	,\sa_snapshot[22].r.part1[7] ,\sa_snapshot[22].r.part1[6] 
	,\sa_snapshot[22].r.part1[5] ,\sa_snapshot[22].r.part1[4] 
	,\sa_snapshot[22].r.part1[3] ,\sa_snapshot[22].r.part1[2] 
	,\sa_snapshot[22].r.part1[1] ,\sa_snapshot[22].r.part1[0] 
	,\sa_snapshot[22].r.part0[31] ,\sa_snapshot[22].r.part0[30] 
	,\sa_snapshot[22].r.part0[29] ,\sa_snapshot[22].r.part0[28] 
	,\sa_snapshot[22].r.part0[27] ,\sa_snapshot[22].r.part0[26] 
	,\sa_snapshot[22].r.part0[25] ,\sa_snapshot[22].r.part0[24] 
	,\sa_snapshot[22].r.part0[23] ,\sa_snapshot[22].r.part0[22] 
	,\sa_snapshot[22].r.part0[21] ,\sa_snapshot[22].r.part0[20] 
	,\sa_snapshot[22].r.part0[19] ,\sa_snapshot[22].r.part0[18] 
	,\sa_snapshot[22].r.part0[17] ,\sa_snapshot[22].r.part0[16] 
	,\sa_snapshot[22].r.part0[15] ,\sa_snapshot[22].r.part0[14] 
	,\sa_snapshot[22].r.part0[13] ,\sa_snapshot[22].r.part0[12] 
	,\sa_snapshot[22].r.part0[11] ,\sa_snapshot[22].r.part0[10] 
	,\sa_snapshot[22].r.part0[9] ,\sa_snapshot[22].r.part0[8] 
	,\sa_snapshot[22].r.part0[7] ,\sa_snapshot[22].r.part0[6] 
	,\sa_snapshot[22].r.part0[5] ,\sa_snapshot[22].r.part0[4] 
	,\sa_snapshot[22].r.part0[3] ,\sa_snapshot[22].r.part0[2] 
	,\sa_snapshot[22].r.part0[1] ,\sa_snapshot[22].r.part0[0] 
	,\sa_snapshot[21].r.part1[31] ,\sa_snapshot[21].r.part1[30] 
	,\sa_snapshot[21].r.part1[29] ,\sa_snapshot[21].r.part1[28] 
	,\sa_snapshot[21].r.part1[27] ,\sa_snapshot[21].r.part1[26] 
	,\sa_snapshot[21].r.part1[25] ,\sa_snapshot[21].r.part1[24] 
	,\sa_snapshot[21].r.part1[23] ,\sa_snapshot[21].r.part1[22] 
	,\sa_snapshot[21].r.part1[21] ,\sa_snapshot[21].r.part1[20] 
	,\sa_snapshot[21].r.part1[19] ,\sa_snapshot[21].r.part1[18] 
	,\sa_snapshot[21].r.part1[17] ,\sa_snapshot[21].r.part1[16] 
	,\sa_snapshot[21].r.part1[15] ,\sa_snapshot[21].r.part1[14] 
	,\sa_snapshot[21].r.part1[13] ,\sa_snapshot[21].r.part1[12] 
	,\sa_snapshot[21].r.part1[11] ,\sa_snapshot[21].r.part1[10] 
	,\sa_snapshot[21].r.part1[9] ,\sa_snapshot[21].r.part1[8] 
	,\sa_snapshot[21].r.part1[7] ,\sa_snapshot[21].r.part1[6] 
	,\sa_snapshot[21].r.part1[5] ,\sa_snapshot[21].r.part1[4] 
	,\sa_snapshot[21].r.part1[3] ,\sa_snapshot[21].r.part1[2] 
	,\sa_snapshot[21].r.part1[1] ,\sa_snapshot[21].r.part1[0] 
	,\sa_snapshot[21].r.part0[31] ,\sa_snapshot[21].r.part0[30] 
	,\sa_snapshot[21].r.part0[29] ,\sa_snapshot[21].r.part0[28] 
	,\sa_snapshot[21].r.part0[27] ,\sa_snapshot[21].r.part0[26] 
	,\sa_snapshot[21].r.part0[25] ,\sa_snapshot[21].r.part0[24] 
	,\sa_snapshot[21].r.part0[23] ,\sa_snapshot[21].r.part0[22] 
	,\sa_snapshot[21].r.part0[21] ,\sa_snapshot[21].r.part0[20] 
	,\sa_snapshot[21].r.part0[19] ,\sa_snapshot[21].r.part0[18] 
	,\sa_snapshot[21].r.part0[17] ,\sa_snapshot[21].r.part0[16] 
	,\sa_snapshot[21].r.part0[15] ,\sa_snapshot[21].r.part0[14] 
	,\sa_snapshot[21].r.part0[13] ,\sa_snapshot[21].r.part0[12] 
	,\sa_snapshot[21].r.part0[11] ,\sa_snapshot[21].r.part0[10] 
	,\sa_snapshot[21].r.part0[9] ,\sa_snapshot[21].r.part0[8] 
	,\sa_snapshot[21].r.part0[7] ,\sa_snapshot[21].r.part0[6] 
	,\sa_snapshot[21].r.part0[5] ,\sa_snapshot[21].r.part0[4] 
	,\sa_snapshot[21].r.part0[3] ,\sa_snapshot[21].r.part0[2] 
	,\sa_snapshot[21].r.part0[1] ,\sa_snapshot[21].r.part0[0] 
	,\sa_snapshot[20].r.part1[31] ,\sa_snapshot[20].r.part1[30] 
	,\sa_snapshot[20].r.part1[29] ,\sa_snapshot[20].r.part1[28] 
	,\sa_snapshot[20].r.part1[27] ,\sa_snapshot[20].r.part1[26] 
	,\sa_snapshot[20].r.part1[25] ,\sa_snapshot[20].r.part1[24] 
	,\sa_snapshot[20].r.part1[23] ,\sa_snapshot[20].r.part1[22] 
	,\sa_snapshot[20].r.part1[21] ,\sa_snapshot[20].r.part1[20] 
	,\sa_snapshot[20].r.part1[19] ,\sa_snapshot[20].r.part1[18] 
	,\sa_snapshot[20].r.part1[17] ,\sa_snapshot[20].r.part1[16] 
	,\sa_snapshot[20].r.part1[15] ,\sa_snapshot[20].r.part1[14] 
	,\sa_snapshot[20].r.part1[13] ,\sa_snapshot[20].r.part1[12] 
	,\sa_snapshot[20].r.part1[11] ,\sa_snapshot[20].r.part1[10] 
	,\sa_snapshot[20].r.part1[9] ,\sa_snapshot[20].r.part1[8] 
	,\sa_snapshot[20].r.part1[7] ,\sa_snapshot[20].r.part1[6] 
	,\sa_snapshot[20].r.part1[5] ,\sa_snapshot[20].r.part1[4] 
	,\sa_snapshot[20].r.part1[3] ,\sa_snapshot[20].r.part1[2] 
	,\sa_snapshot[20].r.part1[1] ,\sa_snapshot[20].r.part1[0] 
	,\sa_snapshot[20].r.part0[31] ,\sa_snapshot[20].r.part0[30] 
	,\sa_snapshot[20].r.part0[29] ,\sa_snapshot[20].r.part0[28] 
	,\sa_snapshot[20].r.part0[27] ,\sa_snapshot[20].r.part0[26] 
	,\sa_snapshot[20].r.part0[25] ,\sa_snapshot[20].r.part0[24] 
	,\sa_snapshot[20].r.part0[23] ,\sa_snapshot[20].r.part0[22] 
	,\sa_snapshot[20].r.part0[21] ,\sa_snapshot[20].r.part0[20] 
	,\sa_snapshot[20].r.part0[19] ,\sa_snapshot[20].r.part0[18] 
	,\sa_snapshot[20].r.part0[17] ,\sa_snapshot[20].r.part0[16] 
	,\sa_snapshot[20].r.part0[15] ,\sa_snapshot[20].r.part0[14] 
	,\sa_snapshot[20].r.part0[13] ,\sa_snapshot[20].r.part0[12] 
	,\sa_snapshot[20].r.part0[11] ,\sa_snapshot[20].r.part0[10] 
	,\sa_snapshot[20].r.part0[9] ,\sa_snapshot[20].r.part0[8] 
	,\sa_snapshot[20].r.part0[7] ,\sa_snapshot[20].r.part0[6] 
	,\sa_snapshot[20].r.part0[5] ,\sa_snapshot[20].r.part0[4] 
	,\sa_snapshot[20].r.part0[3] ,\sa_snapshot[20].r.part0[2] 
	,\sa_snapshot[20].r.part0[1] ,\sa_snapshot[20].r.part0[0] 
	,\sa_snapshot[19].r.part1[31] ,\sa_snapshot[19].r.part1[30] 
	,\sa_snapshot[19].r.part1[29] ,\sa_snapshot[19].r.part1[28] 
	,\sa_snapshot[19].r.part1[27] ,\sa_snapshot[19].r.part1[26] 
	,\sa_snapshot[19].r.part1[25] ,\sa_snapshot[19].r.part1[24] 
	,\sa_snapshot[19].r.part1[23] ,\sa_snapshot[19].r.part1[22] 
	,\sa_snapshot[19].r.part1[21] ,\sa_snapshot[19].r.part1[20] 
	,\sa_snapshot[19].r.part1[19] ,\sa_snapshot[19].r.part1[18] 
	,\sa_snapshot[19].r.part1[17] ,\sa_snapshot[19].r.part1[16] 
	,\sa_snapshot[19].r.part1[15] ,\sa_snapshot[19].r.part1[14] 
	,\sa_snapshot[19].r.part1[13] ,\sa_snapshot[19].r.part1[12] 
	,\sa_snapshot[19].r.part1[11] ,\sa_snapshot[19].r.part1[10] 
	,\sa_snapshot[19].r.part1[9] ,\sa_snapshot[19].r.part1[8] 
	,\sa_snapshot[19].r.part1[7] ,\sa_snapshot[19].r.part1[6] 
	,\sa_snapshot[19].r.part1[5] ,\sa_snapshot[19].r.part1[4] 
	,\sa_snapshot[19].r.part1[3] ,\sa_snapshot[19].r.part1[2] 
	,\sa_snapshot[19].r.part1[1] ,\sa_snapshot[19].r.part1[0] 
	,\sa_snapshot[19].r.part0[31] ,\sa_snapshot[19].r.part0[30] 
	,\sa_snapshot[19].r.part0[29] ,\sa_snapshot[19].r.part0[28] 
	,\sa_snapshot[19].r.part0[27] ,\sa_snapshot[19].r.part0[26] 
	,\sa_snapshot[19].r.part0[25] ,\sa_snapshot[19].r.part0[24] 
	,\sa_snapshot[19].r.part0[23] ,\sa_snapshot[19].r.part0[22] 
	,\sa_snapshot[19].r.part0[21] ,\sa_snapshot[19].r.part0[20] 
	,\sa_snapshot[19].r.part0[19] ,\sa_snapshot[19].r.part0[18] 
	,\sa_snapshot[19].r.part0[17] ,\sa_snapshot[19].r.part0[16] 
	,\sa_snapshot[19].r.part0[15] ,\sa_snapshot[19].r.part0[14] 
	,\sa_snapshot[19].r.part0[13] ,\sa_snapshot[19].r.part0[12] 
	,\sa_snapshot[19].r.part0[11] ,\sa_snapshot[19].r.part0[10] 
	,\sa_snapshot[19].r.part0[9] ,\sa_snapshot[19].r.part0[8] 
	,\sa_snapshot[19].r.part0[7] ,\sa_snapshot[19].r.part0[6] 
	,\sa_snapshot[19].r.part0[5] ,\sa_snapshot[19].r.part0[4] 
	,\sa_snapshot[19].r.part0[3] ,\sa_snapshot[19].r.part0[2] 
	,\sa_snapshot[19].r.part0[1] ,\sa_snapshot[19].r.part0[0] 
	,\sa_snapshot[18].r.part1[31] ,\sa_snapshot[18].r.part1[30] 
	,\sa_snapshot[18].r.part1[29] ,\sa_snapshot[18].r.part1[28] 
	,\sa_snapshot[18].r.part1[27] ,\sa_snapshot[18].r.part1[26] 
	,\sa_snapshot[18].r.part1[25] ,\sa_snapshot[18].r.part1[24] 
	,\sa_snapshot[18].r.part1[23] ,\sa_snapshot[18].r.part1[22] 
	,\sa_snapshot[18].r.part1[21] ,\sa_snapshot[18].r.part1[20] 
	,\sa_snapshot[18].r.part1[19] ,\sa_snapshot[18].r.part1[18] 
	,\sa_snapshot[18].r.part1[17] ,\sa_snapshot[18].r.part1[16] 
	,\sa_snapshot[18].r.part1[15] ,\sa_snapshot[18].r.part1[14] 
	,\sa_snapshot[18].r.part1[13] ,\sa_snapshot[18].r.part1[12] 
	,\sa_snapshot[18].r.part1[11] ,\sa_snapshot[18].r.part1[10] 
	,\sa_snapshot[18].r.part1[9] ,\sa_snapshot[18].r.part1[8] 
	,\sa_snapshot[18].r.part1[7] ,\sa_snapshot[18].r.part1[6] 
	,\sa_snapshot[18].r.part1[5] ,\sa_snapshot[18].r.part1[4] 
	,\sa_snapshot[18].r.part1[3] ,\sa_snapshot[18].r.part1[2] 
	,\sa_snapshot[18].r.part1[1] ,\sa_snapshot[18].r.part1[0] 
	,\sa_snapshot[18].r.part0[31] ,\sa_snapshot[18].r.part0[30] 
	,\sa_snapshot[18].r.part0[29] ,\sa_snapshot[18].r.part0[28] 
	,\sa_snapshot[18].r.part0[27] ,\sa_snapshot[18].r.part0[26] 
	,\sa_snapshot[18].r.part0[25] ,\sa_snapshot[18].r.part0[24] 
	,\sa_snapshot[18].r.part0[23] ,\sa_snapshot[18].r.part0[22] 
	,\sa_snapshot[18].r.part0[21] ,\sa_snapshot[18].r.part0[20] 
	,\sa_snapshot[18].r.part0[19] ,\sa_snapshot[18].r.part0[18] 
	,\sa_snapshot[18].r.part0[17] ,\sa_snapshot[18].r.part0[16] 
	,\sa_snapshot[18].r.part0[15] ,\sa_snapshot[18].r.part0[14] 
	,\sa_snapshot[18].r.part0[13] ,\sa_snapshot[18].r.part0[12] 
	,\sa_snapshot[18].r.part0[11] ,\sa_snapshot[18].r.part0[10] 
	,\sa_snapshot[18].r.part0[9] ,\sa_snapshot[18].r.part0[8] 
	,\sa_snapshot[18].r.part0[7] ,\sa_snapshot[18].r.part0[6] 
	,\sa_snapshot[18].r.part0[5] ,\sa_snapshot[18].r.part0[4] 
	,\sa_snapshot[18].r.part0[3] ,\sa_snapshot[18].r.part0[2] 
	,\sa_snapshot[18].r.part0[1] ,\sa_snapshot[18].r.part0[0] 
	,\sa_snapshot[17].r.part1[31] ,\sa_snapshot[17].r.part1[30] 
	,\sa_snapshot[17].r.part1[29] ,\sa_snapshot[17].r.part1[28] 
	,\sa_snapshot[17].r.part1[27] ,\sa_snapshot[17].r.part1[26] 
	,\sa_snapshot[17].r.part1[25] ,\sa_snapshot[17].r.part1[24] 
	,\sa_snapshot[17].r.part1[23] ,\sa_snapshot[17].r.part1[22] 
	,\sa_snapshot[17].r.part1[21] ,\sa_snapshot[17].r.part1[20] 
	,\sa_snapshot[17].r.part1[19] ,\sa_snapshot[17].r.part1[18] 
	,\sa_snapshot[17].r.part1[17] ,\sa_snapshot[17].r.part1[16] 
	,\sa_snapshot[17].r.part1[15] ,\sa_snapshot[17].r.part1[14] 
	,\sa_snapshot[17].r.part1[13] ,\sa_snapshot[17].r.part1[12] 
	,\sa_snapshot[17].r.part1[11] ,\sa_snapshot[17].r.part1[10] 
	,\sa_snapshot[17].r.part1[9] ,\sa_snapshot[17].r.part1[8] 
	,\sa_snapshot[17].r.part1[7] ,\sa_snapshot[17].r.part1[6] 
	,\sa_snapshot[17].r.part1[5] ,\sa_snapshot[17].r.part1[4] 
	,\sa_snapshot[17].r.part1[3] ,\sa_snapshot[17].r.part1[2] 
	,\sa_snapshot[17].r.part1[1] ,\sa_snapshot[17].r.part1[0] 
	,\sa_snapshot[17].r.part0[31] ,\sa_snapshot[17].r.part0[30] 
	,\sa_snapshot[17].r.part0[29] ,\sa_snapshot[17].r.part0[28] 
	,\sa_snapshot[17].r.part0[27] ,\sa_snapshot[17].r.part0[26] 
	,\sa_snapshot[17].r.part0[25] ,\sa_snapshot[17].r.part0[24] 
	,\sa_snapshot[17].r.part0[23] ,\sa_snapshot[17].r.part0[22] 
	,\sa_snapshot[17].r.part0[21] ,\sa_snapshot[17].r.part0[20] 
	,\sa_snapshot[17].r.part0[19] ,\sa_snapshot[17].r.part0[18] 
	,\sa_snapshot[17].r.part0[17] ,\sa_snapshot[17].r.part0[16] 
	,\sa_snapshot[17].r.part0[15] ,\sa_snapshot[17].r.part0[14] 
	,\sa_snapshot[17].r.part0[13] ,\sa_snapshot[17].r.part0[12] 
	,\sa_snapshot[17].r.part0[11] ,\sa_snapshot[17].r.part0[10] 
	,\sa_snapshot[17].r.part0[9] ,\sa_snapshot[17].r.part0[8] 
	,\sa_snapshot[17].r.part0[7] ,\sa_snapshot[17].r.part0[6] 
	,\sa_snapshot[17].r.part0[5] ,\sa_snapshot[17].r.part0[4] 
	,\sa_snapshot[17].r.part0[3] ,\sa_snapshot[17].r.part0[2] 
	,\sa_snapshot[17].r.part0[1] ,\sa_snapshot[17].r.part0[0] 
	,\sa_snapshot[16].r.part1[31] ,\sa_snapshot[16].r.part1[30] 
	,\sa_snapshot[16].r.part1[29] ,\sa_snapshot[16].r.part1[28] 
	,\sa_snapshot[16].r.part1[27] ,\sa_snapshot[16].r.part1[26] 
	,\sa_snapshot[16].r.part1[25] ,\sa_snapshot[16].r.part1[24] 
	,\sa_snapshot[16].r.part1[23] ,\sa_snapshot[16].r.part1[22] 
	,\sa_snapshot[16].r.part1[21] ,\sa_snapshot[16].r.part1[20] 
	,\sa_snapshot[16].r.part1[19] ,\sa_snapshot[16].r.part1[18] 
	,\sa_snapshot[16].r.part1[17] ,\sa_snapshot[16].r.part1[16] 
	,\sa_snapshot[16].r.part1[15] ,\sa_snapshot[16].r.part1[14] 
	,\sa_snapshot[16].r.part1[13] ,\sa_snapshot[16].r.part1[12] 
	,\sa_snapshot[16].r.part1[11] ,\sa_snapshot[16].r.part1[10] 
	,\sa_snapshot[16].r.part1[9] ,\sa_snapshot[16].r.part1[8] 
	,\sa_snapshot[16].r.part1[7] ,\sa_snapshot[16].r.part1[6] 
	,\sa_snapshot[16].r.part1[5] ,\sa_snapshot[16].r.part1[4] 
	,\sa_snapshot[16].r.part1[3] ,\sa_snapshot[16].r.part1[2] 
	,\sa_snapshot[16].r.part1[1] ,\sa_snapshot[16].r.part1[0] 
	,\sa_snapshot[16].r.part0[31] ,\sa_snapshot[16].r.part0[30] 
	,\sa_snapshot[16].r.part0[29] ,\sa_snapshot[16].r.part0[28] 
	,\sa_snapshot[16].r.part0[27] ,\sa_snapshot[16].r.part0[26] 
	,\sa_snapshot[16].r.part0[25] ,\sa_snapshot[16].r.part0[24] 
	,\sa_snapshot[16].r.part0[23] ,\sa_snapshot[16].r.part0[22] 
	,\sa_snapshot[16].r.part0[21] ,\sa_snapshot[16].r.part0[20] 
	,\sa_snapshot[16].r.part0[19] ,\sa_snapshot[16].r.part0[18] 
	,\sa_snapshot[16].r.part0[17] ,\sa_snapshot[16].r.part0[16] 
	,\sa_snapshot[16].r.part0[15] ,\sa_snapshot[16].r.part0[14] 
	,\sa_snapshot[16].r.part0[13] ,\sa_snapshot[16].r.part0[12] 
	,\sa_snapshot[16].r.part0[11] ,\sa_snapshot[16].r.part0[10] 
	,\sa_snapshot[16].r.part0[9] ,\sa_snapshot[16].r.part0[8] 
	,\sa_snapshot[16].r.part0[7] ,\sa_snapshot[16].r.part0[6] 
	,\sa_snapshot[16].r.part0[5] ,\sa_snapshot[16].r.part0[4] 
	,\sa_snapshot[16].r.part0[3] ,\sa_snapshot[16].r.part0[2] 
	,\sa_snapshot[16].r.part0[1] ,\sa_snapshot[16].r.part0[0] 
	,\sa_snapshot[15].r.part1[31] ,\sa_snapshot[15].r.part1[30] 
	,\sa_snapshot[15].r.part1[29] ,\sa_snapshot[15].r.part1[28] 
	,\sa_snapshot[15].r.part1[27] ,\sa_snapshot[15].r.part1[26] 
	,\sa_snapshot[15].r.part1[25] ,\sa_snapshot[15].r.part1[24] 
	,\sa_snapshot[15].r.part1[23] ,\sa_snapshot[15].r.part1[22] 
	,\sa_snapshot[15].r.part1[21] ,\sa_snapshot[15].r.part1[20] 
	,\sa_snapshot[15].r.part1[19] ,\sa_snapshot[15].r.part1[18] 
	,\sa_snapshot[15].r.part1[17] ,\sa_snapshot[15].r.part1[16] 
	,\sa_snapshot[15].r.part1[15] ,\sa_snapshot[15].r.part1[14] 
	,\sa_snapshot[15].r.part1[13] ,\sa_snapshot[15].r.part1[12] 
	,\sa_snapshot[15].r.part1[11] ,\sa_snapshot[15].r.part1[10] 
	,\sa_snapshot[15].r.part1[9] ,\sa_snapshot[15].r.part1[8] 
	,\sa_snapshot[15].r.part1[7] ,\sa_snapshot[15].r.part1[6] 
	,\sa_snapshot[15].r.part1[5] ,\sa_snapshot[15].r.part1[4] 
	,\sa_snapshot[15].r.part1[3] ,\sa_snapshot[15].r.part1[2] 
	,\sa_snapshot[15].r.part1[1] ,\sa_snapshot[15].r.part1[0] 
	,\sa_snapshot[15].r.part0[31] ,\sa_snapshot[15].r.part0[30] 
	,\sa_snapshot[15].r.part0[29] ,\sa_snapshot[15].r.part0[28] 
	,\sa_snapshot[15].r.part0[27] ,\sa_snapshot[15].r.part0[26] 
	,\sa_snapshot[15].r.part0[25] ,\sa_snapshot[15].r.part0[24] 
	,\sa_snapshot[15].r.part0[23] ,\sa_snapshot[15].r.part0[22] 
	,\sa_snapshot[15].r.part0[21] ,\sa_snapshot[15].r.part0[20] 
	,\sa_snapshot[15].r.part0[19] ,\sa_snapshot[15].r.part0[18] 
	,\sa_snapshot[15].r.part0[17] ,\sa_snapshot[15].r.part0[16] 
	,\sa_snapshot[15].r.part0[15] ,\sa_snapshot[15].r.part0[14] 
	,\sa_snapshot[15].r.part0[13] ,\sa_snapshot[15].r.part0[12] 
	,\sa_snapshot[15].r.part0[11] ,\sa_snapshot[15].r.part0[10] 
	,\sa_snapshot[15].r.part0[9] ,\sa_snapshot[15].r.part0[8] 
	,\sa_snapshot[15].r.part0[7] ,\sa_snapshot[15].r.part0[6] 
	,\sa_snapshot[15].r.part0[5] ,\sa_snapshot[15].r.part0[4] 
	,\sa_snapshot[15].r.part0[3] ,\sa_snapshot[15].r.part0[2] 
	,\sa_snapshot[15].r.part0[1] ,\sa_snapshot[15].r.part0[0] 
	,\sa_snapshot[14].r.part1[31] ,\sa_snapshot[14].r.part1[30] 
	,\sa_snapshot[14].r.part1[29] ,\sa_snapshot[14].r.part1[28] 
	,\sa_snapshot[14].r.part1[27] ,\sa_snapshot[14].r.part1[26] 
	,\sa_snapshot[14].r.part1[25] ,\sa_snapshot[14].r.part1[24] 
	,\sa_snapshot[14].r.part1[23] ,\sa_snapshot[14].r.part1[22] 
	,\sa_snapshot[14].r.part1[21] ,\sa_snapshot[14].r.part1[20] 
	,\sa_snapshot[14].r.part1[19] ,\sa_snapshot[14].r.part1[18] 
	,\sa_snapshot[14].r.part1[17] ,\sa_snapshot[14].r.part1[16] 
	,\sa_snapshot[14].r.part1[15] ,\sa_snapshot[14].r.part1[14] 
	,\sa_snapshot[14].r.part1[13] ,\sa_snapshot[14].r.part1[12] 
	,\sa_snapshot[14].r.part1[11] ,\sa_snapshot[14].r.part1[10] 
	,\sa_snapshot[14].r.part1[9] ,\sa_snapshot[14].r.part1[8] 
	,\sa_snapshot[14].r.part1[7] ,\sa_snapshot[14].r.part1[6] 
	,\sa_snapshot[14].r.part1[5] ,\sa_snapshot[14].r.part1[4] 
	,\sa_snapshot[14].r.part1[3] ,\sa_snapshot[14].r.part1[2] 
	,\sa_snapshot[14].r.part1[1] ,\sa_snapshot[14].r.part1[0] 
	,\sa_snapshot[14].r.part0[31] ,\sa_snapshot[14].r.part0[30] 
	,\sa_snapshot[14].r.part0[29] ,\sa_snapshot[14].r.part0[28] 
	,\sa_snapshot[14].r.part0[27] ,\sa_snapshot[14].r.part0[26] 
	,\sa_snapshot[14].r.part0[25] ,\sa_snapshot[14].r.part0[24] 
	,\sa_snapshot[14].r.part0[23] ,\sa_snapshot[14].r.part0[22] 
	,\sa_snapshot[14].r.part0[21] ,\sa_snapshot[14].r.part0[20] 
	,\sa_snapshot[14].r.part0[19] ,\sa_snapshot[14].r.part0[18] 
	,\sa_snapshot[14].r.part0[17] ,\sa_snapshot[14].r.part0[16] 
	,\sa_snapshot[14].r.part0[15] ,\sa_snapshot[14].r.part0[14] 
	,\sa_snapshot[14].r.part0[13] ,\sa_snapshot[14].r.part0[12] 
	,\sa_snapshot[14].r.part0[11] ,\sa_snapshot[14].r.part0[10] 
	,\sa_snapshot[14].r.part0[9] ,\sa_snapshot[14].r.part0[8] 
	,\sa_snapshot[14].r.part0[7] ,\sa_snapshot[14].r.part0[6] 
	,\sa_snapshot[14].r.part0[5] ,\sa_snapshot[14].r.part0[4] 
	,\sa_snapshot[14].r.part0[3] ,\sa_snapshot[14].r.part0[2] 
	,\sa_snapshot[14].r.part0[1] ,\sa_snapshot[14].r.part0[0] 
	,\sa_snapshot[13].r.part1[31] ,\sa_snapshot[13].r.part1[30] 
	,\sa_snapshot[13].r.part1[29] ,\sa_snapshot[13].r.part1[28] 
	,\sa_snapshot[13].r.part1[27] ,\sa_snapshot[13].r.part1[26] 
	,\sa_snapshot[13].r.part1[25] ,\sa_snapshot[13].r.part1[24] 
	,\sa_snapshot[13].r.part1[23] ,\sa_snapshot[13].r.part1[22] 
	,\sa_snapshot[13].r.part1[21] ,\sa_snapshot[13].r.part1[20] 
	,\sa_snapshot[13].r.part1[19] ,\sa_snapshot[13].r.part1[18] 
	,\sa_snapshot[13].r.part1[17] ,\sa_snapshot[13].r.part1[16] 
	,\sa_snapshot[13].r.part1[15] ,\sa_snapshot[13].r.part1[14] 
	,\sa_snapshot[13].r.part1[13] ,\sa_snapshot[13].r.part1[12] 
	,\sa_snapshot[13].r.part1[11] ,\sa_snapshot[13].r.part1[10] 
	,\sa_snapshot[13].r.part1[9] ,\sa_snapshot[13].r.part1[8] 
	,\sa_snapshot[13].r.part1[7] ,\sa_snapshot[13].r.part1[6] 
	,\sa_snapshot[13].r.part1[5] ,\sa_snapshot[13].r.part1[4] 
	,\sa_snapshot[13].r.part1[3] ,\sa_snapshot[13].r.part1[2] 
	,\sa_snapshot[13].r.part1[1] ,\sa_snapshot[13].r.part1[0] 
	,\sa_snapshot[13].r.part0[31] ,\sa_snapshot[13].r.part0[30] 
	,\sa_snapshot[13].r.part0[29] ,\sa_snapshot[13].r.part0[28] 
	,\sa_snapshot[13].r.part0[27] ,\sa_snapshot[13].r.part0[26] 
	,\sa_snapshot[13].r.part0[25] ,\sa_snapshot[13].r.part0[24] 
	,\sa_snapshot[13].r.part0[23] ,\sa_snapshot[13].r.part0[22] 
	,\sa_snapshot[13].r.part0[21] ,\sa_snapshot[13].r.part0[20] 
	,\sa_snapshot[13].r.part0[19] ,\sa_snapshot[13].r.part0[18] 
	,\sa_snapshot[13].r.part0[17] ,\sa_snapshot[13].r.part0[16] 
	,\sa_snapshot[13].r.part0[15] ,\sa_snapshot[13].r.part0[14] 
	,\sa_snapshot[13].r.part0[13] ,\sa_snapshot[13].r.part0[12] 
	,\sa_snapshot[13].r.part0[11] ,\sa_snapshot[13].r.part0[10] 
	,\sa_snapshot[13].r.part0[9] ,\sa_snapshot[13].r.part0[8] 
	,\sa_snapshot[13].r.part0[7] ,\sa_snapshot[13].r.part0[6] 
	,\sa_snapshot[13].r.part0[5] ,\sa_snapshot[13].r.part0[4] 
	,\sa_snapshot[13].r.part0[3] ,\sa_snapshot[13].r.part0[2] 
	,\sa_snapshot[13].r.part0[1] ,\sa_snapshot[13].r.part0[0] 
	,\sa_snapshot[12].r.part1[31] ,\sa_snapshot[12].r.part1[30] 
	,\sa_snapshot[12].r.part1[29] ,\sa_snapshot[12].r.part1[28] 
	,\sa_snapshot[12].r.part1[27] ,\sa_snapshot[12].r.part1[26] 
	,\sa_snapshot[12].r.part1[25] ,\sa_snapshot[12].r.part1[24] 
	,\sa_snapshot[12].r.part1[23] ,\sa_snapshot[12].r.part1[22] 
	,\sa_snapshot[12].r.part1[21] ,\sa_snapshot[12].r.part1[20] 
	,\sa_snapshot[12].r.part1[19] ,\sa_snapshot[12].r.part1[18] 
	,\sa_snapshot[12].r.part1[17] ,\sa_snapshot[12].r.part1[16] 
	,\sa_snapshot[12].r.part1[15] ,\sa_snapshot[12].r.part1[14] 
	,\sa_snapshot[12].r.part1[13] ,\sa_snapshot[12].r.part1[12] 
	,\sa_snapshot[12].r.part1[11] ,\sa_snapshot[12].r.part1[10] 
	,\sa_snapshot[12].r.part1[9] ,\sa_snapshot[12].r.part1[8] 
	,\sa_snapshot[12].r.part1[7] ,\sa_snapshot[12].r.part1[6] 
	,\sa_snapshot[12].r.part1[5] ,\sa_snapshot[12].r.part1[4] 
	,\sa_snapshot[12].r.part1[3] ,\sa_snapshot[12].r.part1[2] 
	,\sa_snapshot[12].r.part1[1] ,\sa_snapshot[12].r.part1[0] 
	,\sa_snapshot[12].r.part0[31] ,\sa_snapshot[12].r.part0[30] 
	,\sa_snapshot[12].r.part0[29] ,\sa_snapshot[12].r.part0[28] 
	,\sa_snapshot[12].r.part0[27] ,\sa_snapshot[12].r.part0[26] 
	,\sa_snapshot[12].r.part0[25] ,\sa_snapshot[12].r.part0[24] 
	,\sa_snapshot[12].r.part0[23] ,\sa_snapshot[12].r.part0[22] 
	,\sa_snapshot[12].r.part0[21] ,\sa_snapshot[12].r.part0[20] 
	,\sa_snapshot[12].r.part0[19] ,\sa_snapshot[12].r.part0[18] 
	,\sa_snapshot[12].r.part0[17] ,\sa_snapshot[12].r.part0[16] 
	,\sa_snapshot[12].r.part0[15] ,\sa_snapshot[12].r.part0[14] 
	,\sa_snapshot[12].r.part0[13] ,\sa_snapshot[12].r.part0[12] 
	,\sa_snapshot[12].r.part0[11] ,\sa_snapshot[12].r.part0[10] 
	,\sa_snapshot[12].r.part0[9] ,\sa_snapshot[12].r.part0[8] 
	,\sa_snapshot[12].r.part0[7] ,\sa_snapshot[12].r.part0[6] 
	,\sa_snapshot[12].r.part0[5] ,\sa_snapshot[12].r.part0[4] 
	,\sa_snapshot[12].r.part0[3] ,\sa_snapshot[12].r.part0[2] 
	,\sa_snapshot[12].r.part0[1] ,\sa_snapshot[12].r.part0[0] 
	,\sa_snapshot[11].r.part1[31] ,\sa_snapshot[11].r.part1[30] 
	,\sa_snapshot[11].r.part1[29] ,\sa_snapshot[11].r.part1[28] 
	,\sa_snapshot[11].r.part1[27] ,\sa_snapshot[11].r.part1[26] 
	,\sa_snapshot[11].r.part1[25] ,\sa_snapshot[11].r.part1[24] 
	,\sa_snapshot[11].r.part1[23] ,\sa_snapshot[11].r.part1[22] 
	,\sa_snapshot[11].r.part1[21] ,\sa_snapshot[11].r.part1[20] 
	,\sa_snapshot[11].r.part1[19] ,\sa_snapshot[11].r.part1[18] 
	,\sa_snapshot[11].r.part1[17] ,\sa_snapshot[11].r.part1[16] 
	,\sa_snapshot[11].r.part1[15] ,\sa_snapshot[11].r.part1[14] 
	,\sa_snapshot[11].r.part1[13] ,\sa_snapshot[11].r.part1[12] 
	,\sa_snapshot[11].r.part1[11] ,\sa_snapshot[11].r.part1[10] 
	,\sa_snapshot[11].r.part1[9] ,\sa_snapshot[11].r.part1[8] 
	,\sa_snapshot[11].r.part1[7] ,\sa_snapshot[11].r.part1[6] 
	,\sa_snapshot[11].r.part1[5] ,\sa_snapshot[11].r.part1[4] 
	,\sa_snapshot[11].r.part1[3] ,\sa_snapshot[11].r.part1[2] 
	,\sa_snapshot[11].r.part1[1] ,\sa_snapshot[11].r.part1[0] 
	,\sa_snapshot[11].r.part0[31] ,\sa_snapshot[11].r.part0[30] 
	,\sa_snapshot[11].r.part0[29] ,\sa_snapshot[11].r.part0[28] 
	,\sa_snapshot[11].r.part0[27] ,\sa_snapshot[11].r.part0[26] 
	,\sa_snapshot[11].r.part0[25] ,\sa_snapshot[11].r.part0[24] 
	,\sa_snapshot[11].r.part0[23] ,\sa_snapshot[11].r.part0[22] 
	,\sa_snapshot[11].r.part0[21] ,\sa_snapshot[11].r.part0[20] 
	,\sa_snapshot[11].r.part0[19] ,\sa_snapshot[11].r.part0[18] 
	,\sa_snapshot[11].r.part0[17] ,\sa_snapshot[11].r.part0[16] 
	,\sa_snapshot[11].r.part0[15] ,\sa_snapshot[11].r.part0[14] 
	,\sa_snapshot[11].r.part0[13] ,\sa_snapshot[11].r.part0[12] 
	,\sa_snapshot[11].r.part0[11] ,\sa_snapshot[11].r.part0[10] 
	,\sa_snapshot[11].r.part0[9] ,\sa_snapshot[11].r.part0[8] 
	,\sa_snapshot[11].r.part0[7] ,\sa_snapshot[11].r.part0[6] 
	,\sa_snapshot[11].r.part0[5] ,\sa_snapshot[11].r.part0[4] 
	,\sa_snapshot[11].r.part0[3] ,\sa_snapshot[11].r.part0[2] 
	,\sa_snapshot[11].r.part0[1] ,\sa_snapshot[11].r.part0[0] 
	,\sa_snapshot[10].r.part1[31] ,\sa_snapshot[10].r.part1[30] 
	,\sa_snapshot[10].r.part1[29] ,\sa_snapshot[10].r.part1[28] 
	,\sa_snapshot[10].r.part1[27] ,\sa_snapshot[10].r.part1[26] 
	,\sa_snapshot[10].r.part1[25] ,\sa_snapshot[10].r.part1[24] 
	,\sa_snapshot[10].r.part1[23] ,\sa_snapshot[10].r.part1[22] 
	,\sa_snapshot[10].r.part1[21] ,\sa_snapshot[10].r.part1[20] 
	,\sa_snapshot[10].r.part1[19] ,\sa_snapshot[10].r.part1[18] 
	,\sa_snapshot[10].r.part1[17] ,\sa_snapshot[10].r.part1[16] 
	,\sa_snapshot[10].r.part1[15] ,\sa_snapshot[10].r.part1[14] 
	,\sa_snapshot[10].r.part1[13] ,\sa_snapshot[10].r.part1[12] 
	,\sa_snapshot[10].r.part1[11] ,\sa_snapshot[10].r.part1[10] 
	,\sa_snapshot[10].r.part1[9] ,\sa_snapshot[10].r.part1[8] 
	,\sa_snapshot[10].r.part1[7] ,\sa_snapshot[10].r.part1[6] 
	,\sa_snapshot[10].r.part1[5] ,\sa_snapshot[10].r.part1[4] 
	,\sa_snapshot[10].r.part1[3] ,\sa_snapshot[10].r.part1[2] 
	,\sa_snapshot[10].r.part1[1] ,\sa_snapshot[10].r.part1[0] 
	,\sa_snapshot[10].r.part0[31] ,\sa_snapshot[10].r.part0[30] 
	,\sa_snapshot[10].r.part0[29] ,\sa_snapshot[10].r.part0[28] 
	,\sa_snapshot[10].r.part0[27] ,\sa_snapshot[10].r.part0[26] 
	,\sa_snapshot[10].r.part0[25] ,\sa_snapshot[10].r.part0[24] 
	,\sa_snapshot[10].r.part0[23] ,\sa_snapshot[10].r.part0[22] 
	,\sa_snapshot[10].r.part0[21] ,\sa_snapshot[10].r.part0[20] 
	,\sa_snapshot[10].r.part0[19] ,\sa_snapshot[10].r.part0[18] 
	,\sa_snapshot[10].r.part0[17] ,\sa_snapshot[10].r.part0[16] 
	,\sa_snapshot[10].r.part0[15] ,\sa_snapshot[10].r.part0[14] 
	,\sa_snapshot[10].r.part0[13] ,\sa_snapshot[10].r.part0[12] 
	,\sa_snapshot[10].r.part0[11] ,\sa_snapshot[10].r.part0[10] 
	,\sa_snapshot[10].r.part0[9] ,\sa_snapshot[10].r.part0[8] 
	,\sa_snapshot[10].r.part0[7] ,\sa_snapshot[10].r.part0[6] 
	,\sa_snapshot[10].r.part0[5] ,\sa_snapshot[10].r.part0[4] 
	,\sa_snapshot[10].r.part0[3] ,\sa_snapshot[10].r.part0[2] 
	,\sa_snapshot[10].r.part0[1] ,\sa_snapshot[10].r.part0[0] 
	,\sa_snapshot[9].r.part1[31] ,\sa_snapshot[9].r.part1[30] 
	,\sa_snapshot[9].r.part1[29] ,\sa_snapshot[9].r.part1[28] 
	,\sa_snapshot[9].r.part1[27] ,\sa_snapshot[9].r.part1[26] 
	,\sa_snapshot[9].r.part1[25] ,\sa_snapshot[9].r.part1[24] 
	,\sa_snapshot[9].r.part1[23] ,\sa_snapshot[9].r.part1[22] 
	,\sa_snapshot[9].r.part1[21] ,\sa_snapshot[9].r.part1[20] 
	,\sa_snapshot[9].r.part1[19] ,\sa_snapshot[9].r.part1[18] 
	,\sa_snapshot[9].r.part1[17] ,\sa_snapshot[9].r.part1[16] 
	,\sa_snapshot[9].r.part1[15] ,\sa_snapshot[9].r.part1[14] 
	,\sa_snapshot[9].r.part1[13] ,\sa_snapshot[9].r.part1[12] 
	,\sa_snapshot[9].r.part1[11] ,\sa_snapshot[9].r.part1[10] 
	,\sa_snapshot[9].r.part1[9] ,\sa_snapshot[9].r.part1[8] 
	,\sa_snapshot[9].r.part1[7] ,\sa_snapshot[9].r.part1[6] 
	,\sa_snapshot[9].r.part1[5] ,\sa_snapshot[9].r.part1[4] 
	,\sa_snapshot[9].r.part1[3] ,\sa_snapshot[9].r.part1[2] 
	,\sa_snapshot[9].r.part1[1] ,\sa_snapshot[9].r.part1[0] 
	,\sa_snapshot[9].r.part0[31] ,\sa_snapshot[9].r.part0[30] 
	,\sa_snapshot[9].r.part0[29] ,\sa_snapshot[9].r.part0[28] 
	,\sa_snapshot[9].r.part0[27] ,\sa_snapshot[9].r.part0[26] 
	,\sa_snapshot[9].r.part0[25] ,\sa_snapshot[9].r.part0[24] 
	,\sa_snapshot[9].r.part0[23] ,\sa_snapshot[9].r.part0[22] 
	,\sa_snapshot[9].r.part0[21] ,\sa_snapshot[9].r.part0[20] 
	,\sa_snapshot[9].r.part0[19] ,\sa_snapshot[9].r.part0[18] 
	,\sa_snapshot[9].r.part0[17] ,\sa_snapshot[9].r.part0[16] 
	,\sa_snapshot[9].r.part0[15] ,\sa_snapshot[9].r.part0[14] 
	,\sa_snapshot[9].r.part0[13] ,\sa_snapshot[9].r.part0[12] 
	,\sa_snapshot[9].r.part0[11] ,\sa_snapshot[9].r.part0[10] 
	,\sa_snapshot[9].r.part0[9] ,\sa_snapshot[9].r.part0[8] 
	,\sa_snapshot[9].r.part0[7] ,\sa_snapshot[9].r.part0[6] 
	,\sa_snapshot[9].r.part0[5] ,\sa_snapshot[9].r.part0[4] 
	,\sa_snapshot[9].r.part0[3] ,\sa_snapshot[9].r.part0[2] 
	,\sa_snapshot[9].r.part0[1] ,\sa_snapshot[9].r.part0[0] 
	,\sa_snapshot[8].r.part1[31] ,\sa_snapshot[8].r.part1[30] 
	,\sa_snapshot[8].r.part1[29] ,\sa_snapshot[8].r.part1[28] 
	,\sa_snapshot[8].r.part1[27] ,\sa_snapshot[8].r.part1[26] 
	,\sa_snapshot[8].r.part1[25] ,\sa_snapshot[8].r.part1[24] 
	,\sa_snapshot[8].r.part1[23] ,\sa_snapshot[8].r.part1[22] 
	,\sa_snapshot[8].r.part1[21] ,\sa_snapshot[8].r.part1[20] 
	,\sa_snapshot[8].r.part1[19] ,\sa_snapshot[8].r.part1[18] 
	,\sa_snapshot[8].r.part1[17] ,\sa_snapshot[8].r.part1[16] 
	,\sa_snapshot[8].r.part1[15] ,\sa_snapshot[8].r.part1[14] 
	,\sa_snapshot[8].r.part1[13] ,\sa_snapshot[8].r.part1[12] 
	,\sa_snapshot[8].r.part1[11] ,\sa_snapshot[8].r.part1[10] 
	,\sa_snapshot[8].r.part1[9] ,\sa_snapshot[8].r.part1[8] 
	,\sa_snapshot[8].r.part1[7] ,\sa_snapshot[8].r.part1[6] 
	,\sa_snapshot[8].r.part1[5] ,\sa_snapshot[8].r.part1[4] 
	,\sa_snapshot[8].r.part1[3] ,\sa_snapshot[8].r.part1[2] 
	,\sa_snapshot[8].r.part1[1] ,\sa_snapshot[8].r.part1[0] 
	,\sa_snapshot[8].r.part0[31] ,\sa_snapshot[8].r.part0[30] 
	,\sa_snapshot[8].r.part0[29] ,\sa_snapshot[8].r.part0[28] 
	,\sa_snapshot[8].r.part0[27] ,\sa_snapshot[8].r.part0[26] 
	,\sa_snapshot[8].r.part0[25] ,\sa_snapshot[8].r.part0[24] 
	,\sa_snapshot[8].r.part0[23] ,\sa_snapshot[8].r.part0[22] 
	,\sa_snapshot[8].r.part0[21] ,\sa_snapshot[8].r.part0[20] 
	,\sa_snapshot[8].r.part0[19] ,\sa_snapshot[8].r.part0[18] 
	,\sa_snapshot[8].r.part0[17] ,\sa_snapshot[8].r.part0[16] 
	,\sa_snapshot[8].r.part0[15] ,\sa_snapshot[8].r.part0[14] 
	,\sa_snapshot[8].r.part0[13] ,\sa_snapshot[8].r.part0[12] 
	,\sa_snapshot[8].r.part0[11] ,\sa_snapshot[8].r.part0[10] 
	,\sa_snapshot[8].r.part0[9] ,\sa_snapshot[8].r.part0[8] 
	,\sa_snapshot[8].r.part0[7] ,\sa_snapshot[8].r.part0[6] 
	,\sa_snapshot[8].r.part0[5] ,\sa_snapshot[8].r.part0[4] 
	,\sa_snapshot[8].r.part0[3] ,\sa_snapshot[8].r.part0[2] 
	,\sa_snapshot[8].r.part0[1] ,\sa_snapshot[8].r.part0[0] 
	,\sa_snapshot[7].r.part1[31] ,\sa_snapshot[7].r.part1[30] 
	,\sa_snapshot[7].r.part1[29] ,\sa_snapshot[7].r.part1[28] 
	,\sa_snapshot[7].r.part1[27] ,\sa_snapshot[7].r.part1[26] 
	,\sa_snapshot[7].r.part1[25] ,\sa_snapshot[7].r.part1[24] 
	,\sa_snapshot[7].r.part1[23] ,\sa_snapshot[7].r.part1[22] 
	,\sa_snapshot[7].r.part1[21] ,\sa_snapshot[7].r.part1[20] 
	,\sa_snapshot[7].r.part1[19] ,\sa_snapshot[7].r.part1[18] 
	,\sa_snapshot[7].r.part1[17] ,\sa_snapshot[7].r.part1[16] 
	,\sa_snapshot[7].r.part1[15] ,\sa_snapshot[7].r.part1[14] 
	,\sa_snapshot[7].r.part1[13] ,\sa_snapshot[7].r.part1[12] 
	,\sa_snapshot[7].r.part1[11] ,\sa_snapshot[7].r.part1[10] 
	,\sa_snapshot[7].r.part1[9] ,\sa_snapshot[7].r.part1[8] 
	,\sa_snapshot[7].r.part1[7] ,\sa_snapshot[7].r.part1[6] 
	,\sa_snapshot[7].r.part1[5] ,\sa_snapshot[7].r.part1[4] 
	,\sa_snapshot[7].r.part1[3] ,\sa_snapshot[7].r.part1[2] 
	,\sa_snapshot[7].r.part1[1] ,\sa_snapshot[7].r.part1[0] 
	,\sa_snapshot[7].r.part0[31] ,\sa_snapshot[7].r.part0[30] 
	,\sa_snapshot[7].r.part0[29] ,\sa_snapshot[7].r.part0[28] 
	,\sa_snapshot[7].r.part0[27] ,\sa_snapshot[7].r.part0[26] 
	,\sa_snapshot[7].r.part0[25] ,\sa_snapshot[7].r.part0[24] 
	,\sa_snapshot[7].r.part0[23] ,\sa_snapshot[7].r.part0[22] 
	,\sa_snapshot[7].r.part0[21] ,\sa_snapshot[7].r.part0[20] 
	,\sa_snapshot[7].r.part0[19] ,\sa_snapshot[7].r.part0[18] 
	,\sa_snapshot[7].r.part0[17] ,\sa_snapshot[7].r.part0[16] 
	,\sa_snapshot[7].r.part0[15] ,\sa_snapshot[7].r.part0[14] 
	,\sa_snapshot[7].r.part0[13] ,\sa_snapshot[7].r.part0[12] 
	,\sa_snapshot[7].r.part0[11] ,\sa_snapshot[7].r.part0[10] 
	,\sa_snapshot[7].r.part0[9] ,\sa_snapshot[7].r.part0[8] 
	,\sa_snapshot[7].r.part0[7] ,\sa_snapshot[7].r.part0[6] 
	,\sa_snapshot[7].r.part0[5] ,\sa_snapshot[7].r.part0[4] 
	,\sa_snapshot[7].r.part0[3] ,\sa_snapshot[7].r.part0[2] 
	,\sa_snapshot[7].r.part0[1] ,\sa_snapshot[7].r.part0[0] 
	,\sa_snapshot[6].r.part1[31] ,\sa_snapshot[6].r.part1[30] 
	,\sa_snapshot[6].r.part1[29] ,\sa_snapshot[6].r.part1[28] 
	,\sa_snapshot[6].r.part1[27] ,\sa_snapshot[6].r.part1[26] 
	,\sa_snapshot[6].r.part1[25] ,\sa_snapshot[6].r.part1[24] 
	,\sa_snapshot[6].r.part1[23] ,\sa_snapshot[6].r.part1[22] 
	,\sa_snapshot[6].r.part1[21] ,\sa_snapshot[6].r.part1[20] 
	,\sa_snapshot[6].r.part1[19] ,\sa_snapshot[6].r.part1[18] 
	,\sa_snapshot[6].r.part1[17] ,\sa_snapshot[6].r.part1[16] 
	,\sa_snapshot[6].r.part1[15] ,\sa_snapshot[6].r.part1[14] 
	,\sa_snapshot[6].r.part1[13] ,\sa_snapshot[6].r.part1[12] 
	,\sa_snapshot[6].r.part1[11] ,\sa_snapshot[6].r.part1[10] 
	,\sa_snapshot[6].r.part1[9] ,\sa_snapshot[6].r.part1[8] 
	,\sa_snapshot[6].r.part1[7] ,\sa_snapshot[6].r.part1[6] 
	,\sa_snapshot[6].r.part1[5] ,\sa_snapshot[6].r.part1[4] 
	,\sa_snapshot[6].r.part1[3] ,\sa_snapshot[6].r.part1[2] 
	,\sa_snapshot[6].r.part1[1] ,\sa_snapshot[6].r.part1[0] 
	,\sa_snapshot[6].r.part0[31] ,\sa_snapshot[6].r.part0[30] 
	,\sa_snapshot[6].r.part0[29] ,\sa_snapshot[6].r.part0[28] 
	,\sa_snapshot[6].r.part0[27] ,\sa_snapshot[6].r.part0[26] 
	,\sa_snapshot[6].r.part0[25] ,\sa_snapshot[6].r.part0[24] 
	,\sa_snapshot[6].r.part0[23] ,\sa_snapshot[6].r.part0[22] 
	,\sa_snapshot[6].r.part0[21] ,\sa_snapshot[6].r.part0[20] 
	,\sa_snapshot[6].r.part0[19] ,\sa_snapshot[6].r.part0[18] 
	,\sa_snapshot[6].r.part0[17] ,\sa_snapshot[6].r.part0[16] 
	,\sa_snapshot[6].r.part0[15] ,\sa_snapshot[6].r.part0[14] 
	,\sa_snapshot[6].r.part0[13] ,\sa_snapshot[6].r.part0[12] 
	,\sa_snapshot[6].r.part0[11] ,\sa_snapshot[6].r.part0[10] 
	,\sa_snapshot[6].r.part0[9] ,\sa_snapshot[6].r.part0[8] 
	,\sa_snapshot[6].r.part0[7] ,\sa_snapshot[6].r.part0[6] 
	,\sa_snapshot[6].r.part0[5] ,\sa_snapshot[6].r.part0[4] 
	,\sa_snapshot[6].r.part0[3] ,\sa_snapshot[6].r.part0[2] 
	,\sa_snapshot[6].r.part0[1] ,\sa_snapshot[6].r.part0[0] 
	,\sa_snapshot[5].r.part1[31] ,\sa_snapshot[5].r.part1[30] 
	,\sa_snapshot[5].r.part1[29] ,\sa_snapshot[5].r.part1[28] 
	,\sa_snapshot[5].r.part1[27] ,\sa_snapshot[5].r.part1[26] 
	,\sa_snapshot[5].r.part1[25] ,\sa_snapshot[5].r.part1[24] 
	,\sa_snapshot[5].r.part1[23] ,\sa_snapshot[5].r.part1[22] 
	,\sa_snapshot[5].r.part1[21] ,\sa_snapshot[5].r.part1[20] 
	,\sa_snapshot[5].r.part1[19] ,\sa_snapshot[5].r.part1[18] 
	,\sa_snapshot[5].r.part1[17] ,\sa_snapshot[5].r.part1[16] 
	,\sa_snapshot[5].r.part1[15] ,\sa_snapshot[5].r.part1[14] 
	,\sa_snapshot[5].r.part1[13] ,\sa_snapshot[5].r.part1[12] 
	,\sa_snapshot[5].r.part1[11] ,\sa_snapshot[5].r.part1[10] 
	,\sa_snapshot[5].r.part1[9] ,\sa_snapshot[5].r.part1[8] 
	,\sa_snapshot[5].r.part1[7] ,\sa_snapshot[5].r.part1[6] 
	,\sa_snapshot[5].r.part1[5] ,\sa_snapshot[5].r.part1[4] 
	,\sa_snapshot[5].r.part1[3] ,\sa_snapshot[5].r.part1[2] 
	,\sa_snapshot[5].r.part1[1] ,\sa_snapshot[5].r.part1[0] 
	,\sa_snapshot[5].r.part0[31] ,\sa_snapshot[5].r.part0[30] 
	,\sa_snapshot[5].r.part0[29] ,\sa_snapshot[5].r.part0[28] 
	,\sa_snapshot[5].r.part0[27] ,\sa_snapshot[5].r.part0[26] 
	,\sa_snapshot[5].r.part0[25] ,\sa_snapshot[5].r.part0[24] 
	,\sa_snapshot[5].r.part0[23] ,\sa_snapshot[5].r.part0[22] 
	,\sa_snapshot[5].r.part0[21] ,\sa_snapshot[5].r.part0[20] 
	,\sa_snapshot[5].r.part0[19] ,\sa_snapshot[5].r.part0[18] 
	,\sa_snapshot[5].r.part0[17] ,\sa_snapshot[5].r.part0[16] 
	,\sa_snapshot[5].r.part0[15] ,\sa_snapshot[5].r.part0[14] 
	,\sa_snapshot[5].r.part0[13] ,\sa_snapshot[5].r.part0[12] 
	,\sa_snapshot[5].r.part0[11] ,\sa_snapshot[5].r.part0[10] 
	,\sa_snapshot[5].r.part0[9] ,\sa_snapshot[5].r.part0[8] 
	,\sa_snapshot[5].r.part0[7] ,\sa_snapshot[5].r.part0[6] 
	,\sa_snapshot[5].r.part0[5] ,\sa_snapshot[5].r.part0[4] 
	,\sa_snapshot[5].r.part0[3] ,\sa_snapshot[5].r.part0[2] 
	,\sa_snapshot[5].r.part0[1] ,\sa_snapshot[5].r.part0[0] 
	,\sa_snapshot[4].r.part1[31] ,\sa_snapshot[4].r.part1[30] 
	,\sa_snapshot[4].r.part1[29] ,\sa_snapshot[4].r.part1[28] 
	,\sa_snapshot[4].r.part1[27] ,\sa_snapshot[4].r.part1[26] 
	,\sa_snapshot[4].r.part1[25] ,\sa_snapshot[4].r.part1[24] 
	,\sa_snapshot[4].r.part1[23] ,\sa_snapshot[4].r.part1[22] 
	,\sa_snapshot[4].r.part1[21] ,\sa_snapshot[4].r.part1[20] 
	,\sa_snapshot[4].r.part1[19] ,\sa_snapshot[4].r.part1[18] 
	,\sa_snapshot[4].r.part1[17] ,\sa_snapshot[4].r.part1[16] 
	,\sa_snapshot[4].r.part1[15] ,\sa_snapshot[4].r.part1[14] 
	,\sa_snapshot[4].r.part1[13] ,\sa_snapshot[4].r.part1[12] 
	,\sa_snapshot[4].r.part1[11] ,\sa_snapshot[4].r.part1[10] 
	,\sa_snapshot[4].r.part1[9] ,\sa_snapshot[4].r.part1[8] 
	,\sa_snapshot[4].r.part1[7] ,\sa_snapshot[4].r.part1[6] 
	,\sa_snapshot[4].r.part1[5] ,\sa_snapshot[4].r.part1[4] 
	,\sa_snapshot[4].r.part1[3] ,\sa_snapshot[4].r.part1[2] 
	,\sa_snapshot[4].r.part1[1] ,\sa_snapshot[4].r.part1[0] 
	,\sa_snapshot[4].r.part0[31] ,\sa_snapshot[4].r.part0[30] 
	,\sa_snapshot[4].r.part0[29] ,\sa_snapshot[4].r.part0[28] 
	,\sa_snapshot[4].r.part0[27] ,\sa_snapshot[4].r.part0[26] 
	,\sa_snapshot[4].r.part0[25] ,\sa_snapshot[4].r.part0[24] 
	,\sa_snapshot[4].r.part0[23] ,\sa_snapshot[4].r.part0[22] 
	,\sa_snapshot[4].r.part0[21] ,\sa_snapshot[4].r.part0[20] 
	,\sa_snapshot[4].r.part0[19] ,\sa_snapshot[4].r.part0[18] 
	,\sa_snapshot[4].r.part0[17] ,\sa_snapshot[4].r.part0[16] 
	,\sa_snapshot[4].r.part0[15] ,\sa_snapshot[4].r.part0[14] 
	,\sa_snapshot[4].r.part0[13] ,\sa_snapshot[4].r.part0[12] 
	,\sa_snapshot[4].r.part0[11] ,\sa_snapshot[4].r.part0[10] 
	,\sa_snapshot[4].r.part0[9] ,\sa_snapshot[4].r.part0[8] 
	,\sa_snapshot[4].r.part0[7] ,\sa_snapshot[4].r.part0[6] 
	,\sa_snapshot[4].r.part0[5] ,\sa_snapshot[4].r.part0[4] 
	,\sa_snapshot[4].r.part0[3] ,\sa_snapshot[4].r.part0[2] 
	,\sa_snapshot[4].r.part0[1] ,\sa_snapshot[4].r.part0[0] 
	,\sa_snapshot[3].r.part1[31] ,\sa_snapshot[3].r.part1[30] 
	,\sa_snapshot[3].r.part1[29] ,\sa_snapshot[3].r.part1[28] 
	,\sa_snapshot[3].r.part1[27] ,\sa_snapshot[3].r.part1[26] 
	,\sa_snapshot[3].r.part1[25] ,\sa_snapshot[3].r.part1[24] 
	,\sa_snapshot[3].r.part1[23] ,\sa_snapshot[3].r.part1[22] 
	,\sa_snapshot[3].r.part1[21] ,\sa_snapshot[3].r.part1[20] 
	,\sa_snapshot[3].r.part1[19] ,\sa_snapshot[3].r.part1[18] 
	,\sa_snapshot[3].r.part1[17] ,\sa_snapshot[3].r.part1[16] 
	,\sa_snapshot[3].r.part1[15] ,\sa_snapshot[3].r.part1[14] 
	,\sa_snapshot[3].r.part1[13] ,\sa_snapshot[3].r.part1[12] 
	,\sa_snapshot[3].r.part1[11] ,\sa_snapshot[3].r.part1[10] 
	,\sa_snapshot[3].r.part1[9] ,\sa_snapshot[3].r.part1[8] 
	,\sa_snapshot[3].r.part1[7] ,\sa_snapshot[3].r.part1[6] 
	,\sa_snapshot[3].r.part1[5] ,\sa_snapshot[3].r.part1[4] 
	,\sa_snapshot[3].r.part1[3] ,\sa_snapshot[3].r.part1[2] 
	,\sa_snapshot[3].r.part1[1] ,\sa_snapshot[3].r.part1[0] 
	,\sa_snapshot[3].r.part0[31] ,\sa_snapshot[3].r.part0[30] 
	,\sa_snapshot[3].r.part0[29] ,\sa_snapshot[3].r.part0[28] 
	,\sa_snapshot[3].r.part0[27] ,\sa_snapshot[3].r.part0[26] 
	,\sa_snapshot[3].r.part0[25] ,\sa_snapshot[3].r.part0[24] 
	,\sa_snapshot[3].r.part0[23] ,\sa_snapshot[3].r.part0[22] 
	,\sa_snapshot[3].r.part0[21] ,\sa_snapshot[3].r.part0[20] 
	,\sa_snapshot[3].r.part0[19] ,\sa_snapshot[3].r.part0[18] 
	,\sa_snapshot[3].r.part0[17] ,\sa_snapshot[3].r.part0[16] 
	,\sa_snapshot[3].r.part0[15] ,\sa_snapshot[3].r.part0[14] 
	,\sa_snapshot[3].r.part0[13] ,\sa_snapshot[3].r.part0[12] 
	,\sa_snapshot[3].r.part0[11] ,\sa_snapshot[3].r.part0[10] 
	,\sa_snapshot[3].r.part0[9] ,\sa_snapshot[3].r.part0[8] 
	,\sa_snapshot[3].r.part0[7] ,\sa_snapshot[3].r.part0[6] 
	,\sa_snapshot[3].r.part0[5] ,\sa_snapshot[3].r.part0[4] 
	,\sa_snapshot[3].r.part0[3] ,\sa_snapshot[3].r.part0[2] 
	,\sa_snapshot[3].r.part0[1] ,\sa_snapshot[3].r.part0[0] 
	,\sa_snapshot[2].r.part1[31] ,\sa_snapshot[2].r.part1[30] 
	,\sa_snapshot[2].r.part1[29] ,\sa_snapshot[2].r.part1[28] 
	,\sa_snapshot[2].r.part1[27] ,\sa_snapshot[2].r.part1[26] 
	,\sa_snapshot[2].r.part1[25] ,\sa_snapshot[2].r.part1[24] 
	,\sa_snapshot[2].r.part1[23] ,\sa_snapshot[2].r.part1[22] 
	,\sa_snapshot[2].r.part1[21] ,\sa_snapshot[2].r.part1[20] 
	,\sa_snapshot[2].r.part1[19] ,\sa_snapshot[2].r.part1[18] 
	,\sa_snapshot[2].r.part1[17] ,\sa_snapshot[2].r.part1[16] 
	,\sa_snapshot[2].r.part1[15] ,\sa_snapshot[2].r.part1[14] 
	,\sa_snapshot[2].r.part1[13] ,\sa_snapshot[2].r.part1[12] 
	,\sa_snapshot[2].r.part1[11] ,\sa_snapshot[2].r.part1[10] 
	,\sa_snapshot[2].r.part1[9] ,\sa_snapshot[2].r.part1[8] 
	,\sa_snapshot[2].r.part1[7] ,\sa_snapshot[2].r.part1[6] 
	,\sa_snapshot[2].r.part1[5] ,\sa_snapshot[2].r.part1[4] 
	,\sa_snapshot[2].r.part1[3] ,\sa_snapshot[2].r.part1[2] 
	,\sa_snapshot[2].r.part1[1] ,\sa_snapshot[2].r.part1[0] 
	,\sa_snapshot[2].r.part0[31] ,\sa_snapshot[2].r.part0[30] 
	,\sa_snapshot[2].r.part0[29] ,\sa_snapshot[2].r.part0[28] 
	,\sa_snapshot[2].r.part0[27] ,\sa_snapshot[2].r.part0[26] 
	,\sa_snapshot[2].r.part0[25] ,\sa_snapshot[2].r.part0[24] 
	,\sa_snapshot[2].r.part0[23] ,\sa_snapshot[2].r.part0[22] 
	,\sa_snapshot[2].r.part0[21] ,\sa_snapshot[2].r.part0[20] 
	,\sa_snapshot[2].r.part0[19] ,\sa_snapshot[2].r.part0[18] 
	,\sa_snapshot[2].r.part0[17] ,\sa_snapshot[2].r.part0[16] 
	,\sa_snapshot[2].r.part0[15] ,\sa_snapshot[2].r.part0[14] 
	,\sa_snapshot[2].r.part0[13] ,\sa_snapshot[2].r.part0[12] 
	,\sa_snapshot[2].r.part0[11] ,\sa_snapshot[2].r.part0[10] 
	,\sa_snapshot[2].r.part0[9] ,\sa_snapshot[2].r.part0[8] 
	,\sa_snapshot[2].r.part0[7] ,\sa_snapshot[2].r.part0[6] 
	,\sa_snapshot[2].r.part0[5] ,\sa_snapshot[2].r.part0[4] 
	,\sa_snapshot[2].r.part0[3] ,\sa_snapshot[2].r.part0[2] 
	,\sa_snapshot[2].r.part0[1] ,\sa_snapshot[2].r.part0[0] 
	,\sa_snapshot[1].r.part1[31] ,\sa_snapshot[1].r.part1[30] 
	,\sa_snapshot[1].r.part1[29] ,\sa_snapshot[1].r.part1[28] 
	,\sa_snapshot[1].r.part1[27] ,\sa_snapshot[1].r.part1[26] 
	,\sa_snapshot[1].r.part1[25] ,\sa_snapshot[1].r.part1[24] 
	,\sa_snapshot[1].r.part1[23] ,\sa_snapshot[1].r.part1[22] 
	,\sa_snapshot[1].r.part1[21] ,\sa_snapshot[1].r.part1[20] 
	,\sa_snapshot[1].r.part1[19] ,\sa_snapshot[1].r.part1[18] 
	,\sa_snapshot[1].r.part1[17] ,\sa_snapshot[1].r.part1[16] 
	,\sa_snapshot[1].r.part1[15] ,\sa_snapshot[1].r.part1[14] 
	,\sa_snapshot[1].r.part1[13] ,\sa_snapshot[1].r.part1[12] 
	,\sa_snapshot[1].r.part1[11] ,\sa_snapshot[1].r.part1[10] 
	,\sa_snapshot[1].r.part1[9] ,\sa_snapshot[1].r.part1[8] 
	,\sa_snapshot[1].r.part1[7] ,\sa_snapshot[1].r.part1[6] 
	,\sa_snapshot[1].r.part1[5] ,\sa_snapshot[1].r.part1[4] 
	,\sa_snapshot[1].r.part1[3] ,\sa_snapshot[1].r.part1[2] 
	,\sa_snapshot[1].r.part1[1] ,\sa_snapshot[1].r.part1[0] 
	,\sa_snapshot[1].r.part0[31] ,\sa_snapshot[1].r.part0[30] 
	,\sa_snapshot[1].r.part0[29] ,\sa_snapshot[1].r.part0[28] 
	,\sa_snapshot[1].r.part0[27] ,\sa_snapshot[1].r.part0[26] 
	,\sa_snapshot[1].r.part0[25] ,\sa_snapshot[1].r.part0[24] 
	,\sa_snapshot[1].r.part0[23] ,\sa_snapshot[1].r.part0[22] 
	,\sa_snapshot[1].r.part0[21] ,\sa_snapshot[1].r.part0[20] 
	,\sa_snapshot[1].r.part0[19] ,\sa_snapshot[1].r.part0[18] 
	,\sa_snapshot[1].r.part0[17] ,\sa_snapshot[1].r.part0[16] 
	,\sa_snapshot[1].r.part0[15] ,\sa_snapshot[1].r.part0[14] 
	,\sa_snapshot[1].r.part0[13] ,\sa_snapshot[1].r.part0[12] 
	,\sa_snapshot[1].r.part0[11] ,\sa_snapshot[1].r.part0[10] 
	,\sa_snapshot[1].r.part0[9] ,\sa_snapshot[1].r.part0[8] 
	,\sa_snapshot[1].r.part0[7] ,\sa_snapshot[1].r.part0[6] 
	,\sa_snapshot[1].r.part0[5] ,\sa_snapshot[1].r.part0[4] 
	,\sa_snapshot[1].r.part0[3] ,\sa_snapshot[1].r.part0[2] 
	,\sa_snapshot[1].r.part0[1] ,\sa_snapshot[1].r.part0[0] 
	,\sa_snapshot[0].r.part1[31] ,\sa_snapshot[0].r.part1[30] 
	,\sa_snapshot[0].r.part1[29] ,\sa_snapshot[0].r.part1[28] 
	,\sa_snapshot[0].r.part1[27] ,\sa_snapshot[0].r.part1[26] 
	,\sa_snapshot[0].r.part1[25] ,\sa_snapshot[0].r.part1[24] 
	,\sa_snapshot[0].r.part1[23] ,\sa_snapshot[0].r.part1[22] 
	,\sa_snapshot[0].r.part1[21] ,\sa_snapshot[0].r.part1[20] 
	,\sa_snapshot[0].r.part1[19] ,\sa_snapshot[0].r.part1[18] 
	,\sa_snapshot[0].r.part1[17] ,\sa_snapshot[0].r.part1[16] 
	,\sa_snapshot[0].r.part1[15] ,\sa_snapshot[0].r.part1[14] 
	,\sa_snapshot[0].r.part1[13] ,\sa_snapshot[0].r.part1[12] 
	,\sa_snapshot[0].r.part1[11] ,\sa_snapshot[0].r.part1[10] 
	,\sa_snapshot[0].r.part1[9] ,\sa_snapshot[0].r.part1[8] 
	,\sa_snapshot[0].r.part1[7] ,\sa_snapshot[0].r.part1[6] 
	,\sa_snapshot[0].r.part1[5] ,\sa_snapshot[0].r.part1[4] 
	,\sa_snapshot[0].r.part1[3] ,\sa_snapshot[0].r.part1[2] 
	,\sa_snapshot[0].r.part1[1] ,\sa_snapshot[0].r.part1[0] 
	,\sa_snapshot[0].r.part0[31] ,\sa_snapshot[0].r.part0[30] 
	,\sa_snapshot[0].r.part0[29] ,\sa_snapshot[0].r.part0[28] 
	,\sa_snapshot[0].r.part0[27] ,\sa_snapshot[0].r.part0[26] 
	,\sa_snapshot[0].r.part0[25] ,\sa_snapshot[0].r.part0[24] 
	,\sa_snapshot[0].r.part0[23] ,\sa_snapshot[0].r.part0[22] 
	,\sa_snapshot[0].r.part0[21] ,\sa_snapshot[0].r.part0[20] 
	,\sa_snapshot[0].r.part0[19] ,\sa_snapshot[0].r.part0[18] 
	,\sa_snapshot[0].r.part0[17] ,\sa_snapshot[0].r.part0[16] 
	,\sa_snapshot[0].r.part0[15] ,\sa_snapshot[0].r.part0[14] 
	,\sa_snapshot[0].r.part0[13] ,\sa_snapshot[0].r.part0[12] 
	,\sa_snapshot[0].r.part0[11] ,\sa_snapshot[0].r.part0[10] 
	,\sa_snapshot[0].r.part0[9] ,\sa_snapshot[0].r.part0[8] 
	,\sa_snapshot[0].r.part0[7] ,\sa_snapshot[0].r.part0[6] 
	,\sa_snapshot[0].r.part0[5] ,\sa_snapshot[0].r.part0[4] 
	,\sa_snapshot[0].r.part0[3] ,\sa_snapshot[0].r.part0[2] 
	,\sa_snapshot[0].r.part0[1] ,\sa_snapshot[0].r.part0[0] ;
input \sa_count[31].r.part1[31] ,\sa_count[31].r.part1[30] 
	,\sa_count[31].r.part1[29] ,\sa_count[31].r.part1[28] 
	,\sa_count[31].r.part1[27] ,\sa_count[31].r.part1[26] 
	,\sa_count[31].r.part1[25] ,\sa_count[31].r.part1[24] 
	,\sa_count[31].r.part1[23] ,\sa_count[31].r.part1[22] 
	,\sa_count[31].r.part1[21] ,\sa_count[31].r.part1[20] 
	,\sa_count[31].r.part1[19] ,\sa_count[31].r.part1[18] 
	,\sa_count[31].r.part1[17] ,\sa_count[31].r.part1[16] 
	,\sa_count[31].r.part1[15] ,\sa_count[31].r.part1[14] 
	,\sa_count[31].r.part1[13] ,\sa_count[31].r.part1[12] 
	,\sa_count[31].r.part1[11] ,\sa_count[31].r.part1[10] 
	,\sa_count[31].r.part1[9] ,\sa_count[31].r.part1[8] 
	,\sa_count[31].r.part1[7] ,\sa_count[31].r.part1[6] 
	,\sa_count[31].r.part1[5] ,\sa_count[31].r.part1[4] 
	,\sa_count[31].r.part1[3] ,\sa_count[31].r.part1[2] 
	,\sa_count[31].r.part1[1] ,\sa_count[31].r.part1[0] 
	,\sa_count[31].r.part0[31] ,\sa_count[31].r.part0[30] 
	,\sa_count[31].r.part0[29] ,\sa_count[31].r.part0[28] 
	,\sa_count[31].r.part0[27] ,\sa_count[31].r.part0[26] 
	,\sa_count[31].r.part0[25] ,\sa_count[31].r.part0[24] 
	,\sa_count[31].r.part0[23] ,\sa_count[31].r.part0[22] 
	,\sa_count[31].r.part0[21] ,\sa_count[31].r.part0[20] 
	,\sa_count[31].r.part0[19] ,\sa_count[31].r.part0[18] 
	,\sa_count[31].r.part0[17] ,\sa_count[31].r.part0[16] 
	,\sa_count[31].r.part0[15] ,\sa_count[31].r.part0[14] 
	,\sa_count[31].r.part0[13] ,\sa_count[31].r.part0[12] 
	,\sa_count[31].r.part0[11] ,\sa_count[31].r.part0[10] 
	,\sa_count[31].r.part0[9] ,\sa_count[31].r.part0[8] 
	,\sa_count[31].r.part0[7] ,\sa_count[31].r.part0[6] 
	,\sa_count[31].r.part0[5] ,\sa_count[31].r.part0[4] 
	,\sa_count[31].r.part0[3] ,\sa_count[31].r.part0[2] 
	,\sa_count[31].r.part0[1] ,\sa_count[31].r.part0[0] 
	,\sa_count[30].r.part1[31] ,\sa_count[30].r.part1[30] 
	,\sa_count[30].r.part1[29] ,\sa_count[30].r.part1[28] 
	,\sa_count[30].r.part1[27] ,\sa_count[30].r.part1[26] 
	,\sa_count[30].r.part1[25] ,\sa_count[30].r.part1[24] 
	,\sa_count[30].r.part1[23] ,\sa_count[30].r.part1[22] 
	,\sa_count[30].r.part1[21] ,\sa_count[30].r.part1[20] 
	,\sa_count[30].r.part1[19] ,\sa_count[30].r.part1[18] 
	,\sa_count[30].r.part1[17] ,\sa_count[30].r.part1[16] 
	,\sa_count[30].r.part1[15] ,\sa_count[30].r.part1[14] 
	,\sa_count[30].r.part1[13] ,\sa_count[30].r.part1[12] 
	,\sa_count[30].r.part1[11] ,\sa_count[30].r.part1[10] 
	,\sa_count[30].r.part1[9] ,\sa_count[30].r.part1[8] 
	,\sa_count[30].r.part1[7] ,\sa_count[30].r.part1[6] 
	,\sa_count[30].r.part1[5] ,\sa_count[30].r.part1[4] 
	,\sa_count[30].r.part1[3] ,\sa_count[30].r.part1[2] 
	,\sa_count[30].r.part1[1] ,\sa_count[30].r.part1[0] 
	,\sa_count[30].r.part0[31] ,\sa_count[30].r.part0[30] 
	,\sa_count[30].r.part0[29] ,\sa_count[30].r.part0[28] 
	,\sa_count[30].r.part0[27] ,\sa_count[30].r.part0[26] 
	,\sa_count[30].r.part0[25] ,\sa_count[30].r.part0[24] 
	,\sa_count[30].r.part0[23] ,\sa_count[30].r.part0[22] 
	,\sa_count[30].r.part0[21] ,\sa_count[30].r.part0[20] 
	,\sa_count[30].r.part0[19] ,\sa_count[30].r.part0[18] 
	,\sa_count[30].r.part0[17] ,\sa_count[30].r.part0[16] 
	,\sa_count[30].r.part0[15] ,\sa_count[30].r.part0[14] 
	,\sa_count[30].r.part0[13] ,\sa_count[30].r.part0[12] 
	,\sa_count[30].r.part0[11] ,\sa_count[30].r.part0[10] 
	,\sa_count[30].r.part0[9] ,\sa_count[30].r.part0[8] 
	,\sa_count[30].r.part0[7] ,\sa_count[30].r.part0[6] 
	,\sa_count[30].r.part0[5] ,\sa_count[30].r.part0[4] 
	,\sa_count[30].r.part0[3] ,\sa_count[30].r.part0[2] 
	,\sa_count[30].r.part0[1] ,\sa_count[30].r.part0[0] 
	,\sa_count[29].r.part1[31] ,\sa_count[29].r.part1[30] 
	,\sa_count[29].r.part1[29] ,\sa_count[29].r.part1[28] 
	,\sa_count[29].r.part1[27] ,\sa_count[29].r.part1[26] 
	,\sa_count[29].r.part1[25] ,\sa_count[29].r.part1[24] 
	,\sa_count[29].r.part1[23] ,\sa_count[29].r.part1[22] 
	,\sa_count[29].r.part1[21] ,\sa_count[29].r.part1[20] 
	,\sa_count[29].r.part1[19] ,\sa_count[29].r.part1[18] 
	,\sa_count[29].r.part1[17] ,\sa_count[29].r.part1[16] 
	,\sa_count[29].r.part1[15] ,\sa_count[29].r.part1[14] 
	,\sa_count[29].r.part1[13] ,\sa_count[29].r.part1[12] 
	,\sa_count[29].r.part1[11] ,\sa_count[29].r.part1[10] 
	,\sa_count[29].r.part1[9] ,\sa_count[29].r.part1[8] 
	,\sa_count[29].r.part1[7] ,\sa_count[29].r.part1[6] 
	,\sa_count[29].r.part1[5] ,\sa_count[29].r.part1[4] 
	,\sa_count[29].r.part1[3] ,\sa_count[29].r.part1[2] 
	,\sa_count[29].r.part1[1] ,\sa_count[29].r.part1[0] 
	,\sa_count[29].r.part0[31] ,\sa_count[29].r.part0[30] 
	,\sa_count[29].r.part0[29] ,\sa_count[29].r.part0[28] 
	,\sa_count[29].r.part0[27] ,\sa_count[29].r.part0[26] 
	,\sa_count[29].r.part0[25] ,\sa_count[29].r.part0[24] 
	,\sa_count[29].r.part0[23] ,\sa_count[29].r.part0[22] 
	,\sa_count[29].r.part0[21] ,\sa_count[29].r.part0[20] 
	,\sa_count[29].r.part0[19] ,\sa_count[29].r.part0[18] 
	,\sa_count[29].r.part0[17] ,\sa_count[29].r.part0[16] 
	,\sa_count[29].r.part0[15] ,\sa_count[29].r.part0[14] 
	,\sa_count[29].r.part0[13] ,\sa_count[29].r.part0[12] 
	,\sa_count[29].r.part0[11] ,\sa_count[29].r.part0[10] 
	,\sa_count[29].r.part0[9] ,\sa_count[29].r.part0[8] 
	,\sa_count[29].r.part0[7] ,\sa_count[29].r.part0[6] 
	,\sa_count[29].r.part0[5] ,\sa_count[29].r.part0[4] 
	,\sa_count[29].r.part0[3] ,\sa_count[29].r.part0[2] 
	,\sa_count[29].r.part0[1] ,\sa_count[29].r.part0[0] 
	,\sa_count[28].r.part1[31] ,\sa_count[28].r.part1[30] 
	,\sa_count[28].r.part1[29] ,\sa_count[28].r.part1[28] 
	,\sa_count[28].r.part1[27] ,\sa_count[28].r.part1[26] 
	,\sa_count[28].r.part1[25] ,\sa_count[28].r.part1[24] 
	,\sa_count[28].r.part1[23] ,\sa_count[28].r.part1[22] 
	,\sa_count[28].r.part1[21] ,\sa_count[28].r.part1[20] 
	,\sa_count[28].r.part1[19] ,\sa_count[28].r.part1[18] 
	,\sa_count[28].r.part1[17] ,\sa_count[28].r.part1[16] 
	,\sa_count[28].r.part1[15] ,\sa_count[28].r.part1[14] 
	,\sa_count[28].r.part1[13] ,\sa_count[28].r.part1[12] 
	,\sa_count[28].r.part1[11] ,\sa_count[28].r.part1[10] 
	,\sa_count[28].r.part1[9] ,\sa_count[28].r.part1[8] 
	,\sa_count[28].r.part1[7] ,\sa_count[28].r.part1[6] 
	,\sa_count[28].r.part1[5] ,\sa_count[28].r.part1[4] 
	,\sa_count[28].r.part1[3] ,\sa_count[28].r.part1[2] 
	,\sa_count[28].r.part1[1] ,\sa_count[28].r.part1[0] 
	,\sa_count[28].r.part0[31] ,\sa_count[28].r.part0[30] 
	,\sa_count[28].r.part0[29] ,\sa_count[28].r.part0[28] 
	,\sa_count[28].r.part0[27] ,\sa_count[28].r.part0[26] 
	,\sa_count[28].r.part0[25] ,\sa_count[28].r.part0[24] 
	,\sa_count[28].r.part0[23] ,\sa_count[28].r.part0[22] 
	,\sa_count[28].r.part0[21] ,\sa_count[28].r.part0[20] 
	,\sa_count[28].r.part0[19] ,\sa_count[28].r.part0[18] 
	,\sa_count[28].r.part0[17] ,\sa_count[28].r.part0[16] 
	,\sa_count[28].r.part0[15] ,\sa_count[28].r.part0[14] 
	,\sa_count[28].r.part0[13] ,\sa_count[28].r.part0[12] 
	,\sa_count[28].r.part0[11] ,\sa_count[28].r.part0[10] 
	,\sa_count[28].r.part0[9] ,\sa_count[28].r.part0[8] 
	,\sa_count[28].r.part0[7] ,\sa_count[28].r.part0[6] 
	,\sa_count[28].r.part0[5] ,\sa_count[28].r.part0[4] 
	,\sa_count[28].r.part0[3] ,\sa_count[28].r.part0[2] 
	,\sa_count[28].r.part0[1] ,\sa_count[28].r.part0[0] 
	,\sa_count[27].r.part1[31] ,\sa_count[27].r.part1[30] 
	,\sa_count[27].r.part1[29] ,\sa_count[27].r.part1[28] 
	,\sa_count[27].r.part1[27] ,\sa_count[27].r.part1[26] 
	,\sa_count[27].r.part1[25] ,\sa_count[27].r.part1[24] 
	,\sa_count[27].r.part1[23] ,\sa_count[27].r.part1[22] 
	,\sa_count[27].r.part1[21] ,\sa_count[27].r.part1[20] 
	,\sa_count[27].r.part1[19] ,\sa_count[27].r.part1[18] 
	,\sa_count[27].r.part1[17] ,\sa_count[27].r.part1[16] 
	,\sa_count[27].r.part1[15] ,\sa_count[27].r.part1[14] 
	,\sa_count[27].r.part1[13] ,\sa_count[27].r.part1[12] 
	,\sa_count[27].r.part1[11] ,\sa_count[27].r.part1[10] 
	,\sa_count[27].r.part1[9] ,\sa_count[27].r.part1[8] 
	,\sa_count[27].r.part1[7] ,\sa_count[27].r.part1[6] 
	,\sa_count[27].r.part1[5] ,\sa_count[27].r.part1[4] 
	,\sa_count[27].r.part1[3] ,\sa_count[27].r.part1[2] 
	,\sa_count[27].r.part1[1] ,\sa_count[27].r.part1[0] 
	,\sa_count[27].r.part0[31] ,\sa_count[27].r.part0[30] 
	,\sa_count[27].r.part0[29] ,\sa_count[27].r.part0[28] 
	,\sa_count[27].r.part0[27] ,\sa_count[27].r.part0[26] 
	,\sa_count[27].r.part0[25] ,\sa_count[27].r.part0[24] 
	,\sa_count[27].r.part0[23] ,\sa_count[27].r.part0[22] 
	,\sa_count[27].r.part0[21] ,\sa_count[27].r.part0[20] 
	,\sa_count[27].r.part0[19] ,\sa_count[27].r.part0[18] 
	,\sa_count[27].r.part0[17] ,\sa_count[27].r.part0[16] 
	,\sa_count[27].r.part0[15] ,\sa_count[27].r.part0[14] 
	,\sa_count[27].r.part0[13] ,\sa_count[27].r.part0[12] 
	,\sa_count[27].r.part0[11] ,\sa_count[27].r.part0[10] 
	,\sa_count[27].r.part0[9] ,\sa_count[27].r.part0[8] 
	,\sa_count[27].r.part0[7] ,\sa_count[27].r.part0[6] 
	,\sa_count[27].r.part0[5] ,\sa_count[27].r.part0[4] 
	,\sa_count[27].r.part0[3] ,\sa_count[27].r.part0[2] 
	,\sa_count[27].r.part0[1] ,\sa_count[27].r.part0[0] 
	,\sa_count[26].r.part1[31] ,\sa_count[26].r.part1[30] 
	,\sa_count[26].r.part1[29] ,\sa_count[26].r.part1[28] 
	,\sa_count[26].r.part1[27] ,\sa_count[26].r.part1[26] 
	,\sa_count[26].r.part1[25] ,\sa_count[26].r.part1[24] 
	,\sa_count[26].r.part1[23] ,\sa_count[26].r.part1[22] 
	,\sa_count[26].r.part1[21] ,\sa_count[26].r.part1[20] 
	,\sa_count[26].r.part1[19] ,\sa_count[26].r.part1[18] 
	,\sa_count[26].r.part1[17] ,\sa_count[26].r.part1[16] 
	,\sa_count[26].r.part1[15] ,\sa_count[26].r.part1[14] 
	,\sa_count[26].r.part1[13] ,\sa_count[26].r.part1[12] 
	,\sa_count[26].r.part1[11] ,\sa_count[26].r.part1[10] 
	,\sa_count[26].r.part1[9] ,\sa_count[26].r.part1[8] 
	,\sa_count[26].r.part1[7] ,\sa_count[26].r.part1[6] 
	,\sa_count[26].r.part1[5] ,\sa_count[26].r.part1[4] 
	,\sa_count[26].r.part1[3] ,\sa_count[26].r.part1[2] 
	,\sa_count[26].r.part1[1] ,\sa_count[26].r.part1[0] 
	,\sa_count[26].r.part0[31] ,\sa_count[26].r.part0[30] 
	,\sa_count[26].r.part0[29] ,\sa_count[26].r.part0[28] 
	,\sa_count[26].r.part0[27] ,\sa_count[26].r.part0[26] 
	,\sa_count[26].r.part0[25] ,\sa_count[26].r.part0[24] 
	,\sa_count[26].r.part0[23] ,\sa_count[26].r.part0[22] 
	,\sa_count[26].r.part0[21] ,\sa_count[26].r.part0[20] 
	,\sa_count[26].r.part0[19] ,\sa_count[26].r.part0[18] 
	,\sa_count[26].r.part0[17] ,\sa_count[26].r.part0[16] 
	,\sa_count[26].r.part0[15] ,\sa_count[26].r.part0[14] 
	,\sa_count[26].r.part0[13] ,\sa_count[26].r.part0[12] 
	,\sa_count[26].r.part0[11] ,\sa_count[26].r.part0[10] 
	,\sa_count[26].r.part0[9] ,\sa_count[26].r.part0[8] 
	,\sa_count[26].r.part0[7] ,\sa_count[26].r.part0[6] 
	,\sa_count[26].r.part0[5] ,\sa_count[26].r.part0[4] 
	,\sa_count[26].r.part0[3] ,\sa_count[26].r.part0[2] 
	,\sa_count[26].r.part0[1] ,\sa_count[26].r.part0[0] 
	,\sa_count[25].r.part1[31] ,\sa_count[25].r.part1[30] 
	,\sa_count[25].r.part1[29] ,\sa_count[25].r.part1[28] 
	,\sa_count[25].r.part1[27] ,\sa_count[25].r.part1[26] 
	,\sa_count[25].r.part1[25] ,\sa_count[25].r.part1[24] 
	,\sa_count[25].r.part1[23] ,\sa_count[25].r.part1[22] 
	,\sa_count[25].r.part1[21] ,\sa_count[25].r.part1[20] 
	,\sa_count[25].r.part1[19] ,\sa_count[25].r.part1[18] 
	,\sa_count[25].r.part1[17] ,\sa_count[25].r.part1[16] 
	,\sa_count[25].r.part1[15] ,\sa_count[25].r.part1[14] 
	,\sa_count[25].r.part1[13] ,\sa_count[25].r.part1[12] 
	,\sa_count[25].r.part1[11] ,\sa_count[25].r.part1[10] 
	,\sa_count[25].r.part1[9] ,\sa_count[25].r.part1[8] 
	,\sa_count[25].r.part1[7] ,\sa_count[25].r.part1[6] 
	,\sa_count[25].r.part1[5] ,\sa_count[25].r.part1[4] 
	,\sa_count[25].r.part1[3] ,\sa_count[25].r.part1[2] 
	,\sa_count[25].r.part1[1] ,\sa_count[25].r.part1[0] 
	,\sa_count[25].r.part0[31] ,\sa_count[25].r.part0[30] 
	,\sa_count[25].r.part0[29] ,\sa_count[25].r.part0[28] 
	,\sa_count[25].r.part0[27] ,\sa_count[25].r.part0[26] 
	,\sa_count[25].r.part0[25] ,\sa_count[25].r.part0[24] 
	,\sa_count[25].r.part0[23] ,\sa_count[25].r.part0[22] 
	,\sa_count[25].r.part0[21] ,\sa_count[25].r.part0[20] 
	,\sa_count[25].r.part0[19] ,\sa_count[25].r.part0[18] 
	,\sa_count[25].r.part0[17] ,\sa_count[25].r.part0[16] 
	,\sa_count[25].r.part0[15] ,\sa_count[25].r.part0[14] 
	,\sa_count[25].r.part0[13] ,\sa_count[25].r.part0[12] 
	,\sa_count[25].r.part0[11] ,\sa_count[25].r.part0[10] 
	,\sa_count[25].r.part0[9] ,\sa_count[25].r.part0[8] 
	,\sa_count[25].r.part0[7] ,\sa_count[25].r.part0[6] 
	,\sa_count[25].r.part0[5] ,\sa_count[25].r.part0[4] 
	,\sa_count[25].r.part0[3] ,\sa_count[25].r.part0[2] 
	,\sa_count[25].r.part0[1] ,\sa_count[25].r.part0[0] 
	,\sa_count[24].r.part1[31] ,\sa_count[24].r.part1[30] 
	,\sa_count[24].r.part1[29] ,\sa_count[24].r.part1[28] 
	,\sa_count[24].r.part1[27] ,\sa_count[24].r.part1[26] 
	,\sa_count[24].r.part1[25] ,\sa_count[24].r.part1[24] 
	,\sa_count[24].r.part1[23] ,\sa_count[24].r.part1[22] 
	,\sa_count[24].r.part1[21] ,\sa_count[24].r.part1[20] 
	,\sa_count[24].r.part1[19] ,\sa_count[24].r.part1[18] 
	,\sa_count[24].r.part1[17] ,\sa_count[24].r.part1[16] 
	,\sa_count[24].r.part1[15] ,\sa_count[24].r.part1[14] 
	,\sa_count[24].r.part1[13] ,\sa_count[24].r.part1[12] 
	,\sa_count[24].r.part1[11] ,\sa_count[24].r.part1[10] 
	,\sa_count[24].r.part1[9] ,\sa_count[24].r.part1[8] 
	,\sa_count[24].r.part1[7] ,\sa_count[24].r.part1[6] 
	,\sa_count[24].r.part1[5] ,\sa_count[24].r.part1[4] 
	,\sa_count[24].r.part1[3] ,\sa_count[24].r.part1[2] 
	,\sa_count[24].r.part1[1] ,\sa_count[24].r.part1[0] 
	,\sa_count[24].r.part0[31] ,\sa_count[24].r.part0[30] 
	,\sa_count[24].r.part0[29] ,\sa_count[24].r.part0[28] 
	,\sa_count[24].r.part0[27] ,\sa_count[24].r.part0[26] 
	,\sa_count[24].r.part0[25] ,\sa_count[24].r.part0[24] 
	,\sa_count[24].r.part0[23] ,\sa_count[24].r.part0[22] 
	,\sa_count[24].r.part0[21] ,\sa_count[24].r.part0[20] 
	,\sa_count[24].r.part0[19] ,\sa_count[24].r.part0[18] 
	,\sa_count[24].r.part0[17] ,\sa_count[24].r.part0[16] 
	,\sa_count[24].r.part0[15] ,\sa_count[24].r.part0[14] 
	,\sa_count[24].r.part0[13] ,\sa_count[24].r.part0[12] 
	,\sa_count[24].r.part0[11] ,\sa_count[24].r.part0[10] 
	,\sa_count[24].r.part0[9] ,\sa_count[24].r.part0[8] 
	,\sa_count[24].r.part0[7] ,\sa_count[24].r.part0[6] 
	,\sa_count[24].r.part0[5] ,\sa_count[24].r.part0[4] 
	,\sa_count[24].r.part0[3] ,\sa_count[24].r.part0[2] 
	,\sa_count[24].r.part0[1] ,\sa_count[24].r.part0[0] 
	,\sa_count[23].r.part1[31] ,\sa_count[23].r.part1[30] 
	,\sa_count[23].r.part1[29] ,\sa_count[23].r.part1[28] 
	,\sa_count[23].r.part1[27] ,\sa_count[23].r.part1[26] 
	,\sa_count[23].r.part1[25] ,\sa_count[23].r.part1[24] 
	,\sa_count[23].r.part1[23] ,\sa_count[23].r.part1[22] 
	,\sa_count[23].r.part1[21] ,\sa_count[23].r.part1[20] 
	,\sa_count[23].r.part1[19] ,\sa_count[23].r.part1[18] 
	,\sa_count[23].r.part1[17] ,\sa_count[23].r.part1[16] 
	,\sa_count[23].r.part1[15] ,\sa_count[23].r.part1[14] 
	,\sa_count[23].r.part1[13] ,\sa_count[23].r.part1[12] 
	,\sa_count[23].r.part1[11] ,\sa_count[23].r.part1[10] 
	,\sa_count[23].r.part1[9] ,\sa_count[23].r.part1[8] 
	,\sa_count[23].r.part1[7] ,\sa_count[23].r.part1[6] 
	,\sa_count[23].r.part1[5] ,\sa_count[23].r.part1[4] 
	,\sa_count[23].r.part1[3] ,\sa_count[23].r.part1[2] 
	,\sa_count[23].r.part1[1] ,\sa_count[23].r.part1[0] 
	,\sa_count[23].r.part0[31] ,\sa_count[23].r.part0[30] 
	,\sa_count[23].r.part0[29] ,\sa_count[23].r.part0[28] 
	,\sa_count[23].r.part0[27] ,\sa_count[23].r.part0[26] 
	,\sa_count[23].r.part0[25] ,\sa_count[23].r.part0[24] 
	,\sa_count[23].r.part0[23] ,\sa_count[23].r.part0[22] 
	,\sa_count[23].r.part0[21] ,\sa_count[23].r.part0[20] 
	,\sa_count[23].r.part0[19] ,\sa_count[23].r.part0[18] 
	,\sa_count[23].r.part0[17] ,\sa_count[23].r.part0[16] 
	,\sa_count[23].r.part0[15] ,\sa_count[23].r.part0[14] 
	,\sa_count[23].r.part0[13] ,\sa_count[23].r.part0[12] 
	,\sa_count[23].r.part0[11] ,\sa_count[23].r.part0[10] 
	,\sa_count[23].r.part0[9] ,\sa_count[23].r.part0[8] 
	,\sa_count[23].r.part0[7] ,\sa_count[23].r.part0[6] 
	,\sa_count[23].r.part0[5] ,\sa_count[23].r.part0[4] 
	,\sa_count[23].r.part0[3] ,\sa_count[23].r.part0[2] 
	,\sa_count[23].r.part0[1] ,\sa_count[23].r.part0[0] 
	,\sa_count[22].r.part1[31] ,\sa_count[22].r.part1[30] 
	,\sa_count[22].r.part1[29] ,\sa_count[22].r.part1[28] 
	,\sa_count[22].r.part1[27] ,\sa_count[22].r.part1[26] 
	,\sa_count[22].r.part1[25] ,\sa_count[22].r.part1[24] 
	,\sa_count[22].r.part1[23] ,\sa_count[22].r.part1[22] 
	,\sa_count[22].r.part1[21] ,\sa_count[22].r.part1[20] 
	,\sa_count[22].r.part1[19] ,\sa_count[22].r.part1[18] 
	,\sa_count[22].r.part1[17] ,\sa_count[22].r.part1[16] 
	,\sa_count[22].r.part1[15] ,\sa_count[22].r.part1[14] 
	,\sa_count[22].r.part1[13] ,\sa_count[22].r.part1[12] 
	,\sa_count[22].r.part1[11] ,\sa_count[22].r.part1[10] 
	,\sa_count[22].r.part1[9] ,\sa_count[22].r.part1[8] 
	,\sa_count[22].r.part1[7] ,\sa_count[22].r.part1[6] 
	,\sa_count[22].r.part1[5] ,\sa_count[22].r.part1[4] 
	,\sa_count[22].r.part1[3] ,\sa_count[22].r.part1[2] 
	,\sa_count[22].r.part1[1] ,\sa_count[22].r.part1[0] 
	,\sa_count[22].r.part0[31] ,\sa_count[22].r.part0[30] 
	,\sa_count[22].r.part0[29] ,\sa_count[22].r.part0[28] 
	,\sa_count[22].r.part0[27] ,\sa_count[22].r.part0[26] 
	,\sa_count[22].r.part0[25] ,\sa_count[22].r.part0[24] 
	,\sa_count[22].r.part0[23] ,\sa_count[22].r.part0[22] 
	,\sa_count[22].r.part0[21] ,\sa_count[22].r.part0[20] 
	,\sa_count[22].r.part0[19] ,\sa_count[22].r.part0[18] 
	,\sa_count[22].r.part0[17] ,\sa_count[22].r.part0[16] 
	,\sa_count[22].r.part0[15] ,\sa_count[22].r.part0[14] 
	,\sa_count[22].r.part0[13] ,\sa_count[22].r.part0[12] 
	,\sa_count[22].r.part0[11] ,\sa_count[22].r.part0[10] 
	,\sa_count[22].r.part0[9] ,\sa_count[22].r.part0[8] 
	,\sa_count[22].r.part0[7] ,\sa_count[22].r.part0[6] 
	,\sa_count[22].r.part0[5] ,\sa_count[22].r.part0[4] 
	,\sa_count[22].r.part0[3] ,\sa_count[22].r.part0[2] 
	,\sa_count[22].r.part0[1] ,\sa_count[22].r.part0[0] 
	,\sa_count[21].r.part1[31] ,\sa_count[21].r.part1[30] 
	,\sa_count[21].r.part1[29] ,\sa_count[21].r.part1[28] 
	,\sa_count[21].r.part1[27] ,\sa_count[21].r.part1[26] 
	,\sa_count[21].r.part1[25] ,\sa_count[21].r.part1[24] 
	,\sa_count[21].r.part1[23] ,\sa_count[21].r.part1[22] 
	,\sa_count[21].r.part1[21] ,\sa_count[21].r.part1[20] 
	,\sa_count[21].r.part1[19] ,\sa_count[21].r.part1[18] 
	,\sa_count[21].r.part1[17] ,\sa_count[21].r.part1[16] 
	,\sa_count[21].r.part1[15] ,\sa_count[21].r.part1[14] 
	,\sa_count[21].r.part1[13] ,\sa_count[21].r.part1[12] 
	,\sa_count[21].r.part1[11] ,\sa_count[21].r.part1[10] 
	,\sa_count[21].r.part1[9] ,\sa_count[21].r.part1[8] 
	,\sa_count[21].r.part1[7] ,\sa_count[21].r.part1[6] 
	,\sa_count[21].r.part1[5] ,\sa_count[21].r.part1[4] 
	,\sa_count[21].r.part1[3] ,\sa_count[21].r.part1[2] 
	,\sa_count[21].r.part1[1] ,\sa_count[21].r.part1[0] 
	,\sa_count[21].r.part0[31] ,\sa_count[21].r.part0[30] 
	,\sa_count[21].r.part0[29] ,\sa_count[21].r.part0[28] 
	,\sa_count[21].r.part0[27] ,\sa_count[21].r.part0[26] 
	,\sa_count[21].r.part0[25] ,\sa_count[21].r.part0[24] 
	,\sa_count[21].r.part0[23] ,\sa_count[21].r.part0[22] 
	,\sa_count[21].r.part0[21] ,\sa_count[21].r.part0[20] 
	,\sa_count[21].r.part0[19] ,\sa_count[21].r.part0[18] 
	,\sa_count[21].r.part0[17] ,\sa_count[21].r.part0[16] 
	,\sa_count[21].r.part0[15] ,\sa_count[21].r.part0[14] 
	,\sa_count[21].r.part0[13] ,\sa_count[21].r.part0[12] 
	,\sa_count[21].r.part0[11] ,\sa_count[21].r.part0[10] 
	,\sa_count[21].r.part0[9] ,\sa_count[21].r.part0[8] 
	,\sa_count[21].r.part0[7] ,\sa_count[21].r.part0[6] 
	,\sa_count[21].r.part0[5] ,\sa_count[21].r.part0[4] 
	,\sa_count[21].r.part0[3] ,\sa_count[21].r.part0[2] 
	,\sa_count[21].r.part0[1] ,\sa_count[21].r.part0[0] 
	,\sa_count[20].r.part1[31] ,\sa_count[20].r.part1[30] 
	,\sa_count[20].r.part1[29] ,\sa_count[20].r.part1[28] 
	,\sa_count[20].r.part1[27] ,\sa_count[20].r.part1[26] 
	,\sa_count[20].r.part1[25] ,\sa_count[20].r.part1[24] 
	,\sa_count[20].r.part1[23] ,\sa_count[20].r.part1[22] 
	,\sa_count[20].r.part1[21] ,\sa_count[20].r.part1[20] 
	,\sa_count[20].r.part1[19] ,\sa_count[20].r.part1[18] 
	,\sa_count[20].r.part1[17] ,\sa_count[20].r.part1[16] 
	,\sa_count[20].r.part1[15] ,\sa_count[20].r.part1[14] 
	,\sa_count[20].r.part1[13] ,\sa_count[20].r.part1[12] 
	,\sa_count[20].r.part1[11] ,\sa_count[20].r.part1[10] 
	,\sa_count[20].r.part1[9] ,\sa_count[20].r.part1[8] 
	,\sa_count[20].r.part1[7] ,\sa_count[20].r.part1[6] 
	,\sa_count[20].r.part1[5] ,\sa_count[20].r.part1[4] 
	,\sa_count[20].r.part1[3] ,\sa_count[20].r.part1[2] 
	,\sa_count[20].r.part1[1] ,\sa_count[20].r.part1[0] 
	,\sa_count[20].r.part0[31] ,\sa_count[20].r.part0[30] 
	,\sa_count[20].r.part0[29] ,\sa_count[20].r.part0[28] 
	,\sa_count[20].r.part0[27] ,\sa_count[20].r.part0[26] 
	,\sa_count[20].r.part0[25] ,\sa_count[20].r.part0[24] 
	,\sa_count[20].r.part0[23] ,\sa_count[20].r.part0[22] 
	,\sa_count[20].r.part0[21] ,\sa_count[20].r.part0[20] 
	,\sa_count[20].r.part0[19] ,\sa_count[20].r.part0[18] 
	,\sa_count[20].r.part0[17] ,\sa_count[20].r.part0[16] 
	,\sa_count[20].r.part0[15] ,\sa_count[20].r.part0[14] 
	,\sa_count[20].r.part0[13] ,\sa_count[20].r.part0[12] 
	,\sa_count[20].r.part0[11] ,\sa_count[20].r.part0[10] 
	,\sa_count[20].r.part0[9] ,\sa_count[20].r.part0[8] 
	,\sa_count[20].r.part0[7] ,\sa_count[20].r.part0[6] 
	,\sa_count[20].r.part0[5] ,\sa_count[20].r.part0[4] 
	,\sa_count[20].r.part0[3] ,\sa_count[20].r.part0[2] 
	,\sa_count[20].r.part0[1] ,\sa_count[20].r.part0[0] 
	,\sa_count[19].r.part1[31] ,\sa_count[19].r.part1[30] 
	,\sa_count[19].r.part1[29] ,\sa_count[19].r.part1[28] 
	,\sa_count[19].r.part1[27] ,\sa_count[19].r.part1[26] 
	,\sa_count[19].r.part1[25] ,\sa_count[19].r.part1[24] 
	,\sa_count[19].r.part1[23] ,\sa_count[19].r.part1[22] 
	,\sa_count[19].r.part1[21] ,\sa_count[19].r.part1[20] 
	,\sa_count[19].r.part1[19] ,\sa_count[19].r.part1[18] 
	,\sa_count[19].r.part1[17] ,\sa_count[19].r.part1[16] 
	,\sa_count[19].r.part1[15] ,\sa_count[19].r.part1[14] 
	,\sa_count[19].r.part1[13] ,\sa_count[19].r.part1[12] 
	,\sa_count[19].r.part1[11] ,\sa_count[19].r.part1[10] 
	,\sa_count[19].r.part1[9] ,\sa_count[19].r.part1[8] 
	,\sa_count[19].r.part1[7] ,\sa_count[19].r.part1[6] 
	,\sa_count[19].r.part1[5] ,\sa_count[19].r.part1[4] 
	,\sa_count[19].r.part1[3] ,\sa_count[19].r.part1[2] 
	,\sa_count[19].r.part1[1] ,\sa_count[19].r.part1[0] 
	,\sa_count[19].r.part0[31] ,\sa_count[19].r.part0[30] 
	,\sa_count[19].r.part0[29] ,\sa_count[19].r.part0[28] 
	,\sa_count[19].r.part0[27] ,\sa_count[19].r.part0[26] 
	,\sa_count[19].r.part0[25] ,\sa_count[19].r.part0[24] 
	,\sa_count[19].r.part0[23] ,\sa_count[19].r.part0[22] 
	,\sa_count[19].r.part0[21] ,\sa_count[19].r.part0[20] 
	,\sa_count[19].r.part0[19] ,\sa_count[19].r.part0[18] 
	,\sa_count[19].r.part0[17] ,\sa_count[19].r.part0[16] 
	,\sa_count[19].r.part0[15] ,\sa_count[19].r.part0[14] 
	,\sa_count[19].r.part0[13] ,\sa_count[19].r.part0[12] 
	,\sa_count[19].r.part0[11] ,\sa_count[19].r.part0[10] 
	,\sa_count[19].r.part0[9] ,\sa_count[19].r.part0[8] 
	,\sa_count[19].r.part0[7] ,\sa_count[19].r.part0[6] 
	,\sa_count[19].r.part0[5] ,\sa_count[19].r.part0[4] 
	,\sa_count[19].r.part0[3] ,\sa_count[19].r.part0[2] 
	,\sa_count[19].r.part0[1] ,\sa_count[19].r.part0[0] 
	,\sa_count[18].r.part1[31] ,\sa_count[18].r.part1[30] 
	,\sa_count[18].r.part1[29] ,\sa_count[18].r.part1[28] 
	,\sa_count[18].r.part1[27] ,\sa_count[18].r.part1[26] 
	,\sa_count[18].r.part1[25] ,\sa_count[18].r.part1[24] 
	,\sa_count[18].r.part1[23] ,\sa_count[18].r.part1[22] 
	,\sa_count[18].r.part1[21] ,\sa_count[18].r.part1[20] 
	,\sa_count[18].r.part1[19] ,\sa_count[18].r.part1[18] 
	,\sa_count[18].r.part1[17] ,\sa_count[18].r.part1[16] 
	,\sa_count[18].r.part1[15] ,\sa_count[18].r.part1[14] 
	,\sa_count[18].r.part1[13] ,\sa_count[18].r.part1[12] 
	,\sa_count[18].r.part1[11] ,\sa_count[18].r.part1[10] 
	,\sa_count[18].r.part1[9] ,\sa_count[18].r.part1[8] 
	,\sa_count[18].r.part1[7] ,\sa_count[18].r.part1[6] 
	,\sa_count[18].r.part1[5] ,\sa_count[18].r.part1[4] 
	,\sa_count[18].r.part1[3] ,\sa_count[18].r.part1[2] 
	,\sa_count[18].r.part1[1] ,\sa_count[18].r.part1[0] 
	,\sa_count[18].r.part0[31] ,\sa_count[18].r.part0[30] 
	,\sa_count[18].r.part0[29] ,\sa_count[18].r.part0[28] 
	,\sa_count[18].r.part0[27] ,\sa_count[18].r.part0[26] 
	,\sa_count[18].r.part0[25] ,\sa_count[18].r.part0[24] 
	,\sa_count[18].r.part0[23] ,\sa_count[18].r.part0[22] 
	,\sa_count[18].r.part0[21] ,\sa_count[18].r.part0[20] 
	,\sa_count[18].r.part0[19] ,\sa_count[18].r.part0[18] 
	,\sa_count[18].r.part0[17] ,\sa_count[18].r.part0[16] 
	,\sa_count[18].r.part0[15] ,\sa_count[18].r.part0[14] 
	,\sa_count[18].r.part0[13] ,\sa_count[18].r.part0[12] 
	,\sa_count[18].r.part0[11] ,\sa_count[18].r.part0[10] 
	,\sa_count[18].r.part0[9] ,\sa_count[18].r.part0[8] 
	,\sa_count[18].r.part0[7] ,\sa_count[18].r.part0[6] 
	,\sa_count[18].r.part0[5] ,\sa_count[18].r.part0[4] 
	,\sa_count[18].r.part0[3] ,\sa_count[18].r.part0[2] 
	,\sa_count[18].r.part0[1] ,\sa_count[18].r.part0[0] 
	,\sa_count[17].r.part1[31] ,\sa_count[17].r.part1[30] 
	,\sa_count[17].r.part1[29] ,\sa_count[17].r.part1[28] 
	,\sa_count[17].r.part1[27] ,\sa_count[17].r.part1[26] 
	,\sa_count[17].r.part1[25] ,\sa_count[17].r.part1[24] 
	,\sa_count[17].r.part1[23] ,\sa_count[17].r.part1[22] 
	,\sa_count[17].r.part1[21] ,\sa_count[17].r.part1[20] 
	,\sa_count[17].r.part1[19] ,\sa_count[17].r.part1[18] 
	,\sa_count[17].r.part1[17] ,\sa_count[17].r.part1[16] 
	,\sa_count[17].r.part1[15] ,\sa_count[17].r.part1[14] 
	,\sa_count[17].r.part1[13] ,\sa_count[17].r.part1[12] 
	,\sa_count[17].r.part1[11] ,\sa_count[17].r.part1[10] 
	,\sa_count[17].r.part1[9] ,\sa_count[17].r.part1[8] 
	,\sa_count[17].r.part1[7] ,\sa_count[17].r.part1[6] 
	,\sa_count[17].r.part1[5] ,\sa_count[17].r.part1[4] 
	,\sa_count[17].r.part1[3] ,\sa_count[17].r.part1[2] 
	,\sa_count[17].r.part1[1] ,\sa_count[17].r.part1[0] 
	,\sa_count[17].r.part0[31] ,\sa_count[17].r.part0[30] 
	,\sa_count[17].r.part0[29] ,\sa_count[17].r.part0[28] 
	,\sa_count[17].r.part0[27] ,\sa_count[17].r.part0[26] 
	,\sa_count[17].r.part0[25] ,\sa_count[17].r.part0[24] 
	,\sa_count[17].r.part0[23] ,\sa_count[17].r.part0[22] 
	,\sa_count[17].r.part0[21] ,\sa_count[17].r.part0[20] 
	,\sa_count[17].r.part0[19] ,\sa_count[17].r.part0[18] 
	,\sa_count[17].r.part0[17] ,\sa_count[17].r.part0[16] 
	,\sa_count[17].r.part0[15] ,\sa_count[17].r.part0[14] 
	,\sa_count[17].r.part0[13] ,\sa_count[17].r.part0[12] 
	,\sa_count[17].r.part0[11] ,\sa_count[17].r.part0[10] 
	,\sa_count[17].r.part0[9] ,\sa_count[17].r.part0[8] 
	,\sa_count[17].r.part0[7] ,\sa_count[17].r.part0[6] 
	,\sa_count[17].r.part0[5] ,\sa_count[17].r.part0[4] 
	,\sa_count[17].r.part0[3] ,\sa_count[17].r.part0[2] 
	,\sa_count[17].r.part0[1] ,\sa_count[17].r.part0[0] 
	,\sa_count[16].r.part1[31] ,\sa_count[16].r.part1[30] 
	,\sa_count[16].r.part1[29] ,\sa_count[16].r.part1[28] 
	,\sa_count[16].r.part1[27] ,\sa_count[16].r.part1[26] 
	,\sa_count[16].r.part1[25] ,\sa_count[16].r.part1[24] 
	,\sa_count[16].r.part1[23] ,\sa_count[16].r.part1[22] 
	,\sa_count[16].r.part1[21] ,\sa_count[16].r.part1[20] 
	,\sa_count[16].r.part1[19] ,\sa_count[16].r.part1[18] 
	,\sa_count[16].r.part1[17] ,\sa_count[16].r.part1[16] 
	,\sa_count[16].r.part1[15] ,\sa_count[16].r.part1[14] 
	,\sa_count[16].r.part1[13] ,\sa_count[16].r.part1[12] 
	,\sa_count[16].r.part1[11] ,\sa_count[16].r.part1[10] 
	,\sa_count[16].r.part1[9] ,\sa_count[16].r.part1[8] 
	,\sa_count[16].r.part1[7] ,\sa_count[16].r.part1[6] 
	,\sa_count[16].r.part1[5] ,\sa_count[16].r.part1[4] 
	,\sa_count[16].r.part1[3] ,\sa_count[16].r.part1[2] 
	,\sa_count[16].r.part1[1] ,\sa_count[16].r.part1[0] 
	,\sa_count[16].r.part0[31] ,\sa_count[16].r.part0[30] 
	,\sa_count[16].r.part0[29] ,\sa_count[16].r.part0[28] 
	,\sa_count[16].r.part0[27] ,\sa_count[16].r.part0[26] 
	,\sa_count[16].r.part0[25] ,\sa_count[16].r.part0[24] 
	,\sa_count[16].r.part0[23] ,\sa_count[16].r.part0[22] 
	,\sa_count[16].r.part0[21] ,\sa_count[16].r.part0[20] 
	,\sa_count[16].r.part0[19] ,\sa_count[16].r.part0[18] 
	,\sa_count[16].r.part0[17] ,\sa_count[16].r.part0[16] 
	,\sa_count[16].r.part0[15] ,\sa_count[16].r.part0[14] 
	,\sa_count[16].r.part0[13] ,\sa_count[16].r.part0[12] 
	,\sa_count[16].r.part0[11] ,\sa_count[16].r.part0[10] 
	,\sa_count[16].r.part0[9] ,\sa_count[16].r.part0[8] 
	,\sa_count[16].r.part0[7] ,\sa_count[16].r.part0[6] 
	,\sa_count[16].r.part0[5] ,\sa_count[16].r.part0[4] 
	,\sa_count[16].r.part0[3] ,\sa_count[16].r.part0[2] 
	,\sa_count[16].r.part0[1] ,\sa_count[16].r.part0[0] 
	,\sa_count[15].r.part1[31] ,\sa_count[15].r.part1[30] 
	,\sa_count[15].r.part1[29] ,\sa_count[15].r.part1[28] 
	,\sa_count[15].r.part1[27] ,\sa_count[15].r.part1[26] 
	,\sa_count[15].r.part1[25] ,\sa_count[15].r.part1[24] 
	,\sa_count[15].r.part1[23] ,\sa_count[15].r.part1[22] 
	,\sa_count[15].r.part1[21] ,\sa_count[15].r.part1[20] 
	,\sa_count[15].r.part1[19] ,\sa_count[15].r.part1[18] 
	,\sa_count[15].r.part1[17] ,\sa_count[15].r.part1[16] 
	,\sa_count[15].r.part1[15] ,\sa_count[15].r.part1[14] 
	,\sa_count[15].r.part1[13] ,\sa_count[15].r.part1[12] 
	,\sa_count[15].r.part1[11] ,\sa_count[15].r.part1[10] 
	,\sa_count[15].r.part1[9] ,\sa_count[15].r.part1[8] 
	,\sa_count[15].r.part1[7] ,\sa_count[15].r.part1[6] 
	,\sa_count[15].r.part1[5] ,\sa_count[15].r.part1[4] 
	,\sa_count[15].r.part1[3] ,\sa_count[15].r.part1[2] 
	,\sa_count[15].r.part1[1] ,\sa_count[15].r.part1[0] 
	,\sa_count[15].r.part0[31] ,\sa_count[15].r.part0[30] 
	,\sa_count[15].r.part0[29] ,\sa_count[15].r.part0[28] 
	,\sa_count[15].r.part0[27] ,\sa_count[15].r.part0[26] 
	,\sa_count[15].r.part0[25] ,\sa_count[15].r.part0[24] 
	,\sa_count[15].r.part0[23] ,\sa_count[15].r.part0[22] 
	,\sa_count[15].r.part0[21] ,\sa_count[15].r.part0[20] 
	,\sa_count[15].r.part0[19] ,\sa_count[15].r.part0[18] 
	,\sa_count[15].r.part0[17] ,\sa_count[15].r.part0[16] 
	,\sa_count[15].r.part0[15] ,\sa_count[15].r.part0[14] 
	,\sa_count[15].r.part0[13] ,\sa_count[15].r.part0[12] 
	,\sa_count[15].r.part0[11] ,\sa_count[15].r.part0[10] 
	,\sa_count[15].r.part0[9] ,\sa_count[15].r.part0[8] 
	,\sa_count[15].r.part0[7] ,\sa_count[15].r.part0[6] 
	,\sa_count[15].r.part0[5] ,\sa_count[15].r.part0[4] 
	,\sa_count[15].r.part0[3] ,\sa_count[15].r.part0[2] 
	,\sa_count[15].r.part0[1] ,\sa_count[15].r.part0[0] 
	,\sa_count[14].r.part1[31] ,\sa_count[14].r.part1[30] 
	,\sa_count[14].r.part1[29] ,\sa_count[14].r.part1[28] 
	,\sa_count[14].r.part1[27] ,\sa_count[14].r.part1[26] 
	,\sa_count[14].r.part1[25] ,\sa_count[14].r.part1[24] 
	,\sa_count[14].r.part1[23] ,\sa_count[14].r.part1[22] 
	,\sa_count[14].r.part1[21] ,\sa_count[14].r.part1[20] 
	,\sa_count[14].r.part1[19] ,\sa_count[14].r.part1[18] 
	,\sa_count[14].r.part1[17] ,\sa_count[14].r.part1[16] 
	,\sa_count[14].r.part1[15] ,\sa_count[14].r.part1[14] 
	,\sa_count[14].r.part1[13] ,\sa_count[14].r.part1[12] 
	,\sa_count[14].r.part1[11] ,\sa_count[14].r.part1[10] 
	,\sa_count[14].r.part1[9] ,\sa_count[14].r.part1[8] 
	,\sa_count[14].r.part1[7] ,\sa_count[14].r.part1[6] 
	,\sa_count[14].r.part1[5] ,\sa_count[14].r.part1[4] 
	,\sa_count[14].r.part1[3] ,\sa_count[14].r.part1[2] 
	,\sa_count[14].r.part1[1] ,\sa_count[14].r.part1[0] 
	,\sa_count[14].r.part0[31] ,\sa_count[14].r.part0[30] 
	,\sa_count[14].r.part0[29] ,\sa_count[14].r.part0[28] 
	,\sa_count[14].r.part0[27] ,\sa_count[14].r.part0[26] 
	,\sa_count[14].r.part0[25] ,\sa_count[14].r.part0[24] 
	,\sa_count[14].r.part0[23] ,\sa_count[14].r.part0[22] 
	,\sa_count[14].r.part0[21] ,\sa_count[14].r.part0[20] 
	,\sa_count[14].r.part0[19] ,\sa_count[14].r.part0[18] 
	,\sa_count[14].r.part0[17] ,\sa_count[14].r.part0[16] 
	,\sa_count[14].r.part0[15] ,\sa_count[14].r.part0[14] 
	,\sa_count[14].r.part0[13] ,\sa_count[14].r.part0[12] 
	,\sa_count[14].r.part0[11] ,\sa_count[14].r.part0[10] 
	,\sa_count[14].r.part0[9] ,\sa_count[14].r.part0[8] 
	,\sa_count[14].r.part0[7] ,\sa_count[14].r.part0[6] 
	,\sa_count[14].r.part0[5] ,\sa_count[14].r.part0[4] 
	,\sa_count[14].r.part0[3] ,\sa_count[14].r.part0[2] 
	,\sa_count[14].r.part0[1] ,\sa_count[14].r.part0[0] 
	,\sa_count[13].r.part1[31] ,\sa_count[13].r.part1[30] 
	,\sa_count[13].r.part1[29] ,\sa_count[13].r.part1[28] 
	,\sa_count[13].r.part1[27] ,\sa_count[13].r.part1[26] 
	,\sa_count[13].r.part1[25] ,\sa_count[13].r.part1[24] 
	,\sa_count[13].r.part1[23] ,\sa_count[13].r.part1[22] 
	,\sa_count[13].r.part1[21] ,\sa_count[13].r.part1[20] 
	,\sa_count[13].r.part1[19] ,\sa_count[13].r.part1[18] 
	,\sa_count[13].r.part1[17] ,\sa_count[13].r.part1[16] 
	,\sa_count[13].r.part1[15] ,\sa_count[13].r.part1[14] 
	,\sa_count[13].r.part1[13] ,\sa_count[13].r.part1[12] 
	,\sa_count[13].r.part1[11] ,\sa_count[13].r.part1[10] 
	,\sa_count[13].r.part1[9] ,\sa_count[13].r.part1[8] 
	,\sa_count[13].r.part1[7] ,\sa_count[13].r.part1[6] 
	,\sa_count[13].r.part1[5] ,\sa_count[13].r.part1[4] 
	,\sa_count[13].r.part1[3] ,\sa_count[13].r.part1[2] 
	,\sa_count[13].r.part1[1] ,\sa_count[13].r.part1[0] 
	,\sa_count[13].r.part0[31] ,\sa_count[13].r.part0[30] 
	,\sa_count[13].r.part0[29] ,\sa_count[13].r.part0[28] 
	,\sa_count[13].r.part0[27] ,\sa_count[13].r.part0[26] 
	,\sa_count[13].r.part0[25] ,\sa_count[13].r.part0[24] 
	,\sa_count[13].r.part0[23] ,\sa_count[13].r.part0[22] 
	,\sa_count[13].r.part0[21] ,\sa_count[13].r.part0[20] 
	,\sa_count[13].r.part0[19] ,\sa_count[13].r.part0[18] 
	,\sa_count[13].r.part0[17] ,\sa_count[13].r.part0[16] 
	,\sa_count[13].r.part0[15] ,\sa_count[13].r.part0[14] 
	,\sa_count[13].r.part0[13] ,\sa_count[13].r.part0[12] 
	,\sa_count[13].r.part0[11] ,\sa_count[13].r.part0[10] 
	,\sa_count[13].r.part0[9] ,\sa_count[13].r.part0[8] 
	,\sa_count[13].r.part0[7] ,\sa_count[13].r.part0[6] 
	,\sa_count[13].r.part0[5] ,\sa_count[13].r.part0[4] 
	,\sa_count[13].r.part0[3] ,\sa_count[13].r.part0[2] 
	,\sa_count[13].r.part0[1] ,\sa_count[13].r.part0[0] 
	,\sa_count[12].r.part1[31] ,\sa_count[12].r.part1[30] 
	,\sa_count[12].r.part1[29] ,\sa_count[12].r.part1[28] 
	,\sa_count[12].r.part1[27] ,\sa_count[12].r.part1[26] 
	,\sa_count[12].r.part1[25] ,\sa_count[12].r.part1[24] 
	,\sa_count[12].r.part1[23] ,\sa_count[12].r.part1[22] 
	,\sa_count[12].r.part1[21] ,\sa_count[12].r.part1[20] 
	,\sa_count[12].r.part1[19] ,\sa_count[12].r.part1[18] 
	,\sa_count[12].r.part1[17] ,\sa_count[12].r.part1[16] 
	,\sa_count[12].r.part1[15] ,\sa_count[12].r.part1[14] 
	,\sa_count[12].r.part1[13] ,\sa_count[12].r.part1[12] 
	,\sa_count[12].r.part1[11] ,\sa_count[12].r.part1[10] 
	,\sa_count[12].r.part1[9] ,\sa_count[12].r.part1[8] 
	,\sa_count[12].r.part1[7] ,\sa_count[12].r.part1[6] 
	,\sa_count[12].r.part1[5] ,\sa_count[12].r.part1[4] 
	,\sa_count[12].r.part1[3] ,\sa_count[12].r.part1[2] 
	,\sa_count[12].r.part1[1] ,\sa_count[12].r.part1[0] 
	,\sa_count[12].r.part0[31] ,\sa_count[12].r.part0[30] 
	,\sa_count[12].r.part0[29] ,\sa_count[12].r.part0[28] 
	,\sa_count[12].r.part0[27] ,\sa_count[12].r.part0[26] 
	,\sa_count[12].r.part0[25] ,\sa_count[12].r.part0[24] 
	,\sa_count[12].r.part0[23] ,\sa_count[12].r.part0[22] 
	,\sa_count[12].r.part0[21] ,\sa_count[12].r.part0[20] 
	,\sa_count[12].r.part0[19] ,\sa_count[12].r.part0[18] 
	,\sa_count[12].r.part0[17] ,\sa_count[12].r.part0[16] 
	,\sa_count[12].r.part0[15] ,\sa_count[12].r.part0[14] 
	,\sa_count[12].r.part0[13] ,\sa_count[12].r.part0[12] 
	,\sa_count[12].r.part0[11] ,\sa_count[12].r.part0[10] 
	,\sa_count[12].r.part0[9] ,\sa_count[12].r.part0[8] 
	,\sa_count[12].r.part0[7] ,\sa_count[12].r.part0[6] 
	,\sa_count[12].r.part0[5] ,\sa_count[12].r.part0[4] 
	,\sa_count[12].r.part0[3] ,\sa_count[12].r.part0[2] 
	,\sa_count[12].r.part0[1] ,\sa_count[12].r.part0[0] 
	,\sa_count[11].r.part1[31] ,\sa_count[11].r.part1[30] 
	,\sa_count[11].r.part1[29] ,\sa_count[11].r.part1[28] 
	,\sa_count[11].r.part1[27] ,\sa_count[11].r.part1[26] 
	,\sa_count[11].r.part1[25] ,\sa_count[11].r.part1[24] 
	,\sa_count[11].r.part1[23] ,\sa_count[11].r.part1[22] 
	,\sa_count[11].r.part1[21] ,\sa_count[11].r.part1[20] 
	,\sa_count[11].r.part1[19] ,\sa_count[11].r.part1[18] 
	,\sa_count[11].r.part1[17] ,\sa_count[11].r.part1[16] 
	,\sa_count[11].r.part1[15] ,\sa_count[11].r.part1[14] 
	,\sa_count[11].r.part1[13] ,\sa_count[11].r.part1[12] 
	,\sa_count[11].r.part1[11] ,\sa_count[11].r.part1[10] 
	,\sa_count[11].r.part1[9] ,\sa_count[11].r.part1[8] 
	,\sa_count[11].r.part1[7] ,\sa_count[11].r.part1[6] 
	,\sa_count[11].r.part1[5] ,\sa_count[11].r.part1[4] 
	,\sa_count[11].r.part1[3] ,\sa_count[11].r.part1[2] 
	,\sa_count[11].r.part1[1] ,\sa_count[11].r.part1[0] 
	,\sa_count[11].r.part0[31] ,\sa_count[11].r.part0[30] 
	,\sa_count[11].r.part0[29] ,\sa_count[11].r.part0[28] 
	,\sa_count[11].r.part0[27] ,\sa_count[11].r.part0[26] 
	,\sa_count[11].r.part0[25] ,\sa_count[11].r.part0[24] 
	,\sa_count[11].r.part0[23] ,\sa_count[11].r.part0[22] 
	,\sa_count[11].r.part0[21] ,\sa_count[11].r.part0[20] 
	,\sa_count[11].r.part0[19] ,\sa_count[11].r.part0[18] 
	,\sa_count[11].r.part0[17] ,\sa_count[11].r.part0[16] 
	,\sa_count[11].r.part0[15] ,\sa_count[11].r.part0[14] 
	,\sa_count[11].r.part0[13] ,\sa_count[11].r.part0[12] 
	,\sa_count[11].r.part0[11] ,\sa_count[11].r.part0[10] 
	,\sa_count[11].r.part0[9] ,\sa_count[11].r.part0[8] 
	,\sa_count[11].r.part0[7] ,\sa_count[11].r.part0[6] 
	,\sa_count[11].r.part0[5] ,\sa_count[11].r.part0[4] 
	,\sa_count[11].r.part0[3] ,\sa_count[11].r.part0[2] 
	,\sa_count[11].r.part0[1] ,\sa_count[11].r.part0[0] 
	,\sa_count[10].r.part1[31] ,\sa_count[10].r.part1[30] 
	,\sa_count[10].r.part1[29] ,\sa_count[10].r.part1[28] 
	,\sa_count[10].r.part1[27] ,\sa_count[10].r.part1[26] 
	,\sa_count[10].r.part1[25] ,\sa_count[10].r.part1[24] 
	,\sa_count[10].r.part1[23] ,\sa_count[10].r.part1[22] 
	,\sa_count[10].r.part1[21] ,\sa_count[10].r.part1[20] 
	,\sa_count[10].r.part1[19] ,\sa_count[10].r.part1[18] 
	,\sa_count[10].r.part1[17] ,\sa_count[10].r.part1[16] 
	,\sa_count[10].r.part1[15] ,\sa_count[10].r.part1[14] 
	,\sa_count[10].r.part1[13] ,\sa_count[10].r.part1[12] 
	,\sa_count[10].r.part1[11] ,\sa_count[10].r.part1[10] 
	,\sa_count[10].r.part1[9] ,\sa_count[10].r.part1[8] 
	,\sa_count[10].r.part1[7] ,\sa_count[10].r.part1[6] 
	,\sa_count[10].r.part1[5] ,\sa_count[10].r.part1[4] 
	,\sa_count[10].r.part1[3] ,\sa_count[10].r.part1[2] 
	,\sa_count[10].r.part1[1] ,\sa_count[10].r.part1[0] 
	,\sa_count[10].r.part0[31] ,\sa_count[10].r.part0[30] 
	,\sa_count[10].r.part0[29] ,\sa_count[10].r.part0[28] 
	,\sa_count[10].r.part0[27] ,\sa_count[10].r.part0[26] 
	,\sa_count[10].r.part0[25] ,\sa_count[10].r.part0[24] 
	,\sa_count[10].r.part0[23] ,\sa_count[10].r.part0[22] 
	,\sa_count[10].r.part0[21] ,\sa_count[10].r.part0[20] 
	,\sa_count[10].r.part0[19] ,\sa_count[10].r.part0[18] 
	,\sa_count[10].r.part0[17] ,\sa_count[10].r.part0[16] 
	,\sa_count[10].r.part0[15] ,\sa_count[10].r.part0[14] 
	,\sa_count[10].r.part0[13] ,\sa_count[10].r.part0[12] 
	,\sa_count[10].r.part0[11] ,\sa_count[10].r.part0[10] 
	,\sa_count[10].r.part0[9] ,\sa_count[10].r.part0[8] 
	,\sa_count[10].r.part0[7] ,\sa_count[10].r.part0[6] 
	,\sa_count[10].r.part0[5] ,\sa_count[10].r.part0[4] 
	,\sa_count[10].r.part0[3] ,\sa_count[10].r.part0[2] 
	,\sa_count[10].r.part0[1] ,\sa_count[10].r.part0[0] 
	,\sa_count[9].r.part1[31] ,\sa_count[9].r.part1[30] 
	,\sa_count[9].r.part1[29] ,\sa_count[9].r.part1[28] 
	,\sa_count[9].r.part1[27] ,\sa_count[9].r.part1[26] 
	,\sa_count[9].r.part1[25] ,\sa_count[9].r.part1[24] 
	,\sa_count[9].r.part1[23] ,\sa_count[9].r.part1[22] 
	,\sa_count[9].r.part1[21] ,\sa_count[9].r.part1[20] 
	,\sa_count[9].r.part1[19] ,\sa_count[9].r.part1[18] 
	,\sa_count[9].r.part1[17] ,\sa_count[9].r.part1[16] 
	,\sa_count[9].r.part1[15] ,\sa_count[9].r.part1[14] 
	,\sa_count[9].r.part1[13] ,\sa_count[9].r.part1[12] 
	,\sa_count[9].r.part1[11] ,\sa_count[9].r.part1[10] 
	,\sa_count[9].r.part1[9] ,\sa_count[9].r.part1[8] 
	,\sa_count[9].r.part1[7] ,\sa_count[9].r.part1[6] 
	,\sa_count[9].r.part1[5] ,\sa_count[9].r.part1[4] 
	,\sa_count[9].r.part1[3] ,\sa_count[9].r.part1[2] 
	,\sa_count[9].r.part1[1] ,\sa_count[9].r.part1[0] 
	,\sa_count[9].r.part0[31] ,\sa_count[9].r.part0[30] 
	,\sa_count[9].r.part0[29] ,\sa_count[9].r.part0[28] 
	,\sa_count[9].r.part0[27] ,\sa_count[9].r.part0[26] 
	,\sa_count[9].r.part0[25] ,\sa_count[9].r.part0[24] 
	,\sa_count[9].r.part0[23] ,\sa_count[9].r.part0[22] 
	,\sa_count[9].r.part0[21] ,\sa_count[9].r.part0[20] 
	,\sa_count[9].r.part0[19] ,\sa_count[9].r.part0[18] 
	,\sa_count[9].r.part0[17] ,\sa_count[9].r.part0[16] 
	,\sa_count[9].r.part0[15] ,\sa_count[9].r.part0[14] 
	,\sa_count[9].r.part0[13] ,\sa_count[9].r.part0[12] 
	,\sa_count[9].r.part0[11] ,\sa_count[9].r.part0[10] 
	,\sa_count[9].r.part0[9] ,\sa_count[9].r.part0[8] 
	,\sa_count[9].r.part0[7] ,\sa_count[9].r.part0[6] 
	,\sa_count[9].r.part0[5] ,\sa_count[9].r.part0[4] 
	,\sa_count[9].r.part0[3] ,\sa_count[9].r.part0[2] 
	,\sa_count[9].r.part0[1] ,\sa_count[9].r.part0[0] 
	,\sa_count[8].r.part1[31] ,\sa_count[8].r.part1[30] 
	,\sa_count[8].r.part1[29] ,\sa_count[8].r.part1[28] 
	,\sa_count[8].r.part1[27] ,\sa_count[8].r.part1[26] 
	,\sa_count[8].r.part1[25] ,\sa_count[8].r.part1[24] 
	,\sa_count[8].r.part1[23] ,\sa_count[8].r.part1[22] 
	,\sa_count[8].r.part1[21] ,\sa_count[8].r.part1[20] 
	,\sa_count[8].r.part1[19] ,\sa_count[8].r.part1[18] 
	,\sa_count[8].r.part1[17] ,\sa_count[8].r.part1[16] 
	,\sa_count[8].r.part1[15] ,\sa_count[8].r.part1[14] 
	,\sa_count[8].r.part1[13] ,\sa_count[8].r.part1[12] 
	,\sa_count[8].r.part1[11] ,\sa_count[8].r.part1[10] 
	,\sa_count[8].r.part1[9] ,\sa_count[8].r.part1[8] 
	,\sa_count[8].r.part1[7] ,\sa_count[8].r.part1[6] 
	,\sa_count[8].r.part1[5] ,\sa_count[8].r.part1[4] 
	,\sa_count[8].r.part1[3] ,\sa_count[8].r.part1[2] 
	,\sa_count[8].r.part1[1] ,\sa_count[8].r.part1[0] 
	,\sa_count[8].r.part0[31] ,\sa_count[8].r.part0[30] 
	,\sa_count[8].r.part0[29] ,\sa_count[8].r.part0[28] 
	,\sa_count[8].r.part0[27] ,\sa_count[8].r.part0[26] 
	,\sa_count[8].r.part0[25] ,\sa_count[8].r.part0[24] 
	,\sa_count[8].r.part0[23] ,\sa_count[8].r.part0[22] 
	,\sa_count[8].r.part0[21] ,\sa_count[8].r.part0[20] 
	,\sa_count[8].r.part0[19] ,\sa_count[8].r.part0[18] 
	,\sa_count[8].r.part0[17] ,\sa_count[8].r.part0[16] 
	,\sa_count[8].r.part0[15] ,\sa_count[8].r.part0[14] 
	,\sa_count[8].r.part0[13] ,\sa_count[8].r.part0[12] 
	,\sa_count[8].r.part0[11] ,\sa_count[8].r.part0[10] 
	,\sa_count[8].r.part0[9] ,\sa_count[8].r.part0[8] 
	,\sa_count[8].r.part0[7] ,\sa_count[8].r.part0[6] 
	,\sa_count[8].r.part0[5] ,\sa_count[8].r.part0[4] 
	,\sa_count[8].r.part0[3] ,\sa_count[8].r.part0[2] 
	,\sa_count[8].r.part0[1] ,\sa_count[8].r.part0[0] 
	,\sa_count[7].r.part1[31] ,\sa_count[7].r.part1[30] 
	,\sa_count[7].r.part1[29] ,\sa_count[7].r.part1[28] 
	,\sa_count[7].r.part1[27] ,\sa_count[7].r.part1[26] 
	,\sa_count[7].r.part1[25] ,\sa_count[7].r.part1[24] 
	,\sa_count[7].r.part1[23] ,\sa_count[7].r.part1[22] 
	,\sa_count[7].r.part1[21] ,\sa_count[7].r.part1[20] 
	,\sa_count[7].r.part1[19] ,\sa_count[7].r.part1[18] 
	,\sa_count[7].r.part1[17] ,\sa_count[7].r.part1[16] 
	,\sa_count[7].r.part1[15] ,\sa_count[7].r.part1[14] 
	,\sa_count[7].r.part1[13] ,\sa_count[7].r.part1[12] 
	,\sa_count[7].r.part1[11] ,\sa_count[7].r.part1[10] 
	,\sa_count[7].r.part1[9] ,\sa_count[7].r.part1[8] 
	,\sa_count[7].r.part1[7] ,\sa_count[7].r.part1[6] 
	,\sa_count[7].r.part1[5] ,\sa_count[7].r.part1[4] 
	,\sa_count[7].r.part1[3] ,\sa_count[7].r.part1[2] 
	,\sa_count[7].r.part1[1] ,\sa_count[7].r.part1[0] 
	,\sa_count[7].r.part0[31] ,\sa_count[7].r.part0[30] 
	,\sa_count[7].r.part0[29] ,\sa_count[7].r.part0[28] 
	,\sa_count[7].r.part0[27] ,\sa_count[7].r.part0[26] 
	,\sa_count[7].r.part0[25] ,\sa_count[7].r.part0[24] 
	,\sa_count[7].r.part0[23] ,\sa_count[7].r.part0[22] 
	,\sa_count[7].r.part0[21] ,\sa_count[7].r.part0[20] 
	,\sa_count[7].r.part0[19] ,\sa_count[7].r.part0[18] 
	,\sa_count[7].r.part0[17] ,\sa_count[7].r.part0[16] 
	,\sa_count[7].r.part0[15] ,\sa_count[7].r.part0[14] 
	,\sa_count[7].r.part0[13] ,\sa_count[7].r.part0[12] 
	,\sa_count[7].r.part0[11] ,\sa_count[7].r.part0[10] 
	,\sa_count[7].r.part0[9] ,\sa_count[7].r.part0[8] 
	,\sa_count[7].r.part0[7] ,\sa_count[7].r.part0[6] 
	,\sa_count[7].r.part0[5] ,\sa_count[7].r.part0[4] 
	,\sa_count[7].r.part0[3] ,\sa_count[7].r.part0[2] 
	,\sa_count[7].r.part0[1] ,\sa_count[7].r.part0[0] 
	,\sa_count[6].r.part1[31] ,\sa_count[6].r.part1[30] 
	,\sa_count[6].r.part1[29] ,\sa_count[6].r.part1[28] 
	,\sa_count[6].r.part1[27] ,\sa_count[6].r.part1[26] 
	,\sa_count[6].r.part1[25] ,\sa_count[6].r.part1[24] 
	,\sa_count[6].r.part1[23] ,\sa_count[6].r.part1[22] 
	,\sa_count[6].r.part1[21] ,\sa_count[6].r.part1[20] 
	,\sa_count[6].r.part1[19] ,\sa_count[6].r.part1[18] 
	,\sa_count[6].r.part1[17] ,\sa_count[6].r.part1[16] 
	,\sa_count[6].r.part1[15] ,\sa_count[6].r.part1[14] 
	,\sa_count[6].r.part1[13] ,\sa_count[6].r.part1[12] 
	,\sa_count[6].r.part1[11] ,\sa_count[6].r.part1[10] 
	,\sa_count[6].r.part1[9] ,\sa_count[6].r.part1[8] 
	,\sa_count[6].r.part1[7] ,\sa_count[6].r.part1[6] 
	,\sa_count[6].r.part1[5] ,\sa_count[6].r.part1[4] 
	,\sa_count[6].r.part1[3] ,\sa_count[6].r.part1[2] 
	,\sa_count[6].r.part1[1] ,\sa_count[6].r.part1[0] 
	,\sa_count[6].r.part0[31] ,\sa_count[6].r.part0[30] 
	,\sa_count[6].r.part0[29] ,\sa_count[6].r.part0[28] 
	,\sa_count[6].r.part0[27] ,\sa_count[6].r.part0[26] 
	,\sa_count[6].r.part0[25] ,\sa_count[6].r.part0[24] 
	,\sa_count[6].r.part0[23] ,\sa_count[6].r.part0[22] 
	,\sa_count[6].r.part0[21] ,\sa_count[6].r.part0[20] 
	,\sa_count[6].r.part0[19] ,\sa_count[6].r.part0[18] 
	,\sa_count[6].r.part0[17] ,\sa_count[6].r.part0[16] 
	,\sa_count[6].r.part0[15] ,\sa_count[6].r.part0[14] 
	,\sa_count[6].r.part0[13] ,\sa_count[6].r.part0[12] 
	,\sa_count[6].r.part0[11] ,\sa_count[6].r.part0[10] 
	,\sa_count[6].r.part0[9] ,\sa_count[6].r.part0[8] 
	,\sa_count[6].r.part0[7] ,\sa_count[6].r.part0[6] 
	,\sa_count[6].r.part0[5] ,\sa_count[6].r.part0[4] 
	,\sa_count[6].r.part0[3] ,\sa_count[6].r.part0[2] 
	,\sa_count[6].r.part0[1] ,\sa_count[6].r.part0[0] 
	,\sa_count[5].r.part1[31] ,\sa_count[5].r.part1[30] 
	,\sa_count[5].r.part1[29] ,\sa_count[5].r.part1[28] 
	,\sa_count[5].r.part1[27] ,\sa_count[5].r.part1[26] 
	,\sa_count[5].r.part1[25] ,\sa_count[5].r.part1[24] 
	,\sa_count[5].r.part1[23] ,\sa_count[5].r.part1[22] 
	,\sa_count[5].r.part1[21] ,\sa_count[5].r.part1[20] 
	,\sa_count[5].r.part1[19] ,\sa_count[5].r.part1[18] 
	,\sa_count[5].r.part1[17] ,\sa_count[5].r.part1[16] 
	,\sa_count[5].r.part1[15] ,\sa_count[5].r.part1[14] 
	,\sa_count[5].r.part1[13] ,\sa_count[5].r.part1[12] 
	,\sa_count[5].r.part1[11] ,\sa_count[5].r.part1[10] 
	,\sa_count[5].r.part1[9] ,\sa_count[5].r.part1[8] 
	,\sa_count[5].r.part1[7] ,\sa_count[5].r.part1[6] 
	,\sa_count[5].r.part1[5] ,\sa_count[5].r.part1[4] 
	,\sa_count[5].r.part1[3] ,\sa_count[5].r.part1[2] 
	,\sa_count[5].r.part1[1] ,\sa_count[5].r.part1[0] 
	,\sa_count[5].r.part0[31] ,\sa_count[5].r.part0[30] 
	,\sa_count[5].r.part0[29] ,\sa_count[5].r.part0[28] 
	,\sa_count[5].r.part0[27] ,\sa_count[5].r.part0[26] 
	,\sa_count[5].r.part0[25] ,\sa_count[5].r.part0[24] 
	,\sa_count[5].r.part0[23] ,\sa_count[5].r.part0[22] 
	,\sa_count[5].r.part0[21] ,\sa_count[5].r.part0[20] 
	,\sa_count[5].r.part0[19] ,\sa_count[5].r.part0[18] 
	,\sa_count[5].r.part0[17] ,\sa_count[5].r.part0[16] 
	,\sa_count[5].r.part0[15] ,\sa_count[5].r.part0[14] 
	,\sa_count[5].r.part0[13] ,\sa_count[5].r.part0[12] 
	,\sa_count[5].r.part0[11] ,\sa_count[5].r.part0[10] 
	,\sa_count[5].r.part0[9] ,\sa_count[5].r.part0[8] 
	,\sa_count[5].r.part0[7] ,\sa_count[5].r.part0[6] 
	,\sa_count[5].r.part0[5] ,\sa_count[5].r.part0[4] 
	,\sa_count[5].r.part0[3] ,\sa_count[5].r.part0[2] 
	,\sa_count[5].r.part0[1] ,\sa_count[5].r.part0[0] 
	,\sa_count[4].r.part1[31] ,\sa_count[4].r.part1[30] 
	,\sa_count[4].r.part1[29] ,\sa_count[4].r.part1[28] 
	,\sa_count[4].r.part1[27] ,\sa_count[4].r.part1[26] 
	,\sa_count[4].r.part1[25] ,\sa_count[4].r.part1[24] 
	,\sa_count[4].r.part1[23] ,\sa_count[4].r.part1[22] 
	,\sa_count[4].r.part1[21] ,\sa_count[4].r.part1[20] 
	,\sa_count[4].r.part1[19] ,\sa_count[4].r.part1[18] 
	,\sa_count[4].r.part1[17] ,\sa_count[4].r.part1[16] 
	,\sa_count[4].r.part1[15] ,\sa_count[4].r.part1[14] 
	,\sa_count[4].r.part1[13] ,\sa_count[4].r.part1[12] 
	,\sa_count[4].r.part1[11] ,\sa_count[4].r.part1[10] 
	,\sa_count[4].r.part1[9] ,\sa_count[4].r.part1[8] 
	,\sa_count[4].r.part1[7] ,\sa_count[4].r.part1[6] 
	,\sa_count[4].r.part1[5] ,\sa_count[4].r.part1[4] 
	,\sa_count[4].r.part1[3] ,\sa_count[4].r.part1[2] 
	,\sa_count[4].r.part1[1] ,\sa_count[4].r.part1[0] 
	,\sa_count[4].r.part0[31] ,\sa_count[4].r.part0[30] 
	,\sa_count[4].r.part0[29] ,\sa_count[4].r.part0[28] 
	,\sa_count[4].r.part0[27] ,\sa_count[4].r.part0[26] 
	,\sa_count[4].r.part0[25] ,\sa_count[4].r.part0[24] 
	,\sa_count[4].r.part0[23] ,\sa_count[4].r.part0[22] 
	,\sa_count[4].r.part0[21] ,\sa_count[4].r.part0[20] 
	,\sa_count[4].r.part0[19] ,\sa_count[4].r.part0[18] 
	,\sa_count[4].r.part0[17] ,\sa_count[4].r.part0[16] 
	,\sa_count[4].r.part0[15] ,\sa_count[4].r.part0[14] 
	,\sa_count[4].r.part0[13] ,\sa_count[4].r.part0[12] 
	,\sa_count[4].r.part0[11] ,\sa_count[4].r.part0[10] 
	,\sa_count[4].r.part0[9] ,\sa_count[4].r.part0[8] 
	,\sa_count[4].r.part0[7] ,\sa_count[4].r.part0[6] 
	,\sa_count[4].r.part0[5] ,\sa_count[4].r.part0[4] 
	,\sa_count[4].r.part0[3] ,\sa_count[4].r.part0[2] 
	,\sa_count[4].r.part0[1] ,\sa_count[4].r.part0[0] 
	,\sa_count[3].r.part1[31] ,\sa_count[3].r.part1[30] 
	,\sa_count[3].r.part1[29] ,\sa_count[3].r.part1[28] 
	,\sa_count[3].r.part1[27] ,\sa_count[3].r.part1[26] 
	,\sa_count[3].r.part1[25] ,\sa_count[3].r.part1[24] 
	,\sa_count[3].r.part1[23] ,\sa_count[3].r.part1[22] 
	,\sa_count[3].r.part1[21] ,\sa_count[3].r.part1[20] 
	,\sa_count[3].r.part1[19] ,\sa_count[3].r.part1[18] 
	,\sa_count[3].r.part1[17] ,\sa_count[3].r.part1[16] 
	,\sa_count[3].r.part1[15] ,\sa_count[3].r.part1[14] 
	,\sa_count[3].r.part1[13] ,\sa_count[3].r.part1[12] 
	,\sa_count[3].r.part1[11] ,\sa_count[3].r.part1[10] 
	,\sa_count[3].r.part1[9] ,\sa_count[3].r.part1[8] 
	,\sa_count[3].r.part1[7] ,\sa_count[3].r.part1[6] 
	,\sa_count[3].r.part1[5] ,\sa_count[3].r.part1[4] 
	,\sa_count[3].r.part1[3] ,\sa_count[3].r.part1[2] 
	,\sa_count[3].r.part1[1] ,\sa_count[3].r.part1[0] 
	,\sa_count[3].r.part0[31] ,\sa_count[3].r.part0[30] 
	,\sa_count[3].r.part0[29] ,\sa_count[3].r.part0[28] 
	,\sa_count[3].r.part0[27] ,\sa_count[3].r.part0[26] 
	,\sa_count[3].r.part0[25] ,\sa_count[3].r.part0[24] 
	,\sa_count[3].r.part0[23] ,\sa_count[3].r.part0[22] 
	,\sa_count[3].r.part0[21] ,\sa_count[3].r.part0[20] 
	,\sa_count[3].r.part0[19] ,\sa_count[3].r.part0[18] 
	,\sa_count[3].r.part0[17] ,\sa_count[3].r.part0[16] 
	,\sa_count[3].r.part0[15] ,\sa_count[3].r.part0[14] 
	,\sa_count[3].r.part0[13] ,\sa_count[3].r.part0[12] 
	,\sa_count[3].r.part0[11] ,\sa_count[3].r.part0[10] 
	,\sa_count[3].r.part0[9] ,\sa_count[3].r.part0[8] 
	,\sa_count[3].r.part0[7] ,\sa_count[3].r.part0[6] 
	,\sa_count[3].r.part0[5] ,\sa_count[3].r.part0[4] 
	,\sa_count[3].r.part0[3] ,\sa_count[3].r.part0[2] 
	,\sa_count[3].r.part0[1] ,\sa_count[3].r.part0[0] 
	,\sa_count[2].r.part1[31] ,\sa_count[2].r.part1[30] 
	,\sa_count[2].r.part1[29] ,\sa_count[2].r.part1[28] 
	,\sa_count[2].r.part1[27] ,\sa_count[2].r.part1[26] 
	,\sa_count[2].r.part1[25] ,\sa_count[2].r.part1[24] 
	,\sa_count[2].r.part1[23] ,\sa_count[2].r.part1[22] 
	,\sa_count[2].r.part1[21] ,\sa_count[2].r.part1[20] 
	,\sa_count[2].r.part1[19] ,\sa_count[2].r.part1[18] 
	,\sa_count[2].r.part1[17] ,\sa_count[2].r.part1[16] 
	,\sa_count[2].r.part1[15] ,\sa_count[2].r.part1[14] 
	,\sa_count[2].r.part1[13] ,\sa_count[2].r.part1[12] 
	,\sa_count[2].r.part1[11] ,\sa_count[2].r.part1[10] 
	,\sa_count[2].r.part1[9] ,\sa_count[2].r.part1[8] 
	,\sa_count[2].r.part1[7] ,\sa_count[2].r.part1[6] 
	,\sa_count[2].r.part1[5] ,\sa_count[2].r.part1[4] 
	,\sa_count[2].r.part1[3] ,\sa_count[2].r.part1[2] 
	,\sa_count[2].r.part1[1] ,\sa_count[2].r.part1[0] 
	,\sa_count[2].r.part0[31] ,\sa_count[2].r.part0[30] 
	,\sa_count[2].r.part0[29] ,\sa_count[2].r.part0[28] 
	,\sa_count[2].r.part0[27] ,\sa_count[2].r.part0[26] 
	,\sa_count[2].r.part0[25] ,\sa_count[2].r.part0[24] 
	,\sa_count[2].r.part0[23] ,\sa_count[2].r.part0[22] 
	,\sa_count[2].r.part0[21] ,\sa_count[2].r.part0[20] 
	,\sa_count[2].r.part0[19] ,\sa_count[2].r.part0[18] 
	,\sa_count[2].r.part0[17] ,\sa_count[2].r.part0[16] 
	,\sa_count[2].r.part0[15] ,\sa_count[2].r.part0[14] 
	,\sa_count[2].r.part0[13] ,\sa_count[2].r.part0[12] 
	,\sa_count[2].r.part0[11] ,\sa_count[2].r.part0[10] 
	,\sa_count[2].r.part0[9] ,\sa_count[2].r.part0[8] 
	,\sa_count[2].r.part0[7] ,\sa_count[2].r.part0[6] 
	,\sa_count[2].r.part0[5] ,\sa_count[2].r.part0[4] 
	,\sa_count[2].r.part0[3] ,\sa_count[2].r.part0[2] 
	,\sa_count[2].r.part0[1] ,\sa_count[2].r.part0[0] 
	,\sa_count[1].r.part1[31] ,\sa_count[1].r.part1[30] 
	,\sa_count[1].r.part1[29] ,\sa_count[1].r.part1[28] 
	,\sa_count[1].r.part1[27] ,\sa_count[1].r.part1[26] 
	,\sa_count[1].r.part1[25] ,\sa_count[1].r.part1[24] 
	,\sa_count[1].r.part1[23] ,\sa_count[1].r.part1[22] 
	,\sa_count[1].r.part1[21] ,\sa_count[1].r.part1[20] 
	,\sa_count[1].r.part1[19] ,\sa_count[1].r.part1[18] 
	,\sa_count[1].r.part1[17] ,\sa_count[1].r.part1[16] 
	,\sa_count[1].r.part1[15] ,\sa_count[1].r.part1[14] 
	,\sa_count[1].r.part1[13] ,\sa_count[1].r.part1[12] 
	,\sa_count[1].r.part1[11] ,\sa_count[1].r.part1[10] 
	,\sa_count[1].r.part1[9] ,\sa_count[1].r.part1[8] 
	,\sa_count[1].r.part1[7] ,\sa_count[1].r.part1[6] 
	,\sa_count[1].r.part1[5] ,\sa_count[1].r.part1[4] 
	,\sa_count[1].r.part1[3] ,\sa_count[1].r.part1[2] 
	,\sa_count[1].r.part1[1] ,\sa_count[1].r.part1[0] 
	,\sa_count[1].r.part0[31] ,\sa_count[1].r.part0[30] 
	,\sa_count[1].r.part0[29] ,\sa_count[1].r.part0[28] 
	,\sa_count[1].r.part0[27] ,\sa_count[1].r.part0[26] 
	,\sa_count[1].r.part0[25] ,\sa_count[1].r.part0[24] 
	,\sa_count[1].r.part0[23] ,\sa_count[1].r.part0[22] 
	,\sa_count[1].r.part0[21] ,\sa_count[1].r.part0[20] 
	,\sa_count[1].r.part0[19] ,\sa_count[1].r.part0[18] 
	,\sa_count[1].r.part0[17] ,\sa_count[1].r.part0[16] 
	,\sa_count[1].r.part0[15] ,\sa_count[1].r.part0[14] 
	,\sa_count[1].r.part0[13] ,\sa_count[1].r.part0[12] 
	,\sa_count[1].r.part0[11] ,\sa_count[1].r.part0[10] 
	,\sa_count[1].r.part0[9] ,\sa_count[1].r.part0[8] 
	,\sa_count[1].r.part0[7] ,\sa_count[1].r.part0[6] 
	,\sa_count[1].r.part0[5] ,\sa_count[1].r.part0[4] 
	,\sa_count[1].r.part0[3] ,\sa_count[1].r.part0[2] 
	,\sa_count[1].r.part0[1] ,\sa_count[1].r.part0[0] 
	,\sa_count[0].r.part1[31] ,\sa_count[0].r.part1[30] 
	,\sa_count[0].r.part1[29] ,\sa_count[0].r.part1[28] 
	,\sa_count[0].r.part1[27] ,\sa_count[0].r.part1[26] 
	,\sa_count[0].r.part1[25] ,\sa_count[0].r.part1[24] 
	,\sa_count[0].r.part1[23] ,\sa_count[0].r.part1[22] 
	,\sa_count[0].r.part1[21] ,\sa_count[0].r.part1[20] 
	,\sa_count[0].r.part1[19] ,\sa_count[0].r.part1[18] 
	,\sa_count[0].r.part1[17] ,\sa_count[0].r.part1[16] 
	,\sa_count[0].r.part1[15] ,\sa_count[0].r.part1[14] 
	,\sa_count[0].r.part1[13] ,\sa_count[0].r.part1[12] 
	,\sa_count[0].r.part1[11] ,\sa_count[0].r.part1[10] 
	,\sa_count[0].r.part1[9] ,\sa_count[0].r.part1[8] 
	,\sa_count[0].r.part1[7] ,\sa_count[0].r.part1[6] 
	,\sa_count[0].r.part1[5] ,\sa_count[0].r.part1[4] 
	,\sa_count[0].r.part1[3] ,\sa_count[0].r.part1[2] 
	,\sa_count[0].r.part1[1] ,\sa_count[0].r.part1[0] 
	,\sa_count[0].r.part0[31] ,\sa_count[0].r.part0[30] 
	,\sa_count[0].r.part0[29] ,\sa_count[0].r.part0[28] 
	,\sa_count[0].r.part0[27] ,\sa_count[0].r.part0[26] 
	,\sa_count[0].r.part0[25] ,\sa_count[0].r.part0[24] 
	,\sa_count[0].r.part0[23] ,\sa_count[0].r.part0[22] 
	,\sa_count[0].r.part0[21] ,\sa_count[0].r.part0[20] 
	,\sa_count[0].r.part0[19] ,\sa_count[0].r.part0[18] 
	,\sa_count[0].r.part0[17] ,\sa_count[0].r.part0[16] 
	,\sa_count[0].r.part0[15] ,\sa_count[0].r.part0[14] 
	,\sa_count[0].r.part0[13] ,\sa_count[0].r.part0[12] 
	,\sa_count[0].r.part0[11] ,\sa_count[0].r.part0[10] 
	,\sa_count[0].r.part0[9] ,\sa_count[0].r.part0[8] 
	,\sa_count[0].r.part0[7] ,\sa_count[0].r.part0[6] 
	,\sa_count[0].r.part0[5] ,\sa_count[0].r.part0[4] 
	,\sa_count[0].r.part0[3] ,\sa_count[0].r.part0[2] 
	,\sa_count[0].r.part0[1] ,\sa_count[0].r.part0[0] ;
input debug_kme_ib_tready;
wire [0:83] _zy_simnet_rbus_ring_o_0_w$;
wire [0:82] _zy_simnet_kme_cceip0_ob_out_1_w$;
wire _zy_simnet_kme_cceip0_ob_in_mod_2_w$;
wire [0:82] _zy_simnet_kme_cceip1_ob_out_3_w$;
wire _zy_simnet_kme_cceip1_ob_in_mod_4_w$;
wire [0:82] _zy_simnet_kme_cceip2_ob_out_5_w$;
wire _zy_simnet_kme_cceip2_ob_in_mod_6_w$;
wire [0:82] _zy_simnet_kme_cceip3_ob_out_7_w$;
wire _zy_simnet_kme_cceip3_ob_in_mod_8_w$;
wire [0:82] _zy_simnet_kme_cddip0_ob_out_9_w$;
wire _zy_simnet_kme_cddip0_ob_in_mod_10_w$;
wire [0:82] _zy_simnet_kme_cddip1_ob_out_11_w$;
wire _zy_simnet_kme_cddip1_ob_in_mod_12_w$;
wire [0:82] _zy_simnet_kme_cddip2_ob_out_13_w$;
wire _zy_simnet_kme_cddip2_ob_in_mod_14_w$;
wire [0:82] _zy_simnet_kme_cddip3_ob_out_15_w$;
wire _zy_simnet_kme_cddip3_ob_in_mod_16_w$;
wire [0:37] _zy_simnet_kim_dout_17_w$;
wire [0:2175] _zy_simnet_labels_18_w$;
wire [0:8] _zy_simnet_tready_override_19_w$;
wire [0:6] _zy_simnet_cceip_encrypt_kop_fifo_override_20_w$;
wire [0:6] _zy_simnet_cceip_validate_kop_fifo_override_21_w$;
wire [0:6] _zy_simnet_cddip_decrypt_kop_fifo_override_22_w$;
wire [0:31] _zy_simnet_sa_global_ctrl_23_w$;
wire _zy_simnet_cio_24;
wire [0:10] _zy_simnet_locl_addr_25_w$;
wire _zy_simnet_locl_wr_strb_26_w$;
wire [0:31] _zy_simnet_locl_wr_data_27_w$;
wire _zy_simnet_locl_rd_strb_28_w$;
wire [0:31] _zy_simnet_locl_rd_data_29_w$;
wire _zy_simnet_locl_ack_30_w$;
wire _zy_simnet_locl_err_ack_31_w$;
wire [0:31] _zy_simnet_tvar_32;
wire [0:24] _zy_simnet_tvar_33;
wire _zy_simnet_tvar_34;
wire _zy_simnet_tvar_35;
wire _zy_simnet_tvar_36;
wire _zy_simnet_tvar_37;
wire [0:31] _zy_simnet_cceip0_out_ia_wdata_38_w$;
wire [0:31] _zy_simnet_cceip0_out_ia_wdata_39_w$;
wire [0:31] _zy_simnet_cceip0_out_ia_wdata_40_w$;
wire [0:12] _zy_simnet_cceip0_out_ia_config_41_w$;
wire [0:11] _zy_simnet_cceip0_out_im_config_42_w$;
wire [0:1] _zy_simnet_dio_43;
wire [0:31] _zy_simnet_cceip1_out_ia_wdata_44_w$;
wire [0:31] _zy_simnet_cceip1_out_ia_wdata_45_w$;
wire [0:31] _zy_simnet_cceip1_out_ia_wdata_46_w$;
wire [0:12] _zy_simnet_cceip1_out_ia_config_47_w$;
wire [0:11] _zy_simnet_cceip1_out_im_config_48_w$;
wire [0:1] _zy_simnet_dio_49;
wire [0:31] _zy_simnet_cceip2_out_ia_wdata_50_w$;
wire [0:31] _zy_simnet_cceip2_out_ia_wdata_51_w$;
wire [0:31] _zy_simnet_cceip2_out_ia_wdata_52_w$;
wire [0:12] _zy_simnet_cceip2_out_ia_config_53_w$;
wire [0:11] _zy_simnet_cceip2_out_im_config_54_w$;
wire [0:1] _zy_simnet_dio_55;
wire [0:31] _zy_simnet_cceip3_out_ia_wdata_56_w$;
wire [0:31] _zy_simnet_cceip3_out_ia_wdata_57_w$;
wire [0:31] _zy_simnet_cceip3_out_ia_wdata_58_w$;
wire [0:12] _zy_simnet_cceip3_out_ia_config_59_w$;
wire [0:11] _zy_simnet_cceip3_out_im_config_60_w$;
wire [0:1] _zy_simnet_dio_61;
wire [0:31] _zy_simnet_cddip0_out_ia_wdata_62_w$;
wire [0:31] _zy_simnet_cddip0_out_ia_wdata_63_w$;
wire [0:31] _zy_simnet_cddip0_out_ia_wdata_64_w$;
wire [0:12] _zy_simnet_cddip0_out_ia_config_65_w$;
wire [0:11] _zy_simnet_cddip0_out_im_config_66_w$;
wire [0:1] _zy_simnet_dio_67;
wire [0:31] _zy_simnet_cddip1_out_ia_wdata_68_w$;
wire [0:31] _zy_simnet_cddip1_out_ia_wdata_69_w$;
wire [0:31] _zy_simnet_cddip1_out_ia_wdata_70_w$;
wire [0:12] _zy_simnet_cddip1_out_ia_config_71_w$;
wire [0:11] _zy_simnet_cddip1_out_im_config_72_w$;
wire [0:1] _zy_simnet_dio_73;
wire [0:31] _zy_simnet_cddip2_out_ia_wdata_74_w$;
wire [0:31] _zy_simnet_cddip2_out_ia_wdata_75_w$;
wire [0:31] _zy_simnet_cddip2_out_ia_wdata_76_w$;
wire [0:12] _zy_simnet_cddip2_out_ia_config_77_w$;
wire [0:11] _zy_simnet_cddip2_out_im_config_78_w$;
wire [0:1] _zy_simnet_dio_79;
wire [0:31] _zy_simnet_cddip3_out_ia_wdata_80_w$;
wire [0:31] _zy_simnet_cddip3_out_ia_wdata_81_w$;
wire [0:31] _zy_simnet_cddip3_out_ia_wdata_82_w$;
wire [0:12] _zy_simnet_cddip3_out_ia_config_83_w$;
wire [0:11] _zy_simnet_cddip3_out_im_config_84_w$;
wire [0:1] _zy_simnet_dio_85;
wire [0:31] _zy_simnet_o_ckv_ia_wdata_part0_86_w$;
wire [0:31] _zy_simnet_o_ckv_ia_wdata_part1_87_w$;
wire [0:18] _zy_simnet_o_ckv_ia_config_88_w$;
wire [0:20] _zy_simnet_o_kim_ia_wdata_part0_89_w$;
wire [0:16] _zy_simnet_o_kim_ia_wdata_part1_90_w$;
wire [0:17] _zy_simnet_o_kim_ia_config_91_w$;
wire [0:15] _zy_simnet_tvar_92;
wire [0:31] _zy_simnet_labels_93_w$;
wire [0:31] _zy_simnet_labels_94_w$;
wire [0:31] _zy_simnet_labels_95_w$;
wire [0:31] _zy_simnet_labels_96_w$;
wire [0:31] _zy_simnet_labels_97_w$;
wire [0:31] _zy_simnet_labels_98_w$;
wire [0:31] _zy_simnet_labels_99_w$;
wire [0:31] _zy_simnet_labels_100_w$;
wire [0:15] _zy_simnet_tvar_101;
wire [0:31] _zy_simnet_labels_102_w$;
wire [0:31] _zy_simnet_labels_103_w$;
wire [0:31] _zy_simnet_labels_104_w$;
wire [0:31] _zy_simnet_labels_105_w$;
wire [0:31] _zy_simnet_labels_106_w$;
wire [0:31] _zy_simnet_labels_107_w$;
wire [0:31] _zy_simnet_labels_108_w$;
wire [0:31] _zy_simnet_labels_109_w$;
wire [0:15] _zy_simnet_tvar_110;
wire [0:31] _zy_simnet_labels_111_w$;
wire [0:31] _zy_simnet_labels_112_w$;
wire [0:31] _zy_simnet_labels_113_w$;
wire [0:31] _zy_simnet_labels_114_w$;
wire [0:31] _zy_simnet_labels_115_w$;
wire [0:31] _zy_simnet_labels_116_w$;
wire [0:31] _zy_simnet_labels_117_w$;
wire [0:31] _zy_simnet_labels_118_w$;
wire [0:15] _zy_simnet_tvar_119;
wire [0:31] _zy_simnet_labels_120_w$;
wire [0:31] _zy_simnet_labels_121_w$;
wire [0:31] _zy_simnet_labels_122_w$;
wire [0:31] _zy_simnet_labels_123_w$;
wire [0:31] _zy_simnet_labels_124_w$;
wire [0:31] _zy_simnet_labels_125_w$;
wire [0:31] _zy_simnet_labels_126_w$;
wire [0:31] _zy_simnet_labels_127_w$;
wire [0:15] _zy_simnet_tvar_128;
wire [0:31] _zy_simnet_labels_129_w$;
wire [0:31] _zy_simnet_labels_130_w$;
wire [0:31] _zy_simnet_labels_131_w$;
wire [0:31] _zy_simnet_labels_132_w$;
wire [0:31] _zy_simnet_labels_133_w$;
wire [0:31] _zy_simnet_labels_134_w$;
wire [0:31] _zy_simnet_labels_135_w$;
wire [0:31] _zy_simnet_labels_136_w$;
wire [0:15] _zy_simnet_tvar_137;
wire [0:31] _zy_simnet_labels_138_w$;
wire [0:31] _zy_simnet_labels_139_w$;
wire [0:31] _zy_simnet_labels_140_w$;
wire [0:31] _zy_simnet_labels_141_w$;
wire [0:31] _zy_simnet_labels_142_w$;
wire [0:31] _zy_simnet_labels_143_w$;
wire [0:31] _zy_simnet_labels_144_w$;
wire [0:31] _zy_simnet_labels_145_w$;
wire [0:15] _zy_simnet_tvar_146;
wire [0:31] _zy_simnet_labels_147_w$;
wire [0:31] _zy_simnet_labels_148_w$;
wire [0:31] _zy_simnet_labels_149_w$;
wire [0:31] _zy_simnet_labels_150_w$;
wire [0:31] _zy_simnet_labels_151_w$;
wire [0:31] _zy_simnet_labels_152_w$;
wire [0:31] _zy_simnet_labels_153_w$;
wire [0:31] _zy_simnet_labels_154_w$;
wire [0:15] _zy_simnet_tvar_155;
wire [0:31] _zy_simnet_labels_156_w$;
wire [0:31] _zy_simnet_labels_157_w$;
wire [0:31] _zy_simnet_labels_158_w$;
wire [0:31] _zy_simnet_labels_159_w$;
wire [0:31] _zy_simnet_labels_160_w$;
wire [0:31] _zy_simnet_labels_161_w$;
wire [0:31] _zy_simnet_labels_162_w$;
wire [0:31] _zy_simnet_labels_163_w$;
wire [0:1] _zy_simnet_o_kdf_drbg_ctrl_164_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_31_0_165_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_63_32_166_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_95_64_167_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_127_96_168_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_159_128_169_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_191_160_170_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_223_192_171_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_255_224_172_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_31_0_173_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_63_32_174_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_95_64_175_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_127_96_176_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_reseed_interval_0_177_w$;
wire [0:15] _zy_simnet_o_kdf_drbg_seed_0_reseed_interval_1_178_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_31_0_179_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_63_32_180_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_95_64_181_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_127_96_182_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_159_128_183_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_191_160_184_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_223_192_185_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_255_224_186_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_31_0_187_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_63_32_188_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_95_64_189_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_127_96_190_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_reseed_interval_0_191_w$;
wire [0:15] _zy_simnet_o_kdf_drbg_seed_1_reseed_interval_1_192_w$;
wire [0:4] _zy_simnet_dio_193;
wire [0:4] _zy_simnet_o_interrupt_mask_194_w$;
wire [0:7] _zy_simnet_o_engine_sticky_status_195_w$;
wire [0:6] _zy_simnet_o_bimc_monitor_mask_196_w$;
wire [0:31] _zy_simnet_o_bimc_ecc_uncorrectable_error_cnt_197_w$;
wire [0:31] _zy_simnet_o_bimc_ecc_correctable_error_cnt_198_w$;
wire [0:31] _zy_simnet_o_bimc_parity_error_cnt_199_w$;
wire [0:31] _zy_simnet_o_bimc_global_config_200_w$;
wire [0:28] _zy_simnet_o_bimc_eccpar_debug_201_w$;
wire [0:10] _zy_simnet_o_bimc_cmd2_202_w$;
wire [0:31] _zy_simnet_o_bimc_cmd1_203_w$;
wire [0:31] _zy_simnet_o_bimc_cmd0_204_w$;
wire [0:9] _zy_simnet_o_bimc_rxcmd2_205_w$;
wire [0:9] _zy_simnet_o_bimc_rxrsp2_206_w$;
wire [0:9] _zy_simnet_o_bimc_pollrsp2_207_w$;
wire [0:9] _zy_simnet_o_bimc_dbgcmd2_208_w$;
wire [0:15] _zy_simnet_dio_209;
wire [0:8] _zy_simnet_tready_override_210_w$;
wire [0:31] _zy_simnet_regs_sa_ctrl_211_w$;
wire [0:31] _zy_simnet_sa_snapshot_ia_wdata_212_w$;
wire [0:31] _zy_simnet_sa_snapshot_ia_wdata_213_w$;
wire [0:8] _zy_simnet_sa_snapshot_ia_config_214_w$;
wire [0:31] _zy_simnet_sa_count_ia_wdata_215_w$;
wire [0:31] _zy_simnet_sa_count_ia_wdata_216_w$;
wire [0:8] _zy_simnet_sa_count_ia_config_217_w$;
wire [0:6] _zy_simnet_cceip_encrypt_kop_fifo_override_218_w$;
wire [0:6] _zy_simnet_cceip_validate_kop_fifo_override_219_w$;
wire [0:6] _zy_simnet_cddip_decrypt_kop_fifo_override_220_w$;
wire [0:31] _zy_simnet_sa_global_ctrl_221_w$;
wire [0:31] _zy_simnet_sa_ctrl_ia_wdata_222_w$;
wire [0:8] _zy_simnet_sa_ctrl_ia_config_223_w$;
wire [0:31] _zy_simnet_blkid_revid_config_224_w$;
wire [0:7] _zy_simnet_revid_wire_225_w$;
wire [0:31] _zy_simnet_tvar_226;
wire [0:19] _zy_simnet_cceip0_out_ia_capability_227_w$;
wire [0:16] _zy_simnet_cceip0_out_ia_status_228_w$;
wire [0:31] _zy_simnet_tvar_229;
wire [0:31] _zy_simnet_tvar_230;
wire [0:31] _zy_simnet_tvar_231;
wire [0:11] _zy_simnet_cceip0_out_im_status_232_w$;
wire [0:1] _zy_simnet_cio_233;
wire [0:19] _zy_simnet_cceip1_out_ia_capability_234_w$;
wire [0:16] _zy_simnet_cceip1_out_ia_status_235_w$;
wire [0:31] _zy_simnet_tvar_236;
wire [0:31] _zy_simnet_tvar_237;
wire [0:31] _zy_simnet_tvar_238;
wire [0:11] _zy_simnet_cceip1_out_im_status_239_w$;
wire [0:1] _zy_simnet_cio_240;
wire [0:19] _zy_simnet_cceip2_out_ia_capability_241_w$;
wire [0:16] _zy_simnet_cceip2_out_ia_status_242_w$;
wire [0:31] _zy_simnet_tvar_243;
wire [0:31] _zy_simnet_tvar_244;
wire [0:31] _zy_simnet_tvar_245;
wire [0:11] _zy_simnet_cceip2_out_im_status_246_w$;
wire [0:1] _zy_simnet_cio_247;
wire [0:19] _zy_simnet_cceip3_out_ia_capability_248_w$;
wire [0:16] _zy_simnet_cceip3_out_ia_status_249_w$;
wire [0:31] _zy_simnet_tvar_250;
wire [0:31] _zy_simnet_tvar_251;
wire [0:31] _zy_simnet_tvar_252;
wire [0:11] _zy_simnet_cceip3_out_im_status_253_w$;
wire [0:1] _zy_simnet_cio_254;
wire [0:19] _zy_simnet_cddip0_out_ia_capability_255_w$;
wire [0:16] _zy_simnet_cddip0_out_ia_status_256_w$;
wire [0:31] _zy_simnet_tvar_257;
wire [0:31] _zy_simnet_tvar_258;
wire [0:31] _zy_simnet_tvar_259;
wire [0:11] _zy_simnet_cddip0_out_im_status_260_w$;
wire [0:1] _zy_simnet_cio_261;
wire [0:19] _zy_simnet_cddip1_out_ia_capability_262_w$;
wire [0:16] _zy_simnet_cddip1_out_ia_status_263_w$;
wire [0:31] _zy_simnet_tvar_264;
wire [0:31] _zy_simnet_tvar_265;
wire [0:31] _zy_simnet_tvar_266;
wire [0:11] _zy_simnet_cddip1_out_im_status_267_w$;
wire [0:1] _zy_simnet_cio_268;
wire [0:19] _zy_simnet_cddip2_out_ia_capability_269_w$;
wire [0:16] _zy_simnet_cddip2_out_ia_status_270_w$;
wire [0:31] _zy_simnet_tvar_271;
wire [0:31] _zy_simnet_tvar_272;
wire [0:31] _zy_simnet_tvar_273;
wire [0:11] _zy_simnet_cddip2_out_im_status_274_w$;
wire [0:1] _zy_simnet_cio_275;
wire [0:19] _zy_simnet_cddip3_out_ia_capability_276_w$;
wire [0:16] _zy_simnet_cddip3_out_ia_status_277_w$;
wire [0:31] _zy_simnet_tvar_278;
wire [0:31] _zy_simnet_tvar_279;
wire [0:31] _zy_simnet_tvar_280;
wire [0:11] _zy_simnet_cddip3_out_im_status_281_w$;
wire [0:1] _zy_simnet_cio_282;
wire [0:19] _zy_simnet_ckv_ia_capability_283_w$;
wire [0:22] _zy_simnet_ckv_ia_status_284_w$;
wire [0:31] _zy_simnet_ckv_ia_rdata_part0_285_w$;
wire [0:31] _zy_simnet_ckv_ia_rdata_part1_286_w$;
wire [0:19] _zy_simnet_kim_ia_capability_287_w$;
wire [0:21] _zy_simnet_kim_ia_status_288_w$;
wire [0:20] _zy_simnet_kim_ia_rdata_part0_289_w$;
wire [0:16] _zy_simnet_kim_ia_rdata_part1_290_w$;
wire [0:1] _zy_simnet_kdf_drbg_ctrl_291_w$;
wire [0:4] _zy_simnet_interrupt_status_292_w$;
wire [0:7] _zy_simnet_engine_sticky_status_293_w$;
wire [0:6] _zy_simnet_bimc_monitor_294_w$;
wire [0:31] _zy_simnet_bimc_ecc_uncorrectable_error_cnt_295_w$;
wire [0:31] _zy_simnet_bimc_ecc_correctable_error_cnt_296_w$;
wire [0:31] _zy_simnet_bimc_parity_error_cnt_297_w$;
wire [0:31] _zy_simnet_bimc_global_config_298_w$;
wire [0:11] _zy_simnet_bimc_memid_299_w$;
wire [0:28] _zy_simnet_bimc_eccpar_debug_300_w$;
wire [0:10] _zy_simnet_bimc_cmd2_301_w$;
wire [0:9] _zy_simnet_bimc_rxcmd2_302_w$;
wire [0:31] _zy_simnet_bimc_rxcmd1_303_w$;
wire [0:31] _zy_simnet_bimc_rxcmd0_304_w$;
wire [0:9] _zy_simnet_bimc_rxrsp2_305_w$;
wire [0:31] _zy_simnet_bimc_rxrsp1_306_w$;
wire [0:31] _zy_simnet_bimc_rxrsp0_307_w$;
wire [0:9] _zy_simnet_bimc_pollrsp2_308_w$;
wire [0:31] _zy_simnet_bimc_pollrsp1_309_w$;
wire [0:31] _zy_simnet_bimc_pollrsp0_310_w$;
wire [0:9] _zy_simnet_bimc_dbgcmd2_311_w$;
wire [0:31] _zy_simnet_bimc_dbgcmd1_312_w$;
wire [0:31] _zy_simnet_bimc_dbgcmd0_313_w$;
wire [0:15] _zy_simnet_im_available_314_w$;
wire [0:15] _zy_simnet_cio_315;
wire [0:8] _zy_simnet_tready_override_316_w$;
wire [0:31] _zy_simnet_regs_sa_ctrl_317_w$;
wire [0:19] _zy_simnet_sa_snapshot_ia_capability_318_w$;
wire [0:12] _zy_simnet_sa_snapshot_ia_status_319_w$;
wire [0:31] _zy_simnet_sa_snapshot_ia_rdata_320_w$;
wire [0:31] _zy_simnet_sa_snapshot_ia_rdata_321_w$;
wire [0:19] _zy_simnet_sa_count_ia_capability_322_w$;
wire [0:12] _zy_simnet_sa_count_ia_status_323_w$;
wire [0:31] _zy_simnet_sa_count_ia_rdata_324_w$;
wire [0:31] _zy_simnet_sa_count_ia_rdata_325_w$;
wire [0:31] _zy_simnet_sa_global_ctrl_326_w$;
wire [0:19] _zy_simnet_sa_ctrl_ia_capability_327_w$;
wire [0:12] _zy_simnet_sa_ctrl_ia_status_328_w$;
wire [0:31] _zy_simnet_sa_ctrl_ia_rdata_329_w$;
wire _zy_simnet_wr_stb_330_w$;
wire _zy_simnet_dio_331;
wire [0:31] _zy_simnet_wr_data_332_w$;
wire [0:10] _zy_simnet_reg_addr_333_w$;
wire [0:15] _zy_simnet_rbus_ring_o_334_w$;
wire _zy_simnet_rbus_ring_o_335_w$;
wire [0:31] _zy_simnet_rbus_ring_o_336_w$;
wire _zy_simnet_rbus_ring_o_337_w$;
wire [0:10] _zy_simnet_locl_addr_338_w$;
wire _zy_simnet_locl_wr_strb_339_w$;
wire [0:31] _zy_simnet_locl_wr_data_340_w$;
wire _zy_simnet_locl_rd_strb_341_w$;
wire [0:31] _zy_simnet_locl_rd_data_342_w$;
wire _zy_simnet_locl_ack_343_w$;
wire _zy_simnet_locl_err_ack_344_w$;
wire [0:31] _zy_simnet_rbus_ring_o_345_w$;
wire _zy_simnet_rbus_ring_o_346_w$;
wire _zy_simnet_rbus_ring_o_347_w$;
wire _zy_simnet_kme_cceip0_ob_in_mod_348_w$;
wire [0:82] _zy_simnet_kme_cceip0_ob_out_post_349_w$;
wire _zy_simnet_cceip0_im_vld_350_w$;
wire _zy_simnet_tvar_351;
wire _zy_simnet_cceip0_im_rdy_352_w$;
wire _zy_simnet_kme_cceip1_ob_in_mod_353_w$;
wire [0:82] _zy_simnet_kme_cceip1_ob_out_post_354_w$;
wire _zy_simnet_cceip1_im_vld_355_w$;
wire _zy_simnet_tvar_356;
wire _zy_simnet_cceip1_im_rdy_357_w$;
wire _zy_simnet_kme_cceip2_ob_in_mod_358_w$;
wire [0:82] _zy_simnet_kme_cceip2_ob_out_post_359_w$;
wire _zy_simnet_cceip2_im_vld_360_w$;
wire _zy_simnet_tvar_361;
wire _zy_simnet_cceip2_im_rdy_362_w$;
wire _zy_simnet_kme_cceip3_ob_in_mod_363_w$;
wire [0:82] _zy_simnet_kme_cceip3_ob_out_post_364_w$;
wire _zy_simnet_cceip3_im_vld_365_w$;
wire _zy_simnet_tvar_366;
wire _zy_simnet_cceip3_im_rdy_367_w$;
wire _zy_simnet_kme_cddip0_ob_in_mod_368_w$;
wire [0:82] _zy_simnet_kme_cddip0_ob_out_post_369_w$;
wire _zy_simnet_cddip0_im_vld_370_w$;
wire _zy_simnet_tvar_371;
wire _zy_simnet_cddip0_im_rdy_372_w$;
wire _zy_simnet_kme_cddip1_ob_in_mod_373_w$;
wire [0:82] _zy_simnet_kme_cddip1_ob_out_post_374_w$;
wire _zy_simnet_cddip1_im_vld_375_w$;
wire _zy_simnet_tvar_376;
wire _zy_simnet_cddip1_im_rdy_377_w$;
wire _zy_simnet_kme_cddip2_ob_in_mod_378_w$;
wire [0:82] _zy_simnet_kme_cddip2_ob_out_post_379_w$;
wire _zy_simnet_cddip2_im_vld_380_w$;
wire _zy_simnet_tvar_381;
wire _zy_simnet_cddip2_im_rdy_382_w$;
wire _zy_simnet_kme_cddip3_ob_in_mod_383_w$;
wire [0:82] _zy_simnet_kme_cddip3_ob_out_post_384_w$;
wire _zy_simnet_cddip3_im_vld_385_w$;
wire _zy_simnet_tvar_386;
wire _zy_simnet_cddip3_im_rdy_387_w$;
wire [0:2] _zy_simnet_cceip0_out_ia_status_388_w$;
wire [0:4] _zy_simnet_cceip0_out_ia_status_389_w$;
wire [0:8] _zy_simnet_cceip0_out_ia_status_390_w$;
wire [0:15] _zy_simnet_cceip0_out_ia_capability_391_w$;
wire [0:3] _zy_simnet_cceip0_out_ia_capability_392_w$;
wire [0:95] _zy_simnet_cceip0_out_ia_rdata_393_w$;
wire _zy_simnet_cceip1_ism_idat_394_w$;
wire _zy_simnet_cceip1_ism_isync_395_w$;
wire _zy_simnet_cceip0_ism_mbe_396_w$;
wire _zy_simnet_cceip0_im_rdy_397_w$;
wire [0:1] _zy_simnet_im_available_kme_cceip0_398_w$;
wire [0:11] _zy_simnet_cceip0_out_im_status_399_w$;
wire [0:10] _zy_simnet_reg_addr_400_w$;
wire [0:3] _zy_simnet_cceip0_out_ia_config_401_w$;
wire [0:8] _zy_simnet_cceip0_out_ia_config_402_w$;
wire _zy_simnet_wr_stb_403_w$;
wire [0:95] _zy_simnet_cceip0_out_ia_wdata_404_w$;
wire _zy_simnet_cio_405;
wire _zy_simnet_cceip0_ism_bimc_isync_406_w$;
wire _zy_simnet_cceip0_ism_bimc_idat_407_w$;
wire [0:95] _zy_simnet_cceip0_im_din_408_w$;
wire _zy_simnet_cceip0_im_vld_409_w$;
wire [0:1] _zy_simnet_im_consumed_kme_cceip0_410_w$;
wire [0:11] _zy_simnet_cceip0_out_im_config_411_w$;
wire [0:2] _zy_simnet_cceip1_out_ia_status_412_w$;
wire [0:4] _zy_simnet_cceip1_out_ia_status_413_w$;
wire [0:8] _zy_simnet_cceip1_out_ia_status_414_w$;
wire [0:15] _zy_simnet_cceip1_out_ia_capability_415_w$;
wire [0:3] _zy_simnet_cceip1_out_ia_capability_416_w$;
wire [0:95] _zy_simnet_cceip1_out_ia_rdata_417_w$;
wire _zy_simnet_cceip2_ism_idat_418_w$;
wire _zy_simnet_cceip2_ism_isync_419_w$;
wire _zy_simnet_cceip1_ism_mbe_420_w$;
wire _zy_simnet_cceip1_im_rdy_421_w$;
wire [0:1] _zy_simnet_im_available_kme_cceip1_422_w$;
wire [0:11] _zy_simnet_cceip1_out_im_status_423_w$;
wire [0:10] _zy_simnet_reg_addr_424_w$;
wire [0:3] _zy_simnet_cceip1_out_ia_config_425_w$;
wire [0:8] _zy_simnet_cceip1_out_ia_config_426_w$;
wire _zy_simnet_wr_stb_427_w$;
wire [0:95] _zy_simnet_cceip1_out_ia_wdata_428_w$;
wire _zy_simnet_cio_429;
wire _zy_simnet_cceip1_ism_isync_430_w$;
wire _zy_simnet_cceip1_ism_idat_431_w$;
wire [0:95] _zy_simnet_cceip1_im_din_432_w$;
wire _zy_simnet_cceip1_im_vld_433_w$;
wire [0:1] _zy_simnet_im_consumed_kme_cceip1_434_w$;
wire [0:11] _zy_simnet_cceip1_out_im_config_435_w$;
wire [0:2] _zy_simnet_cceip2_out_ia_status_436_w$;
wire [0:4] _zy_simnet_cceip2_out_ia_status_437_w$;
wire [0:8] _zy_simnet_cceip2_out_ia_status_438_w$;
wire [0:15] _zy_simnet_cceip2_out_ia_capability_439_w$;
wire [0:3] _zy_simnet_cceip2_out_ia_capability_440_w$;
wire [0:95] _zy_simnet_cceip2_out_ia_rdata_441_w$;
wire _zy_simnet_cceip3_ism_idat_442_w$;
wire _zy_simnet_cceip3_ism_isync_443_w$;
wire _zy_simnet_cceip2_ism_mbe_444_w$;
wire _zy_simnet_cceip2_im_rdy_445_w$;
wire [0:1] _zy_simnet_im_available_kme_cceip2_446_w$;
wire [0:11] _zy_simnet_cceip2_out_im_status_447_w$;
wire [0:10] _zy_simnet_reg_addr_448_w$;
wire [0:3] _zy_simnet_cceip2_out_ia_config_449_w$;
wire [0:8] _zy_simnet_cceip2_out_ia_config_450_w$;
wire _zy_simnet_wr_stb_451_w$;
wire [0:95] _zy_simnet_cceip2_out_ia_wdata_452_w$;
wire _zy_simnet_cio_453;
wire _zy_simnet_cceip2_ism_isync_454_w$;
wire _zy_simnet_cceip2_ism_idat_455_w$;
wire [0:95] _zy_simnet_cceip2_im_din_456_w$;
wire _zy_simnet_cceip2_im_vld_457_w$;
wire [0:1] _zy_simnet_im_consumed_kme_cceip2_458_w$;
wire [0:11] _zy_simnet_cceip2_out_im_config_459_w$;
wire [0:2] _zy_simnet_cceip3_out_ia_status_460_w$;
wire [0:4] _zy_simnet_cceip3_out_ia_status_461_w$;
wire [0:8] _zy_simnet_cceip3_out_ia_status_462_w$;
wire [0:15] _zy_simnet_cceip3_out_ia_capability_463_w$;
wire [0:3] _zy_simnet_cceip3_out_ia_capability_464_w$;
wire [0:95] _zy_simnet_cceip3_out_ia_rdata_465_w$;
wire _zy_simnet_cddip0_ism_idat_466_w$;
wire _zy_simnet_cddip0_ism_isync_467_w$;
wire _zy_simnet_cceip3_ism_mbe_468_w$;
wire _zy_simnet_cceip3_im_rdy_469_w$;
wire [0:1] _zy_simnet_im_available_kme_cceip3_470_w$;
wire [0:11] _zy_simnet_cceip3_out_im_status_471_w$;
wire [0:10] _zy_simnet_reg_addr_472_w$;
wire [0:3] _zy_simnet_cceip3_out_ia_config_473_w$;
wire [0:8] _zy_simnet_cceip3_out_ia_config_474_w$;
wire _zy_simnet_wr_stb_475_w$;
wire [0:95] _zy_simnet_cceip3_out_ia_wdata_476_w$;
wire _zy_simnet_cio_477;
wire _zy_simnet_cceip3_ism_isync_478_w$;
wire _zy_simnet_cceip3_ism_idat_479_w$;
wire [0:95] _zy_simnet_cceip3_im_din_480_w$;
wire _zy_simnet_cceip3_im_vld_481_w$;
wire [0:1] _zy_simnet_im_consumed_kme_cceip3_482_w$;
wire [0:11] _zy_simnet_cceip3_out_im_config_483_w$;
wire [0:2] _zy_simnet_cddip0_out_ia_status_484_w$;
wire [0:4] _zy_simnet_cddip0_out_ia_status_485_w$;
wire [0:8] _zy_simnet_cddip0_out_ia_status_486_w$;
wire [0:15] _zy_simnet_cddip0_out_ia_capability_487_w$;
wire [0:3] _zy_simnet_cddip0_out_ia_capability_488_w$;
wire [0:95] _zy_simnet_cddip0_out_ia_rdata_489_w$;
wire _zy_simnet_cddip1_ism_idat_490_w$;
wire _zy_simnet_cddip1_ism_isync_491_w$;
wire _zy_simnet_cddip0_ism_mbe_492_w$;
wire _zy_simnet_cddip0_im_rdy_493_w$;
wire [0:1] _zy_simnet_im_available_kme_cddip0_494_w$;
wire [0:11] _zy_simnet_cddip0_out_im_status_495_w$;
wire [0:10] _zy_simnet_reg_addr_496_w$;
wire [0:3] _zy_simnet_cddip0_out_ia_config_497_w$;
wire [0:8] _zy_simnet_cddip0_out_ia_config_498_w$;
wire _zy_simnet_wr_stb_499_w$;
wire [0:95] _zy_simnet_cddip0_out_ia_wdata_500_w$;
wire _zy_simnet_cio_501;
wire _zy_simnet_cddip0_ism_isync_502_w$;
wire _zy_simnet_cddip0_ism_idat_503_w$;
wire [0:95] _zy_simnet_cddip0_im_din_504_w$;
wire _zy_simnet_cddip0_im_vld_505_w$;
wire [0:1] _zy_simnet_im_consumed_kme_cddip0_506_w$;
wire [0:11] _zy_simnet_cddip0_out_im_config_507_w$;
wire [0:2] _zy_simnet_cddip1_out_ia_status_508_w$;
wire [0:4] _zy_simnet_cddip1_out_ia_status_509_w$;
wire [0:8] _zy_simnet_cddip1_out_ia_status_510_w$;
wire [0:15] _zy_simnet_cddip1_out_ia_capability_511_w$;
wire [0:3] _zy_simnet_cddip1_out_ia_capability_512_w$;
wire [0:95] _zy_simnet_cddip1_out_ia_rdata_513_w$;
wire _zy_simnet_cddip2_ism_idat_514_w$;
wire _zy_simnet_cddip2_ism_isync_515_w$;
wire _zy_simnet_cddip1_ism_mbe_516_w$;
wire _zy_simnet_cddip1_im_rdy_517_w$;
wire [0:1] _zy_simnet_im_available_kme_cddip1_518_w$;
wire [0:11] _zy_simnet_cddip1_out_im_status_519_w$;
wire [0:10] _zy_simnet_reg_addr_520_w$;
wire [0:3] _zy_simnet_cddip1_out_ia_config_521_w$;
wire [0:8] _zy_simnet_cddip1_out_ia_config_522_w$;
wire _zy_simnet_wr_stb_523_w$;
wire [0:95] _zy_simnet_cddip1_out_ia_wdata_524_w$;
wire _zy_simnet_cio_525;
wire _zy_simnet_cddip1_ism_isync_526_w$;
wire _zy_simnet_cddip1_ism_idat_527_w$;
wire [0:95] _zy_simnet_cddip1_im_din_528_w$;
wire _zy_simnet_cddip1_im_vld_529_w$;
wire [0:1] _zy_simnet_im_consumed_kme_cddip1_530_w$;
wire [0:11] _zy_simnet_cddip1_out_im_config_531_w$;
wire [0:2] _zy_simnet_cddip2_out_ia_status_532_w$;
wire [0:4] _zy_simnet_cddip2_out_ia_status_533_w$;
wire [0:8] _zy_simnet_cddip2_out_ia_status_534_w$;
wire [0:15] _zy_simnet_cddip2_out_ia_capability_535_w$;
wire [0:3] _zy_simnet_cddip2_out_ia_capability_536_w$;
wire [0:95] _zy_simnet_cddip2_out_ia_rdata_537_w$;
wire _zy_simnet_cddip3_ism_idat_538_w$;
wire _zy_simnet_cddip3_ism_isync_539_w$;
wire _zy_simnet_cddip2_ism_mbe_540_w$;
wire _zy_simnet_cddip2_im_rdy_541_w$;
wire [0:1] _zy_simnet_im_available_kme_cddip2_542_w$;
wire [0:11] _zy_simnet_cddip2_out_im_status_543_w$;
wire [0:10] _zy_simnet_reg_addr_544_w$;
wire [0:3] _zy_simnet_cddip2_out_ia_config_545_w$;
wire [0:8] _zy_simnet_cddip2_out_ia_config_546_w$;
wire _zy_simnet_wr_stb_547_w$;
wire [0:95] _zy_simnet_cddip2_out_ia_wdata_548_w$;
wire _zy_simnet_cio_549;
wire _zy_simnet_cddip2_ism_isync_550_w$;
wire _zy_simnet_cddip2_ism_idat_551_w$;
wire [0:95] _zy_simnet_cddip2_im_din_552_w$;
wire _zy_simnet_cddip2_im_vld_553_w$;
wire [0:1] _zy_simnet_im_consumed_kme_cddip2_554_w$;
wire [0:11] _zy_simnet_cddip2_out_im_config_555_w$;
wire [0:2] _zy_simnet_cddip3_out_ia_status_556_w$;
wire [0:4] _zy_simnet_cddip3_out_ia_status_557_w$;
wire [0:8] _zy_simnet_cddip3_out_ia_status_558_w$;
wire [0:15] _zy_simnet_cddip3_out_ia_capability_559_w$;
wire [0:3] _zy_simnet_cddip3_out_ia_capability_560_w$;
wire [0:95] _zy_simnet_cddip3_out_ia_rdata_561_w$;
wire _zy_simnet_cddip3_ism_odat_562_w$;
wire _zy_simnet_cddip3_ism_osync_563_w$;
wire _zy_simnet_cddip3_ism_mbe_564_w$;
wire _zy_simnet_cddip3_im_rdy_565_w$;
wire [0:1] _zy_simnet_im_available_kme_cddip3_566_w$;
wire [0:11] _zy_simnet_cddip3_out_im_status_567_w$;
wire [0:10] _zy_simnet_reg_addr_568_w$;
wire [0:3] _zy_simnet_cddip3_out_ia_config_569_w$;
wire [0:8] _zy_simnet_cddip3_out_ia_config_570_w$;
wire _zy_simnet_wr_stb_571_w$;
wire [0:95] _zy_simnet_cddip3_out_ia_wdata_572_w$;
wire _zy_simnet_cio_573;
wire _zy_simnet_cddip3_ism_isync_574_w$;
wire _zy_simnet_cddip3_ism_idat_575_w$;
wire [0:95] _zy_simnet_cddip3_im_din_576_w$;
wire _zy_simnet_cddip3_im_vld_577_w$;
wire [0:1] _zy_simnet_im_consumed_kme_cddip3_578_w$;
wire [0:11] _zy_simnet_cddip3_out_im_config_579_w$;
wire [0:3] _zy_simnet_ckv_cmnd_op_580_w$;
wire [0:14] _zy_simnet_ckv_cmnd_addr_581_w$;
wire [0:63] _zy_simnet_ckv_wr_dat_582_w$;
wire [0:19] _zy_simnet_ckv_ia_capability_583_w$;
wire [0:31] _zy_simnet_ckv_ia_rdata_part0_584_w$;
wire [0:31] _zy_simnet_ckv_ia_rdata_part1_585_w$;
wire [0:22] _zy_simnet_ckv_ia_status_586_w$;
wire [0:3] _zy_simnet_kim_cmnd_op_587_w$;
wire [0:13] _zy_simnet_kim_cmnd_addr_588_w$;
wire [0:37] _zy_simnet_kim_wr_dat_589_w$;
wire [0:19] _zy_simnet_kim_ia_capability_590_w$;
wire [0:20] _zy_simnet_kim_ia_rdata_part0_591_w$;
wire [0:16] _zy_simnet_kim_ia_rdata_part1_592_w$;
wire [0:21] _zy_simnet_kim_ia_status_593_w$;
wire [0:7] _zy_simnet_engine_sticky_status_594_w$;
wire _zy_simnet_disable_ckv_kim_ism_reads_595_w$;
wire _zy_simnet_send_kme_ib_beat_596_w$;
wire [0:82] _zy_simnet_kme_cceip0_ob_out_597_w$;
wire [0:82] _zy_simnet_kme_cceip1_ob_out_598_w$;
wire [0:82] _zy_simnet_kme_cceip2_ob_out_599_w$;
wire [0:82] _zy_simnet_kme_cceip3_ob_out_600_w$;
wire [0:82] _zy_simnet_kme_cddip0_ob_out_601_w$;
wire [0:82] _zy_simnet_kme_cddip1_ob_out_602_w$;
wire [0:82] _zy_simnet_kme_cddip2_ob_out_603_w$;
wire [0:82] _zy_simnet_kme_cddip3_ob_out_604_w$;
wire _zy_simnet_axi_term_bimc_isync_605_w$;
wire _zy_simnet_axi_term_bimc_idat_606_w$;
wire [0:2] _zy_simnet_ckv_stat_code_607_w$;
wire [0:4] _zy_simnet_ckv_stat_datawords_608_w$;
wire [0:14] _zy_simnet_ckv_stat_addr_609_w$;
wire [0:3] _zy_simnet_ckv_capability_type_610_w$;
wire [0:15] _zy_simnet_ckv_capability_lst_611_w$;
wire [0:63] _zy_simnet_ckv_rd_dat_612_w$;
wire [0:18] _zy_simnet_o_ckv_ia_config_613_w$;
wire [0:31] _zy_simnet_o_ckv_ia_wdata_part0_614_w$;
wire [0:31] _zy_simnet_o_ckv_ia_wdata_part1_615_w$;
wire [0:2] _zy_simnet_kim_stat_code_616_w$;
wire [0:4] _zy_simnet_kim_stat_datawords_617_w$;
wire [0:13] _zy_simnet_kim_stat_addr_618_w$;
wire [0:3] _zy_simnet_kim_capability_type_619_w$;
wire [0:15] _zy_simnet_kim_capability_lst_620_w$;
wire [0:37] _zy_simnet_kim_rd_dat_621_w$;
wire [0:17] _zy_simnet_o_kim_ia_config_622_w$;
wire [0:20] _zy_simnet_o_kim_ia_wdata_part0_623_w$;
wire [0:16] _zy_simnet_o_kim_ia_wdata_part1_624_w$;
wire _zy_simnet_wr_stb_625_w$;
wire [0:31] _zy_simnet_wr_data_626_w$;
wire [0:10] _zy_simnet_reg_addr_627_w$;
wire [0:7] _zy_simnet_o_engine_sticky_status_628_w$;
wire _zy_simnet_o_disable_ckv_kim_ism_reads_629_w$;
wire _zy_simnet_o_send_kme_ib_beat_630_w$;
wire [0:95] _zy_simnet_cceip0_out_ia_wdata_631_w$;
wire [0:8] _zy_simnet_tready_override_632_w$;
wire [0:82] _zy_simnet_kme_cceip0_ob_out_post_633_w$;
wire [0:82] _zy_simnet_kme_cceip1_ob_out_post_634_w$;
wire [0:82] _zy_simnet_kme_cceip2_ob_out_post_635_w$;
wire [0:82] _zy_simnet_kme_cceip3_ob_out_post_636_w$;
wire [0:82] _zy_simnet_kme_cddip0_ob_out_post_637_w$;
wire [0:82] _zy_simnet_kme_cddip1_ob_out_post_638_w$;
wire [0:82] _zy_simnet_kme_cddip2_ob_out_post_639_w$;
wire [0:82] _zy_simnet_kme_cddip3_ob_out_post_640_w$;
wire _zy_simnet_cddip3_ism_osync_641_w$;
wire _zy_simnet_cddip3_ism_odat_642_w$;
wire [0:10] _zy_simnet_reg_addr_643_w$;
wire [0:3] _zy_simnet_ckv_cmnd_op_644_w$;
wire [0:14] _zy_simnet_ckv_cmnd_addr_645_w$;
wire [0:2] _zy_simnet_ckv_stat_code_646_w$;
wire [0:4] _zy_simnet_ckv_stat_datawords_647_w$;
wire [0:14] _zy_simnet_ckv_stat_addr_648_w$;
wire [0:15] _zy_simnet_ckv_capability_lst_649_w$;
wire [0:3] _zy_simnet_ckv_capability_type_650_w$;
wire _zy_simnet_wr_stb_651_w$;
wire [0:63] _zy_simnet_ckv_wr_dat_652_w$;
wire [0:63] _zy_simnet_ckv_rd_dat_653_w$;
wire _zy_simnet_cio_654;
wire _zy_simnet_ckv_bimc_isync_655_w$;
wire _zy_simnet_ckv_bimc_idat_656_w$;
wire _zy_simnet_cceip0_ism_bimc_idat_657_w$;
wire _zy_simnet_cceip0_ism_bimc_isync_658_w$;
wire _zy_simnet_cio_659;
wire [0:63] _zy_simnet_cio_660;
wire [0:63] _zy_simnet_cio_661;
wire _zy_simnet_dio_662;
wire [0:10] _zy_simnet_reg_addr_663_w$;
wire [0:3] _zy_simnet_kim_cmnd_op_664_w$;
wire [0:13] _zy_simnet_kim_cmnd_addr_665_w$;
wire [0:2] _zy_simnet_kim_stat_code_666_w$;
wire [0:4] _zy_simnet_kim_stat_datawords_667_w$;
wire [0:13] _zy_simnet_kim_stat_addr_668_w$;
wire [0:15] _zy_simnet_kim_capability_lst_669_w$;
wire [0:3] _zy_simnet_kim_capability_type_670_w$;
wire _zy_simnet_wr_stb_671_w$;
wire [0:37] _zy_simnet_kim_wr_dat_672_w$;
wire [0:37] _zy_simnet_kim_rd_dat_673_w$;
wire _zy_simnet_cio_674;
wire _zy_simnet_kim_bimc_isync_675_w$;
wire _zy_simnet_kim_bimc_idat_676_w$;
wire _zy_simnet_ckv_bimc_idat_677_w$;
wire _zy_simnet_ckv_bimc_isync_678_w$;
wire _zy_simnet_cio_679;
wire [0:37] _zy_simnet_cio_680;
wire [0:37] _zy_simnet_cio_681;
wire [0:37] _zy_simnet_kim_dout_682_w$;
wire _zy_simnet_dio_683;
wire _zy_simnet_set_drbg_expired_int_684_w$;
wire [0:1] _zy_simnet_kdf_drbg_ctrl_685_w$;
wire _zy_simnet_wr_stb_686_w$;
wire [0:31] _zy_simnet_wr_data_687_w$;
wire [0:10] _zy_simnet_reg_addr_688_w$;
wire [0:1] _zy_simnet_o_kdf_drbg_ctrl_689_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_reseed_interval_0_690_w$;
wire [0:15] _zy_simnet_o_kdf_drbg_seed_0_reseed_interval_1_691_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_127_96_692_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_159_128_693_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_191_160_694_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_223_192_695_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_255_224_696_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_31_0_697_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_63_32_698_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_key_95_64_699_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_127_96_700_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_31_0_701_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_63_32_702_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_0_state_value_95_64_703_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_reseed_interval_0_704_w$;
wire [0:15] _zy_simnet_o_kdf_drbg_seed_1_reseed_interval_1_705_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_127_96_706_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_159_128_707_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_191_160_708_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_223_192_709_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_255_224_710_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_31_0_711_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_63_32_712_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_key_95_64_713_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_127_96_714_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_31_0_715_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_63_32_716_w$;
wire [0:31] _zy_simnet_o_kdf_drbg_seed_1_state_value_95_64_717_w$;
wire _zy_simnet_dio_718;
wire _zy_simnet_bimc_interrupt_719_w$;
wire _zy_simnet_kim_bimc_idat_720_w$;
wire _zy_simnet_kim_bimc_isync_721_w$;
wire _zy_simnet_axi_term_bimc_idat_722_w$;
wire _zy_simnet_axi_term_bimc_isync_723_w$;
wire [0:6] _zy_simnet_o_bimc_monitor_mask_724_w$;
wire [0:31] _zy_simnet_o_bimc_ecc_uncorrectable_error_cnt_725_w$;
wire [0:31] _zy_simnet_o_bimc_ecc_correctable_error_cnt_726_w$;
wire [0:31] _zy_simnet_o_bimc_parity_error_cnt_727_w$;
wire [0:31] _zy_simnet_o_bimc_global_config_728_w$;
wire [0:28] _zy_simnet_o_bimc_eccpar_debug_729_w$;
wire [0:10] _zy_simnet_o_bimc_cmd2_730_w$;
wire [0:31] _zy_simnet_o_bimc_cmd1_731_w$;
wire [0:31] _zy_simnet_o_bimc_cmd0_732_w$;
wire [0:9] _zy_simnet_o_bimc_rxcmd2_733_w$;
wire [0:9] _zy_simnet_o_bimc_rxrsp2_734_w$;
wire [0:9] _zy_simnet_o_bimc_pollrsp2_735_w$;
wire [0:9] _zy_simnet_o_bimc_dbgcmd2_736_w$;
wire [0:6] _zy_simnet_bimc_monitor_737_w$;
wire [0:31] _zy_simnet_bimc_ecc_uncorrectable_error_cnt_738_w$;
wire [0:31] _zy_simnet_bimc_ecc_correctable_error_cnt_739_w$;
wire [0:31] _zy_simnet_bimc_parity_error_cnt_740_w$;
wire [0:31] _zy_simnet_bimc_global_config_741_w$;
wire [0:11] _zy_simnet_bimc_memid_742_w$;
wire [0:28] _zy_simnet_bimc_eccpar_debug_743_w$;
wire [0:10] _zy_simnet_bimc_cmd2_744_w$;
wire [0:9] _zy_simnet_bimc_rxcmd2_745_w$;
wire [0:31] _zy_simnet_bimc_rxcmd1_746_w$;
wire [0:31] _zy_simnet_bimc_rxcmd0_747_w$;
wire [0:9] _zy_simnet_bimc_rxrsp2_748_w$;
wire [0:31] _zy_simnet_bimc_rxrsp1_749_w$;
wire [0:31] _zy_simnet_bimc_rxrsp0_750_w$;
wire [0:9] _zy_simnet_bimc_pollrsp2_751_w$;
wire [0:31] _zy_simnet_bimc_pollrsp1_752_w$;
wire [0:31] _zy_simnet_bimc_pollrsp0_753_w$;
wire [0:9] _zy_simnet_bimc_dbgcmd2_754_w$;
wire [0:31] _zy_simnet_bimc_dbgcmd1_755_w$;
wire [0:31] _zy_simnet_bimc_dbgcmd0_756_w$;
wire [0:4] _zy_simnet_interrupt_status_757_w$;
wire _zy_simnet_set_drbg_expired_int_758_w$;
wire _zy_simnet_cceip0_ism_mbe_759_w$;
wire _zy_simnet_cceip1_ism_mbe_760_w$;
wire _zy_simnet_cceip2_ism_mbe_761_w$;
wire _zy_simnet_cceip3_ism_mbe_762_w$;
wire _zy_simnet_cddip0_ism_mbe_763_w$;
wire _zy_simnet_cddip1_ism_mbe_764_w$;
wire _zy_simnet_cddip2_ism_mbe_765_w$;
wire _zy_simnet_cddip3_ism_mbe_766_w$;
wire _zy_simnet_bimc_interrupt_767_w$;
wire _zy_simnet_wr_stb_768_w$;
wire [0:31] _zy_simnet_wr_data_769_w$;
wire [0:10] _zy_simnet_reg_addr_770_w$;
wire [0:4] _zy_simnet_o_interrupt_mask_771_w$;
wire [0:2] _zy_simnet_sa_snapshot_ia_status_772_w$;
wire [0:4] _zy_simnet_sa_snapshot_ia_status_773_w$;
wire [0:4] _zy_simnet_sa_snapshot_ia_status_774_w$;
wire [0:15] _zy_simnet_sa_snapshot_ia_capability_775_w$;
wire [0:3] _zy_simnet_sa_snapshot_ia_capability_776_w$;
wire [0:63] _zy_simnet_sa_snapshot_ia_rdata_777_w$;
wire [0:10] _zy_simnet_reg_addr_778_w$;
wire [0:3] _zy_simnet_sa_snapshot_ia_config_779_w$;
wire [0:4] _zy_simnet_sa_snapshot_ia_config_780_w$;
wire _zy_simnet_wr_stb_781_w$;
wire [0:63] _zy_simnet_sa_snapshot_ia_wdata_782_w$;
wire [0:2] _zy_simnet_sa_count_ia_status_783_w$;
wire [0:4] _zy_simnet_sa_count_ia_status_784_w$;
wire [0:4] _zy_simnet_sa_count_ia_status_785_w$;
wire [0:15] _zy_simnet_sa_count_ia_capability_786_w$;
wire [0:3] _zy_simnet_sa_count_ia_capability_787_w$;
wire [0:63] _zy_simnet_sa_count_ia_rdata_788_w$;
wire [0:10] _zy_simnet_reg_addr_789_w$;
wire [0:3] _zy_simnet_sa_count_ia_config_790_w$;
wire [0:4] _zy_simnet_sa_count_ia_config_791_w$;
wire _zy_simnet_wr_stb_792_w$;
wire [0:63] _zy_simnet_sa_count_ia_wdata_793_w$;
wire [0:2] _zy_simnet_sa_ctrl_ia_status_794_w$;
wire [0:4] _zy_simnet_sa_ctrl_ia_status_795_w$;
wire [0:4] _zy_simnet_sa_ctrl_ia_status_796_w$;
wire [0:15] _zy_simnet_sa_ctrl_ia_capability_797_w$;
wire [0:3] _zy_simnet_sa_ctrl_ia_capability_798_w$;
wire [0:31] _zy_simnet_sa_ctrl_ia_rdata_799_w$;
wire [0:10] _zy_simnet_reg_addr_800_w$;
wire [0:3] _zy_simnet_sa_ctrl_ia_config_801_w$;
wire [0:4] _zy_simnet_sa_ctrl_ia_config_802_w$;
wire _zy_simnet_wr_stb_803_w$;
wire [0:31] _zy_simnet_sa_ctrl_ia_wdata_804_w$;
wire axi_term_bimc_idat;
wire axi_term_bimc_isync;
wire [10:0] bimc_cmd2;
wire [31:0] bimc_dbgcmd0;
wire [31:0] bimc_dbgcmd1;
wire [9:0] bimc_dbgcmd2;
wire [31:0] bimc_ecc_correctable_error_cnt;
wire [31:0] bimc_ecc_uncorrectable_error_cnt;
wire [28:0] bimc_eccpar_debug;
wire [31:0] bimc_global_config;
wire bimc_interrupt;
wire [11:0] bimc_memid;
wire [6:0] bimc_monitor;
wire [31:0] bimc_parity_error_cnt;
wire [31:0] bimc_pollrsp0;
wire [31:0] bimc_pollrsp1;
wire [9:0] bimc_pollrsp2;
wire [31:0] bimc_rxcmd0;
wire [31:0] bimc_rxcmd1;
wire [9:0] bimc_rxcmd2;
wire [31:0] bimc_rxrsp0;
wire [31:0] bimc_rxrsp1;
wire [9:0] bimc_rxrsp2;
wire cceip0_im_rdy;
wire cceip0_ism_bimc_idat;
wire cceip0_ism_bimc_isync;
wire cceip0_ism_mbe;
wire cceip1_im_rdy;
wire cceip1_ism_idat;
wire cceip1_ism_isync;
wire cceip1_ism_mbe;
wire cceip2_im_rdy;
wire cceip2_ism_idat;
wire cceip2_ism_isync;
wire cceip2_ism_mbe;
wire cceip3_im_rdy;
wire cceip3_ism_idat;
wire cceip3_ism_isync;
wire cceip3_ism_mbe;
wire cddip0_im_rdy;
wire cddip0_ism_idat;
wire cddip0_ism_isync;
wire cddip0_ism_mbe;
wire cddip1_im_rdy;
wire cddip1_ism_idat;
wire cddip1_ism_isync;
wire cddip1_ism_mbe;
wire cddip2_im_rdy;
wire cddip2_ism_idat;
wire cddip2_ism_isync;
wire cddip2_ism_mbe;
wire cddip3_im_rdy;
wire cddip3_ism_idat;
wire cddip3_ism_isync;
wire cddip3_ism_mbe;
wire cddip3_ism_odat;
wire cddip3_ism_osync;
wire ckv_bimc_idat;
wire ckv_bimc_isync;
wire [15:0] ckv_capability_lst;
wire [3:0] ckv_capability_type;
wire [14:0] ckv_cmnd_addr;
wire [3:0] ckv_cmnd_op;
wire [19:0] ckv_ia_capability;
wire [31:0] ckv_ia_rdata_part0;
wire [31:0] ckv_ia_rdata_part1;
wire [22:0] ckv_ia_status;
wire [63:0] ckv_rd_dat;
wire [14:0] ckv_stat_addr;
wire [2:0] ckv_stat_code;
wire [4:0] ckv_stat_datawords;
wire [63:0] ckv_wr_dat;
wire disable_ckv_kim_ism_reads;
wire [7:0] engine_sticky_status;
wire [4:0] interrupt_status;
wire [1:0] kdf_drbg_ctrl;
wire kim_bimc_idat;
wire kim_bimc_isync;
wire [15:0] kim_capability_lst;
wire [3:0] kim_capability_type;
wire [13:0] kim_cmnd_addr;
wire [3:0] kim_cmnd_op;
wire [19:0] kim_ia_capability;
wire [20:0] kim_ia_rdata_part0;
wire [16:0] kim_ia_rdata_part1;
wire [21:0] kim_ia_status;
wire [37:0] kim_rd_dat;
wire [13:0] kim_stat_addr;
wire [2:0] kim_stat_code;
wire [4:0] kim_stat_datawords;
wire [37:0] kim_wr_dat;
wire locl_ack;
wire locl_err_ack;
wire [31:0] locl_rd_data;
wire locl_rd_strb;
wire locl_wr_strb;
wire [31:0] o_bimc_cmd0;
wire [31:0] o_bimc_cmd1;
wire [10:0] o_bimc_cmd2;
wire [9:0] o_bimc_dbgcmd2;
wire [31:0] o_bimc_ecc_correctable_error_cnt;
wire [31:0] o_bimc_ecc_uncorrectable_error_cnt;
wire [28:0] o_bimc_eccpar_debug;
wire [31:0] o_bimc_global_config;
wire [6:0] o_bimc_monitor_mask;
wire [31:0] o_bimc_parity_error_cnt;
wire [9:0] o_bimc_pollrsp2;
wire [9:0] o_bimc_rxcmd2;
wire [9:0] o_bimc_rxrsp2;
wire [18:0] o_ckv_ia_config;
wire [31:0] o_ckv_ia_wdata_part0;
wire [31:0] o_ckv_ia_wdata_part1;
wire o_disable_ckv_kim_ism_reads;
wire [7:0] o_engine_sticky_status;
wire [4:0] o_interrupt_mask;
wire [1:0] o_kdf_drbg_ctrl;
wire [31:0] o_kdf_drbg_seed_0_reseed_interval_0;
wire [15:0] o_kdf_drbg_seed_0_reseed_interval_1;
wire [31:0] o_kdf_drbg_seed_0_state_key_127_96;
wire [31:0] o_kdf_drbg_seed_0_state_key_159_128;
wire [31:0] o_kdf_drbg_seed_0_state_key_191_160;
wire [31:0] o_kdf_drbg_seed_0_state_key_223_192;
wire [31:0] o_kdf_drbg_seed_0_state_key_255_224;
wire [31:0] o_kdf_drbg_seed_0_state_key_31_0;
wire [31:0] o_kdf_drbg_seed_0_state_key_63_32;
wire [31:0] o_kdf_drbg_seed_0_state_key_95_64;
wire [31:0] o_kdf_drbg_seed_0_state_value_127_96;
wire [31:0] o_kdf_drbg_seed_0_state_value_31_0;
wire [31:0] o_kdf_drbg_seed_0_state_value_63_32;
wire [31:0] o_kdf_drbg_seed_0_state_value_95_64;
wire [31:0] o_kdf_drbg_seed_1_reseed_interval_0;
wire [15:0] o_kdf_drbg_seed_1_reseed_interval_1;
wire [31:0] o_kdf_drbg_seed_1_state_key_127_96;
wire [31:0] o_kdf_drbg_seed_1_state_key_159_128;
wire [31:0] o_kdf_drbg_seed_1_state_key_191_160;
wire [31:0] o_kdf_drbg_seed_1_state_key_223_192;
wire [31:0] o_kdf_drbg_seed_1_state_key_255_224;
wire [31:0] o_kdf_drbg_seed_1_state_key_31_0;
wire [31:0] o_kdf_drbg_seed_1_state_key_63_32;
wire [31:0] o_kdf_drbg_seed_1_state_key_95_64;
wire [31:0] o_kdf_drbg_seed_1_state_value_127_96;
wire [31:0] o_kdf_drbg_seed_1_state_value_31_0;
wire [31:0] o_kdf_drbg_seed_1_state_value_63_32;
wire [31:0] o_kdf_drbg_seed_1_state_value_95_64;
wire [17:0] o_kim_ia_config;
wire [20:0] o_kim_ia_wdata_part0;
wire [16:0] o_kim_ia_wdata_part1;
wire o_send_kme_ib_beat;
wire o_tready_override_val;
wire [31:0] regs_sa_ctrl;
wire send_kme_ib_beat;
wire set_drbg_expired_int;
wire [31:0] wr_data;
wire wr_stb;
wire [10:0] reg_addr;
wire [10:0] locl_addr;
wire [31:0] locl_wr_data;
wire [31:0] spare;
wire [95:0] cceip0_out_ia_wdata;
wire [12:0] cceip0_out_ia_config;
wire [95:0] cceip0_out_ia_rdata;
wire [16:0] cceip0_out_ia_status;
wire [19:0] cceip0_out_ia_capability;
wire [11:0] cceip0_out_im_status;
wire [11:0] cceip0_out_im_config;
wire [95:0] cddip0_out_ia_wdata;
wire [12:0] cddip0_out_ia_config;
wire [95:0] cddip0_out_ia_rdata;
wire [16:0] cddip0_out_ia_status;
wire [19:0] cddip0_out_ia_capability;
wire [11:0] cddip0_out_im_status;
wire [11:0] cddip0_out_im_config;
wire [95:0] cceip1_out_ia_wdata;
wire [12:0] cceip1_out_ia_config;
wire [95:0] cceip1_out_ia_rdata;
wire [16:0] cceip1_out_ia_status;
wire [19:0] cceip1_out_ia_capability;
wire [11:0] cceip1_out_im_status;
wire [11:0] cceip1_out_im_config;
wire [95:0] cddip1_out_ia_wdata;
wire [12:0] cddip1_out_ia_config;
wire [95:0] cddip1_out_ia_rdata;
wire [16:0] cddip1_out_ia_status;
wire [19:0] cddip1_out_ia_capability;
wire [11:0] cddip1_out_im_status;
wire [11:0] cddip1_out_im_config;
wire [95:0] cceip2_out_ia_wdata;
wire [12:0] cceip2_out_ia_config;
wire [95:0] cceip2_out_ia_rdata;
wire [16:0] cceip2_out_ia_status;
wire [19:0] cceip2_out_ia_capability;
wire [11:0] cceip2_out_im_status;
wire [11:0] cceip2_out_im_config;
wire [95:0] cddip2_out_ia_wdata;
wire [12:0] cddip2_out_ia_config;
wire [95:0] cddip2_out_ia_rdata;
wire [16:0] cddip2_out_ia_status;
wire [19:0] cddip2_out_ia_capability;
wire [11:0] cddip2_out_im_status;
wire [11:0] cddip2_out_im_config;
wire [95:0] cceip3_out_ia_wdata;
wire [12:0] cceip3_out_ia_config;
wire [95:0] cceip3_out_ia_rdata;
wire [16:0] cceip3_out_ia_status;
wire [19:0] cceip3_out_ia_capability;
wire [11:0] cceip3_out_im_status;
wire [11:0] cceip3_out_im_config;
wire [95:0] cddip3_out_ia_wdata;
wire [12:0] cddip3_out_ia_config;
wire [95:0] cddip3_out_ia_rdata;
wire [16:0] cddip3_out_ia_status;
wire [19:0] cddip3_out_ia_capability;
wire [11:0] cddip3_out_im_status;
wire [11:0] cddip3_out_im_config;
wire [63:0] sa_snapshot_ia_wdata;
wire [63:0] sa_snapshot_ia_rdata;
wire [8:0] sa_snapshot_ia_config;
wire [12:0] sa_snapshot_ia_status;
wire [19:0] sa_snapshot_ia_capability;
wire [63:0] sa_count_ia_wdata;
wire [63:0] sa_count_ia_rdata;
wire [8:0] sa_count_ia_config;
wire [12:0] sa_count_ia_status;
wire [19:0] sa_count_ia_capability;
wire [31:0] sa_ctrl_ia_wdata;
wire [31:0] sa_ctrl_ia_rdata;
wire [8:0] sa_ctrl_ia_config;
wire [12:0] sa_ctrl_ia_status;
wire [19:0] sa_ctrl_ia_capability;
wire [95:0] cceip0_im_din;
wire cceip0_im_vld;
wire [95:0] cddip0_im_din;
wire cddip0_im_vld;
wire [95:0] cceip1_im_din;
wire cceip1_im_vld;
wire [95:0] cddip1_im_din;
wire cddip1_im_vld;
wire [95:0] cceip2_im_din;
wire cceip2_im_vld;
wire [95:0] cddip2_im_din;
wire cddip2_im_vld;
wire [95:0] cceip3_im_din;
wire cceip3_im_vld;
wire [95:0] cddip3_im_din;
wire cddip3_im_vld;
wire [15:0] im_available;
wire [1:0] im_consumed_kme_cceip0;
wire [1:0] im_available_kme_cceip0;
wire [1:0] im_consumed_kme_cddip0;
wire [1:0] im_available_kme_cddip0;
wire [1:0] im_consumed_kme_cceip1;
wire [1:0] im_available_kme_cceip1;
wire [1:0] im_consumed_kme_cddip1;
wire [1:0] im_available_kme_cddip1;
wire [1:0] im_consumed_kme_cceip2;
wire [1:0] im_available_kme_cceip2;
wire [1:0] im_consumed_kme_cddip2;
wire [1:0] im_available_kme_cddip2;
wire [1:0] im_consumed_kme_cceip3;
wire [1:0] im_available_kme_cceip3;
wire [1:0] im_consumed_kme_cddip3;
wire [1:0] im_available_kme_cddip3;
wire [82:0] kme_cceip0_ob_out_post;
wire [82:0] kme_cceip1_ob_out_post;
wire [82:0] kme_cceip2_ob_out_post;
wire [82:0] kme_cceip3_ob_out_post;
wire [82:0] kme_cddip0_ob_out_post;
wire [82:0] kme_cddip1_ob_out_post;
wire [82:0] kme_cddip2_ob_out_post;
wire [82:0] kme_cddip3_ob_out_post;
wire [31:0] blkid_revid_config;
wire [7:0] revid_wire;
supply1 n1;
supply0 n2;
wire [19:0] \ckv_ia_capability.r.part0 ;
wire [3:0] \ckv_ia_capability.f.mem_type ;
wire \ckv_ia_capability.f.ack_error ;
wire \ckv_ia_capability.f.sim_tmo ;
wire [3:0] \ckv_ia_capability.f.reserved_op ;
wire \ckv_ia_capability.f.compare ;
wire \ckv_ia_capability.f.set_init_start ;
wire \ckv_ia_capability.f.initialize_inc ;
wire \ckv_ia_capability.f.initialize ;
wire \ckv_ia_capability.f.reset ;
wire \ckv_ia_capability.f.disabled ;
wire \ckv_ia_capability.f.enable ;
wire \ckv_ia_capability.f.write ;
wire \ckv_ia_capability.f.read ;
wire \ckv_ia_capability.f.nop ;
wire [22:0] \ckv_ia_status.r.part0 ;
wire [2:0] \ckv_ia_status.f.code ;
wire [4:0] \ckv_ia_status.f.datawords ;
wire [14:0] \ckv_ia_status.f.addr ;
wire [19:0] \kim_ia_capability.r.part0 ;
wire [3:0] \kim_ia_capability.f.mem_type ;
wire \kim_ia_capability.f.ack_error ;
wire \kim_ia_capability.f.sim_tmo ;
wire [3:0] \kim_ia_capability.f.reserved_op ;
wire \kim_ia_capability.f.compare ;
wire \kim_ia_capability.f.set_init_start ;
wire \kim_ia_capability.f.initialize_inc ;
wire \kim_ia_capability.f.initialize ;
wire \kim_ia_capability.f.reset ;
wire \kim_ia_capability.f.disabled ;
wire \kim_ia_capability.f.enable ;
wire \kim_ia_capability.f.write ;
wire \kim_ia_capability.f.read ;
wire \kim_ia_capability.f.nop ;
wire [21:0] \kim_ia_status.r.part0 ;
wire [2:0] \kim_ia_status.f.code ;
wire [4:0] \kim_ia_status.f.datawords ;
wire [13:0] \kim_ia_status.f.addr ;
wire [31:0] \spare.r.part0 ;
wire [31:0] \spare.f.spare ;
wire [31:0] \cceip0_out_ia_wdata.r.part2 ;
wire [31:0] \cceip0_out_ia_wdata.r.part1 ;
wire [31:0] \cceip0_out_ia_wdata.r.part0 ;
wire [31:0] \cceip0_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cceip0_out_ia_wdata.f.tdata_lo ;
wire \cceip0_out_ia_wdata.f.eob ;
wire [7:0] \cceip0_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cceip0_out_ia_wdata.f.unused1 ;
wire \cceip0_out_ia_wdata.f.tid ;
wire [7:0] \cceip0_out_ia_wdata.f.tuser ;
wire [5:0] \cceip0_out_ia_wdata.f.unused0 ;
wire [12:0] \cceip0_out_ia_config.r.part0 ;
wire [3:0] \cceip0_out_ia_config.f.op ;
wire [8:0] \cceip0_out_ia_config.f.addr ;
wire [31:0] \cceip0_out_ia_rdata.r.part2 ;
wire [31:0] \cceip0_out_ia_rdata.r.part1 ;
wire [31:0] \cceip0_out_ia_rdata.r.part0 ;
wire [31:0] \cceip0_out_ia_rdata.f.tdata_hi ;
wire [31:0] \cceip0_out_ia_rdata.f.tdata_lo ;
wire \cceip0_out_ia_rdata.f.eob ;
wire [7:0] \cceip0_out_ia_rdata.f.bytes_vld ;
wire [7:0] \cceip0_out_ia_rdata.f.unused1 ;
wire \cceip0_out_ia_rdata.f.tid ;
wire [7:0] \cceip0_out_ia_rdata.f.tuser ;
wire [5:0] \cceip0_out_ia_rdata.f.unused0 ;
wire [16:0] \cceip0_out_ia_status.r.part0 ;
wire [2:0] \cceip0_out_ia_status.f.code ;
wire [4:0] \cceip0_out_ia_status.f.datawords ;
wire [8:0] \cceip0_out_ia_status.f.addr ;
wire [19:0] \cceip0_out_ia_capability.r.part0 ;
wire [3:0] \cceip0_out_ia_capability.f.mem_type ;
wire \cceip0_out_ia_capability.f.ack_error ;
wire \cceip0_out_ia_capability.f.sim_tmo ;
wire [3:0] \cceip0_out_ia_capability.f.reserved_op ;
wire \cceip0_out_ia_capability.f.compare ;
wire \cceip0_out_ia_capability.f.set_init_start ;
wire \cceip0_out_ia_capability.f.initialize_inc ;
wire \cceip0_out_ia_capability.f.initialize ;
wire \cceip0_out_ia_capability.f.reset ;
wire \cceip0_out_ia_capability.f.disabled ;
wire \cceip0_out_ia_capability.f.enable ;
wire \cceip0_out_ia_capability.f.write ;
wire \cceip0_out_ia_capability.f.read ;
wire \cceip0_out_ia_capability.f.nop ;
wire [11:0] \cceip0_out_im_status.r.part0 ;
wire \cceip0_out_im_status.f.bank_hi ;
wire \cceip0_out_im_status.f.bank_lo ;
wire \cceip0_out_im_status.f.overflow ;
wire [8:0] \cceip0_out_im_status.f.wr_pointer ;
wire [11:0] \cceip0_out_im_config.r.part0 ;
wire [1:0] \cceip0_out_im_config.f.mode ;
wire [9:0] \cceip0_out_im_config.f.wr_credit_config ;
wire [31:0] \cddip0_out_ia_wdata.r.part2 ;
wire [31:0] \cddip0_out_ia_wdata.r.part1 ;
wire [31:0] \cddip0_out_ia_wdata.r.part0 ;
wire [31:0] \cddip0_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cddip0_out_ia_wdata.f.tdata_lo ;
wire \cddip0_out_ia_wdata.f.eob ;
wire [7:0] \cddip0_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cddip0_out_ia_wdata.f.unused1 ;
wire \cddip0_out_ia_wdata.f.tid ;
wire [7:0] \cddip0_out_ia_wdata.f.tuser ;
wire [5:0] \cddip0_out_ia_wdata.f.unused0 ;
wire [12:0] \cddip0_out_ia_config.r.part0 ;
wire [3:0] \cddip0_out_ia_config.f.op ;
wire [8:0] \cddip0_out_ia_config.f.addr ;
wire [31:0] \cddip0_out_ia_rdata.r.part2 ;
wire [31:0] \cddip0_out_ia_rdata.r.part1 ;
wire [31:0] \cddip0_out_ia_rdata.r.part0 ;
wire [31:0] \cddip0_out_ia_rdata.f.tdata_hi ;
wire [31:0] \cddip0_out_ia_rdata.f.tdata_lo ;
wire \cddip0_out_ia_rdata.f.eob ;
wire [7:0] \cddip0_out_ia_rdata.f.bytes_vld ;
wire [7:0] \cddip0_out_ia_rdata.f.unused1 ;
wire \cddip0_out_ia_rdata.f.tid ;
wire [7:0] \cddip0_out_ia_rdata.f.tuser ;
wire [5:0] \cddip0_out_ia_rdata.f.unused0 ;
wire [16:0] \cddip0_out_ia_status.r.part0 ;
wire [2:0] \cddip0_out_ia_status.f.code ;
wire [4:0] \cddip0_out_ia_status.f.datawords ;
wire [8:0] \cddip0_out_ia_status.f.addr ;
wire [19:0] \cddip0_out_ia_capability.r.part0 ;
wire [3:0] \cddip0_out_ia_capability.f.mem_type ;
wire \cddip0_out_ia_capability.f.ack_error ;
wire \cddip0_out_ia_capability.f.sim_tmo ;
wire [3:0] \cddip0_out_ia_capability.f.reserved_op ;
wire \cddip0_out_ia_capability.f.compare ;
wire \cddip0_out_ia_capability.f.set_init_start ;
wire \cddip0_out_ia_capability.f.initialize_inc ;
wire \cddip0_out_ia_capability.f.initialize ;
wire \cddip0_out_ia_capability.f.reset ;
wire \cddip0_out_ia_capability.f.disabled ;
wire \cddip0_out_ia_capability.f.enable ;
wire \cddip0_out_ia_capability.f.write ;
wire \cddip0_out_ia_capability.f.read ;
wire \cddip0_out_ia_capability.f.nop ;
wire [11:0] \cddip0_out_im_status.r.part0 ;
wire \cddip0_out_im_status.f.bank_hi ;
wire \cddip0_out_im_status.f.bank_lo ;
wire \cddip0_out_im_status.f.overflow ;
wire [8:0] \cddip0_out_im_status.f.wr_pointer ;
wire [11:0] \cddip0_out_im_config.r.part0 ;
wire [1:0] \cddip0_out_im_config.f.mode ;
wire [9:0] \cddip0_out_im_config.f.wr_credit_config ;
wire [31:0] \cceip1_out_ia_wdata.r.part2 ;
wire [31:0] \cceip1_out_ia_wdata.r.part1 ;
wire [31:0] \cceip1_out_ia_wdata.r.part0 ;
wire [31:0] \cceip1_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cceip1_out_ia_wdata.f.tdata_lo ;
wire \cceip1_out_ia_wdata.f.eob ;
wire [7:0] \cceip1_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cceip1_out_ia_wdata.f.unused1 ;
wire \cceip1_out_ia_wdata.f.tid ;
wire [7:0] \cceip1_out_ia_wdata.f.tuser ;
wire [5:0] \cceip1_out_ia_wdata.f.unused0 ;
wire [12:0] \cceip1_out_ia_config.r.part0 ;
wire [3:0] \cceip1_out_ia_config.f.op ;
wire [8:0] \cceip1_out_ia_config.f.addr ;
wire [31:0] \cceip1_out_ia_rdata.r.part2 ;
wire [31:0] \cceip1_out_ia_rdata.r.part1 ;
wire [31:0] \cceip1_out_ia_rdata.r.part0 ;
wire [31:0] \cceip1_out_ia_rdata.f.tdata_hi ;
wire [31:0] \cceip1_out_ia_rdata.f.tdata_lo ;
wire \cceip1_out_ia_rdata.f.eob ;
wire [7:0] \cceip1_out_ia_rdata.f.bytes_vld ;
wire [7:0] \cceip1_out_ia_rdata.f.unused1 ;
wire \cceip1_out_ia_rdata.f.tid ;
wire [7:0] \cceip1_out_ia_rdata.f.tuser ;
wire [5:0] \cceip1_out_ia_rdata.f.unused0 ;
wire [16:0] \cceip1_out_ia_status.r.part0 ;
wire [2:0] \cceip1_out_ia_status.f.code ;
wire [4:0] \cceip1_out_ia_status.f.datawords ;
wire [8:0] \cceip1_out_ia_status.f.addr ;
wire [19:0] \cceip1_out_ia_capability.r.part0 ;
wire [3:0] \cceip1_out_ia_capability.f.mem_type ;
wire \cceip1_out_ia_capability.f.ack_error ;
wire \cceip1_out_ia_capability.f.sim_tmo ;
wire [3:0] \cceip1_out_ia_capability.f.reserved_op ;
wire \cceip1_out_ia_capability.f.compare ;
wire \cceip1_out_ia_capability.f.set_init_start ;
wire \cceip1_out_ia_capability.f.initialize_inc ;
wire \cceip1_out_ia_capability.f.initialize ;
wire \cceip1_out_ia_capability.f.reset ;
wire \cceip1_out_ia_capability.f.disabled ;
wire \cceip1_out_ia_capability.f.enable ;
wire \cceip1_out_ia_capability.f.write ;
wire \cceip1_out_ia_capability.f.read ;
wire \cceip1_out_ia_capability.f.nop ;
wire [11:0] \cceip1_out_im_status.r.part0 ;
wire \cceip1_out_im_status.f.bank_hi ;
wire \cceip1_out_im_status.f.bank_lo ;
wire \cceip1_out_im_status.f.overflow ;
wire [8:0] \cceip1_out_im_status.f.wr_pointer ;
wire [11:0] \cceip1_out_im_config.r.part0 ;
wire [1:0] \cceip1_out_im_config.f.mode ;
wire [9:0] \cceip1_out_im_config.f.wr_credit_config ;
wire [31:0] \cddip1_out_ia_wdata.r.part2 ;
wire [31:0] \cddip1_out_ia_wdata.r.part1 ;
wire [31:0] \cddip1_out_ia_wdata.r.part0 ;
wire [31:0] \cddip1_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cddip1_out_ia_wdata.f.tdata_lo ;
wire \cddip1_out_ia_wdata.f.eob ;
wire [7:0] \cddip1_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cddip1_out_ia_wdata.f.unused1 ;
wire \cddip1_out_ia_wdata.f.tid ;
wire [7:0] \cddip1_out_ia_wdata.f.tuser ;
wire [5:0] \cddip1_out_ia_wdata.f.unused0 ;
wire [12:0] \cddip1_out_ia_config.r.part0 ;
wire [3:0] \cddip1_out_ia_config.f.op ;
wire [8:0] \cddip1_out_ia_config.f.addr ;
wire [31:0] \cddip1_out_ia_rdata.r.part2 ;
wire [31:0] \cddip1_out_ia_rdata.r.part1 ;
wire [31:0] \cddip1_out_ia_rdata.r.part0 ;
wire [31:0] \cddip1_out_ia_rdata.f.tdata_hi ;
wire [31:0] \cddip1_out_ia_rdata.f.tdata_lo ;
wire \cddip1_out_ia_rdata.f.eob ;
wire [7:0] \cddip1_out_ia_rdata.f.bytes_vld ;
wire [7:0] \cddip1_out_ia_rdata.f.unused1 ;
wire \cddip1_out_ia_rdata.f.tid ;
wire [7:0] \cddip1_out_ia_rdata.f.tuser ;
wire [5:0] \cddip1_out_ia_rdata.f.unused0 ;
wire [16:0] \cddip1_out_ia_status.r.part0 ;
wire [2:0] \cddip1_out_ia_status.f.code ;
wire [4:0] \cddip1_out_ia_status.f.datawords ;
wire [8:0] \cddip1_out_ia_status.f.addr ;
wire [19:0] \cddip1_out_ia_capability.r.part0 ;
wire [3:0] \cddip1_out_ia_capability.f.mem_type ;
wire \cddip1_out_ia_capability.f.ack_error ;
wire \cddip1_out_ia_capability.f.sim_tmo ;
wire [3:0] \cddip1_out_ia_capability.f.reserved_op ;
wire \cddip1_out_ia_capability.f.compare ;
wire \cddip1_out_ia_capability.f.set_init_start ;
wire \cddip1_out_ia_capability.f.initialize_inc ;
wire \cddip1_out_ia_capability.f.initialize ;
wire \cddip1_out_ia_capability.f.reset ;
wire \cddip1_out_ia_capability.f.disabled ;
wire \cddip1_out_ia_capability.f.enable ;
wire \cddip1_out_ia_capability.f.write ;
wire \cddip1_out_ia_capability.f.read ;
wire \cddip1_out_ia_capability.f.nop ;
wire [11:0] \cddip1_out_im_status.r.part0 ;
wire \cddip1_out_im_status.f.bank_hi ;
wire \cddip1_out_im_status.f.bank_lo ;
wire \cddip1_out_im_status.f.overflow ;
wire [8:0] \cddip1_out_im_status.f.wr_pointer ;
wire [11:0] \cddip1_out_im_config.r.part0 ;
wire [1:0] \cddip1_out_im_config.f.mode ;
wire [9:0] \cddip1_out_im_config.f.wr_credit_config ;
wire [31:0] \cceip2_out_ia_wdata.r.part2 ;
wire [31:0] \cceip2_out_ia_wdata.r.part1 ;
wire [31:0] \cceip2_out_ia_wdata.r.part0 ;
wire [31:0] \cceip2_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cceip2_out_ia_wdata.f.tdata_lo ;
wire \cceip2_out_ia_wdata.f.eob ;
wire [7:0] \cceip2_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cceip2_out_ia_wdata.f.unused1 ;
wire \cceip2_out_ia_wdata.f.tid ;
wire [7:0] \cceip2_out_ia_wdata.f.tuser ;
wire [5:0] \cceip2_out_ia_wdata.f.unused0 ;
wire [12:0] \cceip2_out_ia_config.r.part0 ;
wire [3:0] \cceip2_out_ia_config.f.op ;
wire [8:0] \cceip2_out_ia_config.f.addr ;
wire [31:0] \cceip2_out_ia_rdata.r.part2 ;
wire [31:0] \cceip2_out_ia_rdata.r.part1 ;
wire [31:0] \cceip2_out_ia_rdata.r.part0 ;
wire [31:0] \cceip2_out_ia_rdata.f.tdata_hi ;
wire [31:0] \cceip2_out_ia_rdata.f.tdata_lo ;
wire \cceip2_out_ia_rdata.f.eob ;
wire [7:0] \cceip2_out_ia_rdata.f.bytes_vld ;
wire [7:0] \cceip2_out_ia_rdata.f.unused1 ;
wire \cceip2_out_ia_rdata.f.tid ;
wire [7:0] \cceip2_out_ia_rdata.f.tuser ;
wire [5:0] \cceip2_out_ia_rdata.f.unused0 ;
wire [16:0] \cceip2_out_ia_status.r.part0 ;
wire [2:0] \cceip2_out_ia_status.f.code ;
wire [4:0] \cceip2_out_ia_status.f.datawords ;
wire [8:0] \cceip2_out_ia_status.f.addr ;
wire [19:0] \cceip2_out_ia_capability.r.part0 ;
wire [3:0] \cceip2_out_ia_capability.f.mem_type ;
wire \cceip2_out_ia_capability.f.ack_error ;
wire \cceip2_out_ia_capability.f.sim_tmo ;
wire [3:0] \cceip2_out_ia_capability.f.reserved_op ;
wire \cceip2_out_ia_capability.f.compare ;
wire \cceip2_out_ia_capability.f.set_init_start ;
wire \cceip2_out_ia_capability.f.initialize_inc ;
wire \cceip2_out_ia_capability.f.initialize ;
wire \cceip2_out_ia_capability.f.reset ;
wire \cceip2_out_ia_capability.f.disabled ;
wire \cceip2_out_ia_capability.f.enable ;
wire \cceip2_out_ia_capability.f.write ;
wire \cceip2_out_ia_capability.f.read ;
wire \cceip2_out_ia_capability.f.nop ;
wire [11:0] \cceip2_out_im_status.r.part0 ;
wire \cceip2_out_im_status.f.bank_hi ;
wire \cceip2_out_im_status.f.bank_lo ;
wire \cceip2_out_im_status.f.overflow ;
wire [8:0] \cceip2_out_im_status.f.wr_pointer ;
wire [11:0] \cceip2_out_im_config.r.part0 ;
wire [1:0] \cceip2_out_im_config.f.mode ;
wire [9:0] \cceip2_out_im_config.f.wr_credit_config ;
wire [31:0] \cddip2_out_ia_wdata.r.part2 ;
wire [31:0] \cddip2_out_ia_wdata.r.part1 ;
wire [31:0] \cddip2_out_ia_wdata.r.part0 ;
wire [31:0] \cddip2_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cddip2_out_ia_wdata.f.tdata_lo ;
wire \cddip2_out_ia_wdata.f.eob ;
wire [7:0] \cddip2_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cddip2_out_ia_wdata.f.unused1 ;
wire \cddip2_out_ia_wdata.f.tid ;
wire [7:0] \cddip2_out_ia_wdata.f.tuser ;
wire [5:0] \cddip2_out_ia_wdata.f.unused0 ;
wire [12:0] \cddip2_out_ia_config.r.part0 ;
wire [3:0] \cddip2_out_ia_config.f.op ;
wire [8:0] \cddip2_out_ia_config.f.addr ;
wire [31:0] \cddip2_out_ia_rdata.r.part2 ;
wire [31:0] \cddip2_out_ia_rdata.r.part1 ;
wire [31:0] \cddip2_out_ia_rdata.r.part0 ;
wire [31:0] \cddip2_out_ia_rdata.f.tdata_hi ;
wire [31:0] \cddip2_out_ia_rdata.f.tdata_lo ;
wire \cddip2_out_ia_rdata.f.eob ;
wire [7:0] \cddip2_out_ia_rdata.f.bytes_vld ;
wire [7:0] \cddip2_out_ia_rdata.f.unused1 ;
wire \cddip2_out_ia_rdata.f.tid ;
wire [7:0] \cddip2_out_ia_rdata.f.tuser ;
wire [5:0] \cddip2_out_ia_rdata.f.unused0 ;
wire [16:0] \cddip2_out_ia_status.r.part0 ;
wire [2:0] \cddip2_out_ia_status.f.code ;
wire [4:0] \cddip2_out_ia_status.f.datawords ;
wire [8:0] \cddip2_out_ia_status.f.addr ;
wire [19:0] \cddip2_out_ia_capability.r.part0 ;
wire [3:0] \cddip2_out_ia_capability.f.mem_type ;
wire \cddip2_out_ia_capability.f.ack_error ;
wire \cddip2_out_ia_capability.f.sim_tmo ;
wire [3:0] \cddip2_out_ia_capability.f.reserved_op ;
wire \cddip2_out_ia_capability.f.compare ;
wire \cddip2_out_ia_capability.f.set_init_start ;
wire \cddip2_out_ia_capability.f.initialize_inc ;
wire \cddip2_out_ia_capability.f.initialize ;
wire \cddip2_out_ia_capability.f.reset ;
wire \cddip2_out_ia_capability.f.disabled ;
wire \cddip2_out_ia_capability.f.enable ;
wire \cddip2_out_ia_capability.f.write ;
wire \cddip2_out_ia_capability.f.read ;
wire \cddip2_out_ia_capability.f.nop ;
wire [11:0] \cddip2_out_im_status.r.part0 ;
wire \cddip2_out_im_status.f.bank_hi ;
wire \cddip2_out_im_status.f.bank_lo ;
wire \cddip2_out_im_status.f.overflow ;
wire [8:0] \cddip2_out_im_status.f.wr_pointer ;
wire [11:0] \cddip2_out_im_config.r.part0 ;
wire [1:0] \cddip2_out_im_config.f.mode ;
wire [9:0] \cddip2_out_im_config.f.wr_credit_config ;
wire [31:0] \cceip3_out_ia_wdata.r.part2 ;
wire [31:0] \cceip3_out_ia_wdata.r.part1 ;
wire [31:0] \cceip3_out_ia_wdata.r.part0 ;
wire [31:0] \cceip3_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cceip3_out_ia_wdata.f.tdata_lo ;
wire \cceip3_out_ia_wdata.f.eob ;
wire [7:0] \cceip3_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cceip3_out_ia_wdata.f.unused1 ;
wire \cceip3_out_ia_wdata.f.tid ;
wire [7:0] \cceip3_out_ia_wdata.f.tuser ;
wire [5:0] \cceip3_out_ia_wdata.f.unused0 ;
wire [12:0] \cceip3_out_ia_config.r.part0 ;
wire [3:0] \cceip3_out_ia_config.f.op ;
wire [8:0] \cceip3_out_ia_config.f.addr ;
wire [31:0] \cceip3_out_ia_rdata.r.part2 ;
wire [31:0] \cceip3_out_ia_rdata.r.part1 ;
wire [31:0] \cceip3_out_ia_rdata.r.part0 ;
wire [31:0] \cceip3_out_ia_rdata.f.tdata_hi ;
wire [31:0] \cceip3_out_ia_rdata.f.tdata_lo ;
wire \cceip3_out_ia_rdata.f.eob ;
wire [7:0] \cceip3_out_ia_rdata.f.bytes_vld ;
wire [7:0] \cceip3_out_ia_rdata.f.unused1 ;
wire \cceip3_out_ia_rdata.f.tid ;
wire [7:0] \cceip3_out_ia_rdata.f.tuser ;
wire [5:0] \cceip3_out_ia_rdata.f.unused0 ;
wire [16:0] \cceip3_out_ia_status.r.part0 ;
wire [2:0] \cceip3_out_ia_status.f.code ;
wire [4:0] \cceip3_out_ia_status.f.datawords ;
wire [8:0] \cceip3_out_ia_status.f.addr ;
wire [19:0] \cceip3_out_ia_capability.r.part0 ;
wire [3:0] \cceip3_out_ia_capability.f.mem_type ;
wire \cceip3_out_ia_capability.f.ack_error ;
wire \cceip3_out_ia_capability.f.sim_tmo ;
wire [3:0] \cceip3_out_ia_capability.f.reserved_op ;
wire \cceip3_out_ia_capability.f.compare ;
wire \cceip3_out_ia_capability.f.set_init_start ;
wire \cceip3_out_ia_capability.f.initialize_inc ;
wire \cceip3_out_ia_capability.f.initialize ;
wire \cceip3_out_ia_capability.f.reset ;
wire \cceip3_out_ia_capability.f.disabled ;
wire \cceip3_out_ia_capability.f.enable ;
wire \cceip3_out_ia_capability.f.write ;
wire \cceip3_out_ia_capability.f.read ;
wire \cceip3_out_ia_capability.f.nop ;
wire [11:0] \cceip3_out_im_status.r.part0 ;
wire \cceip3_out_im_status.f.bank_hi ;
wire \cceip3_out_im_status.f.bank_lo ;
wire \cceip3_out_im_status.f.overflow ;
wire [8:0] \cceip3_out_im_status.f.wr_pointer ;
wire [11:0] \cceip3_out_im_config.r.part0 ;
wire [1:0] \cceip3_out_im_config.f.mode ;
wire [9:0] \cceip3_out_im_config.f.wr_credit_config ;
wire [31:0] \cddip3_out_ia_wdata.r.part2 ;
wire [31:0] \cddip3_out_ia_wdata.r.part1 ;
wire [31:0] \cddip3_out_ia_wdata.r.part0 ;
wire [31:0] \cddip3_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cddip3_out_ia_wdata.f.tdata_lo ;
wire \cddip3_out_ia_wdata.f.eob ;
wire [7:0] \cddip3_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cddip3_out_ia_wdata.f.unused1 ;
wire \cddip3_out_ia_wdata.f.tid ;
wire [7:0] \cddip3_out_ia_wdata.f.tuser ;
wire [5:0] \cddip3_out_ia_wdata.f.unused0 ;
wire [12:0] \cddip3_out_ia_config.r.part0 ;
wire [3:0] \cddip3_out_ia_config.f.op ;
wire [8:0] \cddip3_out_ia_config.f.addr ;
wire [31:0] \cddip3_out_ia_rdata.r.part2 ;
wire [31:0] \cddip3_out_ia_rdata.r.part1 ;
wire [31:0] \cddip3_out_ia_rdata.r.part0 ;
wire [31:0] \cddip3_out_ia_rdata.f.tdata_hi ;
wire [31:0] \cddip3_out_ia_rdata.f.tdata_lo ;
wire \cddip3_out_ia_rdata.f.eob ;
wire [7:0] \cddip3_out_ia_rdata.f.bytes_vld ;
wire [7:0] \cddip3_out_ia_rdata.f.unused1 ;
wire \cddip3_out_ia_rdata.f.tid ;
wire [7:0] \cddip3_out_ia_rdata.f.tuser ;
wire [5:0] \cddip3_out_ia_rdata.f.unused0 ;
wire [16:0] \cddip3_out_ia_status.r.part0 ;
wire [2:0] \cddip3_out_ia_status.f.code ;
wire [4:0] \cddip3_out_ia_status.f.datawords ;
wire [8:0] \cddip3_out_ia_status.f.addr ;
wire [19:0] \cddip3_out_ia_capability.r.part0 ;
wire [3:0] \cddip3_out_ia_capability.f.mem_type ;
wire \cddip3_out_ia_capability.f.ack_error ;
wire \cddip3_out_ia_capability.f.sim_tmo ;
wire [3:0] \cddip3_out_ia_capability.f.reserved_op ;
wire \cddip3_out_ia_capability.f.compare ;
wire \cddip3_out_ia_capability.f.set_init_start ;
wire \cddip3_out_ia_capability.f.initialize_inc ;
wire \cddip3_out_ia_capability.f.initialize ;
wire \cddip3_out_ia_capability.f.reset ;
wire \cddip3_out_ia_capability.f.disabled ;
wire \cddip3_out_ia_capability.f.enable ;
wire \cddip3_out_ia_capability.f.write ;
wire \cddip3_out_ia_capability.f.read ;
wire \cddip3_out_ia_capability.f.nop ;
wire [11:0] \cddip3_out_im_status.r.part0 ;
wire \cddip3_out_im_status.f.bank_hi ;
wire \cddip3_out_im_status.f.bank_lo ;
wire \cddip3_out_im_status.f.overflow ;
wire [8:0] \cddip3_out_im_status.f.wr_pointer ;
wire [11:0] \cddip3_out_im_config.r.part0 ;
wire [1:0] \cddip3_out_im_config.f.mode ;
wire [9:0] \cddip3_out_im_config.f.wr_credit_config ;
wire [31:0] \sa_snapshot_ia_wdata.r.part1 ;
wire [31:0] \sa_snapshot_ia_wdata.r.part0 ;
wire [13:0] \sa_snapshot_ia_wdata.f.unused ;
wire [17:0] \sa_snapshot_ia_wdata.f.upper ;
wire [31:0] \sa_snapshot_ia_wdata.f.lower ;
wire [31:0] \sa_snapshot_ia_rdata.r.part1 ;
wire [31:0] \sa_snapshot_ia_rdata.r.part0 ;
wire [13:0] \sa_snapshot_ia_rdata.f.unused ;
wire [17:0] \sa_snapshot_ia_rdata.f.upper ;
wire [31:0] \sa_snapshot_ia_rdata.f.lower ;
wire [8:0] \sa_snapshot_ia_config.r.part0 ;
wire [3:0] \sa_snapshot_ia_config.f.op ;
wire [4:0] \sa_snapshot_ia_config.f.addr ;
wire [12:0] \sa_snapshot_ia_status.r.part0 ;
wire [2:0] \sa_snapshot_ia_status.f.code ;
wire [4:0] \sa_snapshot_ia_status.f.datawords ;
wire [4:0] \sa_snapshot_ia_status.f.addr ;
wire [19:0] \sa_snapshot_ia_capability.r.part0 ;
wire [3:0] \sa_snapshot_ia_capability.f.mem_type ;
wire \sa_snapshot_ia_capability.f.ack_error ;
wire \sa_snapshot_ia_capability.f.sim_tmo ;
wire [3:0] \sa_snapshot_ia_capability.f.reserved_op ;
wire \sa_snapshot_ia_capability.f.compare ;
wire \sa_snapshot_ia_capability.f.set_init_start ;
wire \sa_snapshot_ia_capability.f.initialize_inc ;
wire \sa_snapshot_ia_capability.f.initialize ;
wire \sa_snapshot_ia_capability.f.reset ;
wire \sa_snapshot_ia_capability.f.disabled ;
wire \sa_snapshot_ia_capability.f.enable ;
wire \sa_snapshot_ia_capability.f.write ;
wire \sa_snapshot_ia_capability.f.read ;
wire \sa_snapshot_ia_capability.f.nop ;
wire [31:0] \sa_count_ia_wdata.r.part1 ;
wire [31:0] \sa_count_ia_wdata.r.part0 ;
wire [13:0] \sa_count_ia_wdata.f.unused ;
wire [17:0] \sa_count_ia_wdata.f.upper ;
wire [31:0] \sa_count_ia_wdata.f.lower ;
wire [31:0] \sa_count_ia_rdata.r.part1 ;
wire [31:0] \sa_count_ia_rdata.r.part0 ;
wire [13:0] \sa_count_ia_rdata.f.unused ;
wire [17:0] \sa_count_ia_rdata.f.upper ;
wire [31:0] \sa_count_ia_rdata.f.lower ;
wire [8:0] \sa_count_ia_config.r.part0 ;
wire [3:0] \sa_count_ia_config.f.op ;
wire [4:0] \sa_count_ia_config.f.addr ;
wire [12:0] \sa_count_ia_status.r.part0 ;
wire [2:0] \sa_count_ia_status.f.code ;
wire [4:0] \sa_count_ia_status.f.datawords ;
wire [4:0] \sa_count_ia_status.f.addr ;
wire [19:0] \sa_count_ia_capability.r.part0 ;
wire [3:0] \sa_count_ia_capability.f.mem_type ;
wire \sa_count_ia_capability.f.ack_error ;
wire \sa_count_ia_capability.f.sim_tmo ;
wire [3:0] \sa_count_ia_capability.f.reserved_op ;
wire \sa_count_ia_capability.f.compare ;
wire \sa_count_ia_capability.f.set_init_start ;
wire \sa_count_ia_capability.f.initialize_inc ;
wire \sa_count_ia_capability.f.initialize ;
wire \sa_count_ia_capability.f.reset ;
wire \sa_count_ia_capability.f.disabled ;
wire \sa_count_ia_capability.f.enable ;
wire \sa_count_ia_capability.f.write ;
wire \sa_count_ia_capability.f.read ;
wire \sa_count_ia_capability.f.nop ;
wire [31:0] \sa_ctrl_ia_wdata.r.part0 ;
wire [26:0] \sa_ctrl_ia_wdata.f.spare ;
wire [4:0] \sa_ctrl_ia_wdata.f.sa_event_sel ;
wire [31:0] \sa_ctrl_ia_rdata.r.part0 ;
wire [26:0] \sa_ctrl_ia_rdata.f.spare ;
wire [4:0] \sa_ctrl_ia_rdata.f.sa_event_sel ;
wire [8:0] \sa_ctrl_ia_config.r.part0 ;
wire [3:0] \sa_ctrl_ia_config.f.op ;
wire [4:0] \sa_ctrl_ia_config.f.addr ;
wire [12:0] \sa_ctrl_ia_status.r.part0 ;
wire [2:0] \sa_ctrl_ia_status.f.code ;
wire [4:0] \sa_ctrl_ia_status.f.datawords ;
wire [4:0] \sa_ctrl_ia_status.f.addr ;
wire [19:0] \sa_ctrl_ia_capability.r.part0 ;
wire [3:0] \sa_ctrl_ia_capability.f.mem_type ;
wire \sa_ctrl_ia_capability.f.ack_error ;
wire \sa_ctrl_ia_capability.f.sim_tmo ;
wire [3:0] \sa_ctrl_ia_capability.f.reserved_op ;
wire \sa_ctrl_ia_capability.f.compare ;
wire \sa_ctrl_ia_capability.f.set_init_start ;
wire \sa_ctrl_ia_capability.f.initialize_inc ;
wire \sa_ctrl_ia_capability.f.initialize ;
wire \sa_ctrl_ia_capability.f.reset ;
wire \sa_ctrl_ia_capability.f.disabled ;
wire \sa_ctrl_ia_capability.f.enable ;
wire \sa_ctrl_ia_capability.f.write ;
wire \sa_ctrl_ia_capability.f.read ;
wire \sa_ctrl_ia_capability.f.nop ;
wire [63:0] \cceip0_im_din.data.data ;
wire \cceip0_im_din.desc.eob ;
wire [7:0] \cceip0_im_din.desc.bytes_vld ;
wire [22:0] \cceip0_im_din.desc.im_meta ;
wire [63:0] \cddip0_im_din.data.data ;
wire \cddip0_im_din.desc.eob ;
wire [7:0] \cddip0_im_din.desc.bytes_vld ;
wire [22:0] \cddip0_im_din.desc.im_meta ;
wire [63:0] \cceip1_im_din.data.data ;
wire \cceip1_im_din.desc.eob ;
wire [7:0] \cceip1_im_din.desc.bytes_vld ;
wire [22:0] \cceip1_im_din.desc.im_meta ;
wire [63:0] \cddip1_im_din.data.data ;
wire \cddip1_im_din.desc.eob ;
wire [7:0] \cddip1_im_din.desc.bytes_vld ;
wire [22:0] \cddip1_im_din.desc.im_meta ;
wire [63:0] \cceip2_im_din.data.data ;
wire \cceip2_im_din.desc.eob ;
wire [7:0] \cceip2_im_din.desc.bytes_vld ;
wire [22:0] \cceip2_im_din.desc.im_meta ;
wire [63:0] \cddip2_im_din.data.data ;
wire \cddip2_im_din.desc.eob ;
wire [7:0] \cddip2_im_din.desc.bytes_vld ;
wire [22:0] \cddip2_im_din.desc.im_meta ;
wire [63:0] \cceip3_im_din.data.data ;
wire \cceip3_im_din.desc.eob ;
wire [7:0] \cceip3_im_din.desc.bytes_vld ;
wire [22:0] \cceip3_im_din.desc.im_meta ;
wire [63:0] \cddip3_im_din.data.data ;
wire \cddip3_im_din.desc.eob ;
wire [7:0] \cddip3_im_din.desc.bytes_vld ;
wire [22:0] \cddip3_im_din.desc.im_meta ;
wire \im_consumed_kme_cceip0.bank_hi ;
wire \im_consumed_kme_cceip0.bank_lo ;
wire \im_available_kme_cceip0.bank_hi ;
wire \im_available_kme_cceip0.bank_lo ;
wire \im_consumed_kme_cddip0.bank_hi ;
wire \im_consumed_kme_cddip0.bank_lo ;
wire \im_available_kme_cddip0.bank_hi ;
wire \im_available_kme_cddip0.bank_lo ;
wire \im_consumed_kme_cceip1.bank_hi ;
wire \im_consumed_kme_cceip1.bank_lo ;
wire \im_available_kme_cceip1.bank_hi ;
wire \im_available_kme_cceip1.bank_lo ;
wire \im_consumed_kme_cddip1.bank_hi ;
wire \im_consumed_kme_cddip1.bank_lo ;
wire \im_available_kme_cddip1.bank_hi ;
wire \im_available_kme_cddip1.bank_lo ;
wire \im_consumed_kme_cceip2.bank_hi ;
wire \im_consumed_kme_cceip2.bank_lo ;
wire \im_available_kme_cceip2.bank_hi ;
wire \im_available_kme_cceip2.bank_lo ;
wire \im_consumed_kme_cddip2.bank_hi ;
wire \im_consumed_kme_cddip2.bank_lo ;
wire \im_available_kme_cddip2.bank_hi ;
wire \im_available_kme_cddip2.bank_lo ;
wire \im_consumed_kme_cceip3.bank_hi ;
wire \im_consumed_kme_cceip3.bank_lo ;
wire \im_available_kme_cceip3.bank_hi ;
wire \im_available_kme_cceip3.bank_lo ;
wire \im_consumed_kme_cddip3.bank_hi ;
wire \im_consumed_kme_cddip3.bank_lo ;
wire \im_available_kme_cddip3.bank_hi ;
wire \im_available_kme_cddip3.bank_lo ;
wire \kme_cceip0_ob_out_post.tvalid ;
wire \kme_cceip0_ob_out_post.tlast ;
wire [0:0] \kme_cceip0_ob_out_post.tid ;
wire [7:0] \kme_cceip0_ob_out_post.tstrb ;
wire [7:0] \kme_cceip0_ob_out_post.tuser ;
wire [63:0] \kme_cceip0_ob_out_post.tdata ;
wire \kme_cceip1_ob_out_post.tvalid ;
wire \kme_cceip1_ob_out_post.tlast ;
wire [0:0] \kme_cceip1_ob_out_post.tid ;
wire [7:0] \kme_cceip1_ob_out_post.tstrb ;
wire [7:0] \kme_cceip1_ob_out_post.tuser ;
wire [63:0] \kme_cceip1_ob_out_post.tdata ;
wire \kme_cceip2_ob_out_post.tvalid ;
wire \kme_cceip2_ob_out_post.tlast ;
wire [0:0] \kme_cceip2_ob_out_post.tid ;
wire [7:0] \kme_cceip2_ob_out_post.tstrb ;
wire [7:0] \kme_cceip2_ob_out_post.tuser ;
wire [63:0] \kme_cceip2_ob_out_post.tdata ;
wire \kme_cceip3_ob_out_post.tvalid ;
wire \kme_cceip3_ob_out_post.tlast ;
wire [0:0] \kme_cceip3_ob_out_post.tid ;
wire [7:0] \kme_cceip3_ob_out_post.tstrb ;
wire [7:0] \kme_cceip3_ob_out_post.tuser ;
wire [63:0] \kme_cceip3_ob_out_post.tdata ;
wire \kme_cddip0_ob_out_post.tvalid ;
wire \kme_cddip0_ob_out_post.tlast ;
wire [0:0] \kme_cddip0_ob_out_post.tid ;
wire [7:0] \kme_cddip0_ob_out_post.tstrb ;
wire [7:0] \kme_cddip0_ob_out_post.tuser ;
wire [63:0] \kme_cddip0_ob_out_post.tdata ;
wire \kme_cddip1_ob_out_post.tvalid ;
wire \kme_cddip1_ob_out_post.tlast ;
wire [0:0] \kme_cddip1_ob_out_post.tid ;
wire [7:0] \kme_cddip1_ob_out_post.tstrb ;
wire [7:0] \kme_cddip1_ob_out_post.tuser ;
wire [63:0] \kme_cddip1_ob_out_post.tdata ;
wire \kme_cddip2_ob_out_post.tvalid ;
wire \kme_cddip2_ob_out_post.tlast ;
wire [0:0] \kme_cddip2_ob_out_post.tid ;
wire [7:0] \kme_cddip2_ob_out_post.tstrb ;
wire [7:0] \kme_cddip2_ob_out_post.tuser ;
wire [63:0] \kme_cddip2_ob_out_post.tdata ;
wire \kme_cddip3_ob_out_post.tvalid ;
wire \kme_cddip3_ob_out_post.tlast ;
wire [0:0] \kme_cddip3_ob_out_post.tid ;
wire [7:0] \kme_cddip3_ob_out_post.tstrb ;
wire [7:0] \kme_cddip3_ob_out_post.tuser ;
wire [63:0] \kme_cddip3_ob_out_post.tdata ;
wire [7:0] \revid_wire.r.part0 ;
wire [7:0] \revid_wire.f.revid ;
tran (rbus_ring_o[83], \rbus_ring_o.addr [15]);
tran (rbus_ring_o[82], \rbus_ring_o.addr [14]);
tran (rbus_ring_o[81], \rbus_ring_o.addr [13]);
tran (rbus_ring_o[80], \rbus_ring_o.addr [12]);
tran (rbus_ring_o[79], \rbus_ring_o.addr [11]);
tran (rbus_ring_o[78], \rbus_ring_o.addr [10]);
tran (rbus_ring_o[77], \rbus_ring_o.addr [9]);
tran (rbus_ring_o[76], \rbus_ring_o.addr [8]);
tran (rbus_ring_o[75], \rbus_ring_o.addr [7]);
tran (rbus_ring_o[74], \rbus_ring_o.addr [6]);
tran (rbus_ring_o[73], \rbus_ring_o.addr [5]);
tran (rbus_ring_o[72], \rbus_ring_o.addr [4]);
tran (rbus_ring_o[71], \rbus_ring_o.addr [3]);
tran (rbus_ring_o[70], \rbus_ring_o.addr [2]);
tran (rbus_ring_o[69], \rbus_ring_o.addr [1]);
tran (rbus_ring_o[68], \rbus_ring_o.addr [0]);
tran (rbus_ring_o[67], \rbus_ring_o.wr_strb );
tran (rbus_ring_o[66], \rbus_ring_o.wr_data [31]);
tran (rbus_ring_o[65], \rbus_ring_o.wr_data [30]);
tran (rbus_ring_o[64], \rbus_ring_o.wr_data [29]);
tran (rbus_ring_o[63], \rbus_ring_o.wr_data [28]);
tran (rbus_ring_o[62], \rbus_ring_o.wr_data [27]);
tran (rbus_ring_o[61], \rbus_ring_o.wr_data [26]);
tran (rbus_ring_o[60], \rbus_ring_o.wr_data [25]);
tran (rbus_ring_o[59], \rbus_ring_o.wr_data [24]);
tran (rbus_ring_o[58], \rbus_ring_o.wr_data [23]);
tran (rbus_ring_o[57], \rbus_ring_o.wr_data [22]);
tran (rbus_ring_o[56], \rbus_ring_o.wr_data [21]);
tran (rbus_ring_o[55], \rbus_ring_o.wr_data [20]);
tran (rbus_ring_o[54], \rbus_ring_o.wr_data [19]);
tran (rbus_ring_o[53], \rbus_ring_o.wr_data [18]);
tran (rbus_ring_o[52], \rbus_ring_o.wr_data [17]);
tran (rbus_ring_o[51], \rbus_ring_o.wr_data [16]);
tran (rbus_ring_o[50], \rbus_ring_o.wr_data [15]);
tran (rbus_ring_o[49], \rbus_ring_o.wr_data [14]);
tran (rbus_ring_o[48], \rbus_ring_o.wr_data [13]);
tran (rbus_ring_o[47], \rbus_ring_o.wr_data [12]);
tran (rbus_ring_o[46], \rbus_ring_o.wr_data [11]);
tran (rbus_ring_o[45], \rbus_ring_o.wr_data [10]);
tran (rbus_ring_o[44], \rbus_ring_o.wr_data [9]);
tran (rbus_ring_o[43], \rbus_ring_o.wr_data [8]);
tran (rbus_ring_o[42], \rbus_ring_o.wr_data [7]);
tran (rbus_ring_o[41], \rbus_ring_o.wr_data [6]);
tran (rbus_ring_o[40], \rbus_ring_o.wr_data [5]);
tran (rbus_ring_o[39], \rbus_ring_o.wr_data [4]);
tran (rbus_ring_o[38], \rbus_ring_o.wr_data [3]);
tran (rbus_ring_o[37], \rbus_ring_o.wr_data [2]);
tran (rbus_ring_o[36], \rbus_ring_o.wr_data [1]);
tran (rbus_ring_o[35], \rbus_ring_o.wr_data [0]);
tran (rbus_ring_o[34], \rbus_ring_o.rd_strb );
tran (rbus_ring_o[33], \rbus_ring_o.rd_data [31]);
tran (rbus_ring_o[32], \rbus_ring_o.rd_data [30]);
tran (rbus_ring_o[31], \rbus_ring_o.rd_data [29]);
tran (rbus_ring_o[30], \rbus_ring_o.rd_data [28]);
tran (rbus_ring_o[29], \rbus_ring_o.rd_data [27]);
tran (rbus_ring_o[28], \rbus_ring_o.rd_data [26]);
tran (rbus_ring_o[27], \rbus_ring_o.rd_data [25]);
tran (rbus_ring_o[26], \rbus_ring_o.rd_data [24]);
tran (rbus_ring_o[25], \rbus_ring_o.rd_data [23]);
tran (rbus_ring_o[24], \rbus_ring_o.rd_data [22]);
tran (rbus_ring_o[23], \rbus_ring_o.rd_data [21]);
tran (rbus_ring_o[22], \rbus_ring_o.rd_data [20]);
tran (rbus_ring_o[21], \rbus_ring_o.rd_data [19]);
tran (rbus_ring_o[20], \rbus_ring_o.rd_data [18]);
tran (rbus_ring_o[19], \rbus_ring_o.rd_data [17]);
tran (rbus_ring_o[18], \rbus_ring_o.rd_data [16]);
tran (rbus_ring_o[17], \rbus_ring_o.rd_data [15]);
tran (rbus_ring_o[16], \rbus_ring_o.rd_data [14]);
tran (rbus_ring_o[15], \rbus_ring_o.rd_data [13]);
tran (rbus_ring_o[14], \rbus_ring_o.rd_data [12]);
tran (rbus_ring_o[13], \rbus_ring_o.rd_data [11]);
tran (rbus_ring_o[12], \rbus_ring_o.rd_data [10]);
tran (rbus_ring_o[11], \rbus_ring_o.rd_data [9]);
tran (rbus_ring_o[10], \rbus_ring_o.rd_data [8]);
tran (rbus_ring_o[9], \rbus_ring_o.rd_data [7]);
tran (rbus_ring_o[8], \rbus_ring_o.rd_data [6]);
tran (rbus_ring_o[7], \rbus_ring_o.rd_data [5]);
tran (rbus_ring_o[6], \rbus_ring_o.rd_data [4]);
tran (rbus_ring_o[5], \rbus_ring_o.rd_data [3]);
tran (rbus_ring_o[4], \rbus_ring_o.rd_data [2]);
tran (rbus_ring_o[3], \rbus_ring_o.rd_data [1]);
tran (rbus_ring_o[2], \rbus_ring_o.rd_data [0]);
tran (rbus_ring_o[1], \rbus_ring_o.ack );
tran (rbus_ring_o[0], \rbus_ring_o.err_ack );
tran (kme_cceip0_ob_out[82], \kme_cceip0_ob_out.tvalid );
tran (kme_cceip0_ob_out[81], \kme_cceip0_ob_out.tlast );
tran (kme_cceip0_ob_out[80], \kme_cceip0_ob_out.tid [0]);
tran (kme_cceip0_ob_out[79], \kme_cceip0_ob_out.tstrb [7]);
tran (kme_cceip0_ob_out[78], \kme_cceip0_ob_out.tstrb [6]);
tran (kme_cceip0_ob_out[77], \kme_cceip0_ob_out.tstrb [5]);
tran (kme_cceip0_ob_out[76], \kme_cceip0_ob_out.tstrb [4]);
tran (kme_cceip0_ob_out[75], \kme_cceip0_ob_out.tstrb [3]);
tran (kme_cceip0_ob_out[74], \kme_cceip0_ob_out.tstrb [2]);
tran (kme_cceip0_ob_out[73], \kme_cceip0_ob_out.tstrb [1]);
tran (kme_cceip0_ob_out[72], \kme_cceip0_ob_out.tstrb [0]);
tran (kme_cceip0_ob_out[71], \kme_cceip0_ob_out.tuser [7]);
tran (kme_cceip0_ob_out[70], \kme_cceip0_ob_out.tuser [6]);
tran (kme_cceip0_ob_out[69], \kme_cceip0_ob_out.tuser [5]);
tran (kme_cceip0_ob_out[68], \kme_cceip0_ob_out.tuser [4]);
tran (kme_cceip0_ob_out[67], \kme_cceip0_ob_out.tuser [3]);
tran (kme_cceip0_ob_out[66], \kme_cceip0_ob_out.tuser [2]);
tran (kme_cceip0_ob_out[65], \kme_cceip0_ob_out.tuser [1]);
tran (kme_cceip0_ob_out[64], \kme_cceip0_ob_out.tuser [0]);
tran (kme_cceip0_ob_out[63], \kme_cceip0_ob_out.tdata [63]);
tran (kme_cceip0_ob_out[62], \kme_cceip0_ob_out.tdata [62]);
tran (kme_cceip0_ob_out[61], \kme_cceip0_ob_out.tdata [61]);
tran (kme_cceip0_ob_out[60], \kme_cceip0_ob_out.tdata [60]);
tran (kme_cceip0_ob_out[59], \kme_cceip0_ob_out.tdata [59]);
tran (kme_cceip0_ob_out[58], \kme_cceip0_ob_out.tdata [58]);
tran (kme_cceip0_ob_out[57], \kme_cceip0_ob_out.tdata [57]);
tran (kme_cceip0_ob_out[56], \kme_cceip0_ob_out.tdata [56]);
tran (kme_cceip0_ob_out[55], \kme_cceip0_ob_out.tdata [55]);
tran (kme_cceip0_ob_out[54], \kme_cceip0_ob_out.tdata [54]);
tran (kme_cceip0_ob_out[53], \kme_cceip0_ob_out.tdata [53]);
tran (kme_cceip0_ob_out[52], \kme_cceip0_ob_out.tdata [52]);
tran (kme_cceip0_ob_out[51], \kme_cceip0_ob_out.tdata [51]);
tran (kme_cceip0_ob_out[50], \kme_cceip0_ob_out.tdata [50]);
tran (kme_cceip0_ob_out[49], \kme_cceip0_ob_out.tdata [49]);
tran (kme_cceip0_ob_out[48], \kme_cceip0_ob_out.tdata [48]);
tran (kme_cceip0_ob_out[47], \kme_cceip0_ob_out.tdata [47]);
tran (kme_cceip0_ob_out[46], \kme_cceip0_ob_out.tdata [46]);
tran (kme_cceip0_ob_out[45], \kme_cceip0_ob_out.tdata [45]);
tran (kme_cceip0_ob_out[44], \kme_cceip0_ob_out.tdata [44]);
tran (kme_cceip0_ob_out[43], \kme_cceip0_ob_out.tdata [43]);
tran (kme_cceip0_ob_out[42], \kme_cceip0_ob_out.tdata [42]);
tran (kme_cceip0_ob_out[41], \kme_cceip0_ob_out.tdata [41]);
tran (kme_cceip0_ob_out[40], \kme_cceip0_ob_out.tdata [40]);
tran (kme_cceip0_ob_out[39], \kme_cceip0_ob_out.tdata [39]);
tran (kme_cceip0_ob_out[38], \kme_cceip0_ob_out.tdata [38]);
tran (kme_cceip0_ob_out[37], \kme_cceip0_ob_out.tdata [37]);
tran (kme_cceip0_ob_out[36], \kme_cceip0_ob_out.tdata [36]);
tran (kme_cceip0_ob_out[35], \kme_cceip0_ob_out.tdata [35]);
tran (kme_cceip0_ob_out[34], \kme_cceip0_ob_out.tdata [34]);
tran (kme_cceip0_ob_out[33], \kme_cceip0_ob_out.tdata [33]);
tran (kme_cceip0_ob_out[32], \kme_cceip0_ob_out.tdata [32]);
tran (kme_cceip0_ob_out[31], \kme_cceip0_ob_out.tdata [31]);
tran (kme_cceip0_ob_out[30], \kme_cceip0_ob_out.tdata [30]);
tran (kme_cceip0_ob_out[29], \kme_cceip0_ob_out.tdata [29]);
tran (kme_cceip0_ob_out[28], \kme_cceip0_ob_out.tdata [28]);
tran (kme_cceip0_ob_out[27], \kme_cceip0_ob_out.tdata [27]);
tran (kme_cceip0_ob_out[26], \kme_cceip0_ob_out.tdata [26]);
tran (kme_cceip0_ob_out[25], \kme_cceip0_ob_out.tdata [25]);
tran (kme_cceip0_ob_out[24], \kme_cceip0_ob_out.tdata [24]);
tran (kme_cceip0_ob_out[23], \kme_cceip0_ob_out.tdata [23]);
tran (kme_cceip0_ob_out[22], \kme_cceip0_ob_out.tdata [22]);
tran (kme_cceip0_ob_out[21], \kme_cceip0_ob_out.tdata [21]);
tran (kme_cceip0_ob_out[20], \kme_cceip0_ob_out.tdata [20]);
tran (kme_cceip0_ob_out[19], \kme_cceip0_ob_out.tdata [19]);
tran (kme_cceip0_ob_out[18], \kme_cceip0_ob_out.tdata [18]);
tran (kme_cceip0_ob_out[17], \kme_cceip0_ob_out.tdata [17]);
tran (kme_cceip0_ob_out[16], \kme_cceip0_ob_out.tdata [16]);
tran (kme_cceip0_ob_out[15], \kme_cceip0_ob_out.tdata [15]);
tran (kme_cceip0_ob_out[14], \kme_cceip0_ob_out.tdata [14]);
tran (kme_cceip0_ob_out[13], \kme_cceip0_ob_out.tdata [13]);
tran (kme_cceip0_ob_out[12], \kme_cceip0_ob_out.tdata [12]);
tran (kme_cceip0_ob_out[11], \kme_cceip0_ob_out.tdata [11]);
tran (kme_cceip0_ob_out[10], \kme_cceip0_ob_out.tdata [10]);
tran (kme_cceip0_ob_out[9], \kme_cceip0_ob_out.tdata [9]);
tran (kme_cceip0_ob_out[8], \kme_cceip0_ob_out.tdata [8]);
tran (kme_cceip0_ob_out[7], \kme_cceip0_ob_out.tdata [7]);
tran (kme_cceip0_ob_out[6], \kme_cceip0_ob_out.tdata [6]);
tran (kme_cceip0_ob_out[5], \kme_cceip0_ob_out.tdata [5]);
tran (kme_cceip0_ob_out[4], \kme_cceip0_ob_out.tdata [4]);
tran (kme_cceip0_ob_out[3], \kme_cceip0_ob_out.tdata [3]);
tran (kme_cceip0_ob_out[2], \kme_cceip0_ob_out.tdata [2]);
tran (kme_cceip0_ob_out[1], \kme_cceip0_ob_out.tdata [1]);
tran (kme_cceip0_ob_out[0], \kme_cceip0_ob_out.tdata [0]);
tran (kme_cceip0_ob_in_mod[0], \kme_cceip0_ob_in_mod.tready );
tran (kme_cceip1_ob_out[82], \kme_cceip1_ob_out.tvalid );
tran (kme_cceip1_ob_out[81], \kme_cceip1_ob_out.tlast );
tran (kme_cceip1_ob_out[80], \kme_cceip1_ob_out.tid [0]);
tran (kme_cceip1_ob_out[79], \kme_cceip1_ob_out.tstrb [7]);
tran (kme_cceip1_ob_out[78], \kme_cceip1_ob_out.tstrb [6]);
tran (kme_cceip1_ob_out[77], \kme_cceip1_ob_out.tstrb [5]);
tran (kme_cceip1_ob_out[76], \kme_cceip1_ob_out.tstrb [4]);
tran (kme_cceip1_ob_out[75], \kme_cceip1_ob_out.tstrb [3]);
tran (kme_cceip1_ob_out[74], \kme_cceip1_ob_out.tstrb [2]);
tran (kme_cceip1_ob_out[73], \kme_cceip1_ob_out.tstrb [1]);
tran (kme_cceip1_ob_out[72], \kme_cceip1_ob_out.tstrb [0]);
tran (kme_cceip1_ob_out[71], \kme_cceip1_ob_out.tuser [7]);
tran (kme_cceip1_ob_out[70], \kme_cceip1_ob_out.tuser [6]);
tran (kme_cceip1_ob_out[69], \kme_cceip1_ob_out.tuser [5]);
tran (kme_cceip1_ob_out[68], \kme_cceip1_ob_out.tuser [4]);
tran (kme_cceip1_ob_out[67], \kme_cceip1_ob_out.tuser [3]);
tran (kme_cceip1_ob_out[66], \kme_cceip1_ob_out.tuser [2]);
tran (kme_cceip1_ob_out[65], \kme_cceip1_ob_out.tuser [1]);
tran (kme_cceip1_ob_out[64], \kme_cceip1_ob_out.tuser [0]);
tran (kme_cceip1_ob_out[63], \kme_cceip1_ob_out.tdata [63]);
tran (kme_cceip1_ob_out[62], \kme_cceip1_ob_out.tdata [62]);
tran (kme_cceip1_ob_out[61], \kme_cceip1_ob_out.tdata [61]);
tran (kme_cceip1_ob_out[60], \kme_cceip1_ob_out.tdata [60]);
tran (kme_cceip1_ob_out[59], \kme_cceip1_ob_out.tdata [59]);
tran (kme_cceip1_ob_out[58], \kme_cceip1_ob_out.tdata [58]);
tran (kme_cceip1_ob_out[57], \kme_cceip1_ob_out.tdata [57]);
tran (kme_cceip1_ob_out[56], \kme_cceip1_ob_out.tdata [56]);
tran (kme_cceip1_ob_out[55], \kme_cceip1_ob_out.tdata [55]);
tran (kme_cceip1_ob_out[54], \kme_cceip1_ob_out.tdata [54]);
tran (kme_cceip1_ob_out[53], \kme_cceip1_ob_out.tdata [53]);
tran (kme_cceip1_ob_out[52], \kme_cceip1_ob_out.tdata [52]);
tran (kme_cceip1_ob_out[51], \kme_cceip1_ob_out.tdata [51]);
tran (kme_cceip1_ob_out[50], \kme_cceip1_ob_out.tdata [50]);
tran (kme_cceip1_ob_out[49], \kme_cceip1_ob_out.tdata [49]);
tran (kme_cceip1_ob_out[48], \kme_cceip1_ob_out.tdata [48]);
tran (kme_cceip1_ob_out[47], \kme_cceip1_ob_out.tdata [47]);
tran (kme_cceip1_ob_out[46], \kme_cceip1_ob_out.tdata [46]);
tran (kme_cceip1_ob_out[45], \kme_cceip1_ob_out.tdata [45]);
tran (kme_cceip1_ob_out[44], \kme_cceip1_ob_out.tdata [44]);
tran (kme_cceip1_ob_out[43], \kme_cceip1_ob_out.tdata [43]);
tran (kme_cceip1_ob_out[42], \kme_cceip1_ob_out.tdata [42]);
tran (kme_cceip1_ob_out[41], \kme_cceip1_ob_out.tdata [41]);
tran (kme_cceip1_ob_out[40], \kme_cceip1_ob_out.tdata [40]);
tran (kme_cceip1_ob_out[39], \kme_cceip1_ob_out.tdata [39]);
tran (kme_cceip1_ob_out[38], \kme_cceip1_ob_out.tdata [38]);
tran (kme_cceip1_ob_out[37], \kme_cceip1_ob_out.tdata [37]);
tran (kme_cceip1_ob_out[36], \kme_cceip1_ob_out.tdata [36]);
tran (kme_cceip1_ob_out[35], \kme_cceip1_ob_out.tdata [35]);
tran (kme_cceip1_ob_out[34], \kme_cceip1_ob_out.tdata [34]);
tran (kme_cceip1_ob_out[33], \kme_cceip1_ob_out.tdata [33]);
tran (kme_cceip1_ob_out[32], \kme_cceip1_ob_out.tdata [32]);
tran (kme_cceip1_ob_out[31], \kme_cceip1_ob_out.tdata [31]);
tran (kme_cceip1_ob_out[30], \kme_cceip1_ob_out.tdata [30]);
tran (kme_cceip1_ob_out[29], \kme_cceip1_ob_out.tdata [29]);
tran (kme_cceip1_ob_out[28], \kme_cceip1_ob_out.tdata [28]);
tran (kme_cceip1_ob_out[27], \kme_cceip1_ob_out.tdata [27]);
tran (kme_cceip1_ob_out[26], \kme_cceip1_ob_out.tdata [26]);
tran (kme_cceip1_ob_out[25], \kme_cceip1_ob_out.tdata [25]);
tran (kme_cceip1_ob_out[24], \kme_cceip1_ob_out.tdata [24]);
tran (kme_cceip1_ob_out[23], \kme_cceip1_ob_out.tdata [23]);
tran (kme_cceip1_ob_out[22], \kme_cceip1_ob_out.tdata [22]);
tran (kme_cceip1_ob_out[21], \kme_cceip1_ob_out.tdata [21]);
tran (kme_cceip1_ob_out[20], \kme_cceip1_ob_out.tdata [20]);
tran (kme_cceip1_ob_out[19], \kme_cceip1_ob_out.tdata [19]);
tran (kme_cceip1_ob_out[18], \kme_cceip1_ob_out.tdata [18]);
tran (kme_cceip1_ob_out[17], \kme_cceip1_ob_out.tdata [17]);
tran (kme_cceip1_ob_out[16], \kme_cceip1_ob_out.tdata [16]);
tran (kme_cceip1_ob_out[15], \kme_cceip1_ob_out.tdata [15]);
tran (kme_cceip1_ob_out[14], \kme_cceip1_ob_out.tdata [14]);
tran (kme_cceip1_ob_out[13], \kme_cceip1_ob_out.tdata [13]);
tran (kme_cceip1_ob_out[12], \kme_cceip1_ob_out.tdata [12]);
tran (kme_cceip1_ob_out[11], \kme_cceip1_ob_out.tdata [11]);
tran (kme_cceip1_ob_out[10], \kme_cceip1_ob_out.tdata [10]);
tran (kme_cceip1_ob_out[9], \kme_cceip1_ob_out.tdata [9]);
tran (kme_cceip1_ob_out[8], \kme_cceip1_ob_out.tdata [8]);
tran (kme_cceip1_ob_out[7], \kme_cceip1_ob_out.tdata [7]);
tran (kme_cceip1_ob_out[6], \kme_cceip1_ob_out.tdata [6]);
tran (kme_cceip1_ob_out[5], \kme_cceip1_ob_out.tdata [5]);
tran (kme_cceip1_ob_out[4], \kme_cceip1_ob_out.tdata [4]);
tran (kme_cceip1_ob_out[3], \kme_cceip1_ob_out.tdata [3]);
tran (kme_cceip1_ob_out[2], \kme_cceip1_ob_out.tdata [2]);
tran (kme_cceip1_ob_out[1], \kme_cceip1_ob_out.tdata [1]);
tran (kme_cceip1_ob_out[0], \kme_cceip1_ob_out.tdata [0]);
tran (kme_cceip1_ob_in_mod[0], \kme_cceip1_ob_in_mod.tready );
tran (kme_cceip2_ob_out[82], \kme_cceip2_ob_out.tvalid );
tran (kme_cceip2_ob_out[81], \kme_cceip2_ob_out.tlast );
tran (kme_cceip2_ob_out[80], \kme_cceip2_ob_out.tid [0]);
tran (kme_cceip2_ob_out[79], \kme_cceip2_ob_out.tstrb [7]);
tran (kme_cceip2_ob_out[78], \kme_cceip2_ob_out.tstrb [6]);
tran (kme_cceip2_ob_out[77], \kme_cceip2_ob_out.tstrb [5]);
tran (kme_cceip2_ob_out[76], \kme_cceip2_ob_out.tstrb [4]);
tran (kme_cceip2_ob_out[75], \kme_cceip2_ob_out.tstrb [3]);
tran (kme_cceip2_ob_out[74], \kme_cceip2_ob_out.tstrb [2]);
tran (kme_cceip2_ob_out[73], \kme_cceip2_ob_out.tstrb [1]);
tran (kme_cceip2_ob_out[72], \kme_cceip2_ob_out.tstrb [0]);
tran (kme_cceip2_ob_out[71], \kme_cceip2_ob_out.tuser [7]);
tran (kme_cceip2_ob_out[70], \kme_cceip2_ob_out.tuser [6]);
tran (kme_cceip2_ob_out[69], \kme_cceip2_ob_out.tuser [5]);
tran (kme_cceip2_ob_out[68], \kme_cceip2_ob_out.tuser [4]);
tran (kme_cceip2_ob_out[67], \kme_cceip2_ob_out.tuser [3]);
tran (kme_cceip2_ob_out[66], \kme_cceip2_ob_out.tuser [2]);
tran (kme_cceip2_ob_out[65], \kme_cceip2_ob_out.tuser [1]);
tran (kme_cceip2_ob_out[64], \kme_cceip2_ob_out.tuser [0]);
tran (kme_cceip2_ob_out[63], \kme_cceip2_ob_out.tdata [63]);
tran (kme_cceip2_ob_out[62], \kme_cceip2_ob_out.tdata [62]);
tran (kme_cceip2_ob_out[61], \kme_cceip2_ob_out.tdata [61]);
tran (kme_cceip2_ob_out[60], \kme_cceip2_ob_out.tdata [60]);
tran (kme_cceip2_ob_out[59], \kme_cceip2_ob_out.tdata [59]);
tran (kme_cceip2_ob_out[58], \kme_cceip2_ob_out.tdata [58]);
tran (kme_cceip2_ob_out[57], \kme_cceip2_ob_out.tdata [57]);
tran (kme_cceip2_ob_out[56], \kme_cceip2_ob_out.tdata [56]);
tran (kme_cceip2_ob_out[55], \kme_cceip2_ob_out.tdata [55]);
tran (kme_cceip2_ob_out[54], \kme_cceip2_ob_out.tdata [54]);
tran (kme_cceip2_ob_out[53], \kme_cceip2_ob_out.tdata [53]);
tran (kme_cceip2_ob_out[52], \kme_cceip2_ob_out.tdata [52]);
tran (kme_cceip2_ob_out[51], \kme_cceip2_ob_out.tdata [51]);
tran (kme_cceip2_ob_out[50], \kme_cceip2_ob_out.tdata [50]);
tran (kme_cceip2_ob_out[49], \kme_cceip2_ob_out.tdata [49]);
tran (kme_cceip2_ob_out[48], \kme_cceip2_ob_out.tdata [48]);
tran (kme_cceip2_ob_out[47], \kme_cceip2_ob_out.tdata [47]);
tran (kme_cceip2_ob_out[46], \kme_cceip2_ob_out.tdata [46]);
tran (kme_cceip2_ob_out[45], \kme_cceip2_ob_out.tdata [45]);
tran (kme_cceip2_ob_out[44], \kme_cceip2_ob_out.tdata [44]);
tran (kme_cceip2_ob_out[43], \kme_cceip2_ob_out.tdata [43]);
tran (kme_cceip2_ob_out[42], \kme_cceip2_ob_out.tdata [42]);
tran (kme_cceip2_ob_out[41], \kme_cceip2_ob_out.tdata [41]);
tran (kme_cceip2_ob_out[40], \kme_cceip2_ob_out.tdata [40]);
tran (kme_cceip2_ob_out[39], \kme_cceip2_ob_out.tdata [39]);
tran (kme_cceip2_ob_out[38], \kme_cceip2_ob_out.tdata [38]);
tran (kme_cceip2_ob_out[37], \kme_cceip2_ob_out.tdata [37]);
tran (kme_cceip2_ob_out[36], \kme_cceip2_ob_out.tdata [36]);
tran (kme_cceip2_ob_out[35], \kme_cceip2_ob_out.tdata [35]);
tran (kme_cceip2_ob_out[34], \kme_cceip2_ob_out.tdata [34]);
tran (kme_cceip2_ob_out[33], \kme_cceip2_ob_out.tdata [33]);
tran (kme_cceip2_ob_out[32], \kme_cceip2_ob_out.tdata [32]);
tran (kme_cceip2_ob_out[31], \kme_cceip2_ob_out.tdata [31]);
tran (kme_cceip2_ob_out[30], \kme_cceip2_ob_out.tdata [30]);
tran (kme_cceip2_ob_out[29], \kme_cceip2_ob_out.tdata [29]);
tran (kme_cceip2_ob_out[28], \kme_cceip2_ob_out.tdata [28]);
tran (kme_cceip2_ob_out[27], \kme_cceip2_ob_out.tdata [27]);
tran (kme_cceip2_ob_out[26], \kme_cceip2_ob_out.tdata [26]);
tran (kme_cceip2_ob_out[25], \kme_cceip2_ob_out.tdata [25]);
tran (kme_cceip2_ob_out[24], \kme_cceip2_ob_out.tdata [24]);
tran (kme_cceip2_ob_out[23], \kme_cceip2_ob_out.tdata [23]);
tran (kme_cceip2_ob_out[22], \kme_cceip2_ob_out.tdata [22]);
tran (kme_cceip2_ob_out[21], \kme_cceip2_ob_out.tdata [21]);
tran (kme_cceip2_ob_out[20], \kme_cceip2_ob_out.tdata [20]);
tran (kme_cceip2_ob_out[19], \kme_cceip2_ob_out.tdata [19]);
tran (kme_cceip2_ob_out[18], \kme_cceip2_ob_out.tdata [18]);
tran (kme_cceip2_ob_out[17], \kme_cceip2_ob_out.tdata [17]);
tran (kme_cceip2_ob_out[16], \kme_cceip2_ob_out.tdata [16]);
tran (kme_cceip2_ob_out[15], \kme_cceip2_ob_out.tdata [15]);
tran (kme_cceip2_ob_out[14], \kme_cceip2_ob_out.tdata [14]);
tran (kme_cceip2_ob_out[13], \kme_cceip2_ob_out.tdata [13]);
tran (kme_cceip2_ob_out[12], \kme_cceip2_ob_out.tdata [12]);
tran (kme_cceip2_ob_out[11], \kme_cceip2_ob_out.tdata [11]);
tran (kme_cceip2_ob_out[10], \kme_cceip2_ob_out.tdata [10]);
tran (kme_cceip2_ob_out[9], \kme_cceip2_ob_out.tdata [9]);
tran (kme_cceip2_ob_out[8], \kme_cceip2_ob_out.tdata [8]);
tran (kme_cceip2_ob_out[7], \kme_cceip2_ob_out.tdata [7]);
tran (kme_cceip2_ob_out[6], \kme_cceip2_ob_out.tdata [6]);
tran (kme_cceip2_ob_out[5], \kme_cceip2_ob_out.tdata [5]);
tran (kme_cceip2_ob_out[4], \kme_cceip2_ob_out.tdata [4]);
tran (kme_cceip2_ob_out[3], \kme_cceip2_ob_out.tdata [3]);
tran (kme_cceip2_ob_out[2], \kme_cceip2_ob_out.tdata [2]);
tran (kme_cceip2_ob_out[1], \kme_cceip2_ob_out.tdata [1]);
tran (kme_cceip2_ob_out[0], \kme_cceip2_ob_out.tdata [0]);
tran (kme_cceip2_ob_in_mod[0], \kme_cceip2_ob_in_mod.tready );
tran (kme_cceip3_ob_out[82], \kme_cceip3_ob_out.tvalid );
tran (kme_cceip3_ob_out[81], \kme_cceip3_ob_out.tlast );
tran (kme_cceip3_ob_out[80], \kme_cceip3_ob_out.tid [0]);
tran (kme_cceip3_ob_out[79], \kme_cceip3_ob_out.tstrb [7]);
tran (kme_cceip3_ob_out[78], \kme_cceip3_ob_out.tstrb [6]);
tran (kme_cceip3_ob_out[77], \kme_cceip3_ob_out.tstrb [5]);
tran (kme_cceip3_ob_out[76], \kme_cceip3_ob_out.tstrb [4]);
tran (kme_cceip3_ob_out[75], \kme_cceip3_ob_out.tstrb [3]);
tran (kme_cceip3_ob_out[74], \kme_cceip3_ob_out.tstrb [2]);
tran (kme_cceip3_ob_out[73], \kme_cceip3_ob_out.tstrb [1]);
tran (kme_cceip3_ob_out[72], \kme_cceip3_ob_out.tstrb [0]);
tran (kme_cceip3_ob_out[71], \kme_cceip3_ob_out.tuser [7]);
tran (kme_cceip3_ob_out[70], \kme_cceip3_ob_out.tuser [6]);
tran (kme_cceip3_ob_out[69], \kme_cceip3_ob_out.tuser [5]);
tran (kme_cceip3_ob_out[68], \kme_cceip3_ob_out.tuser [4]);
tran (kme_cceip3_ob_out[67], \kme_cceip3_ob_out.tuser [3]);
tran (kme_cceip3_ob_out[66], \kme_cceip3_ob_out.tuser [2]);
tran (kme_cceip3_ob_out[65], \kme_cceip3_ob_out.tuser [1]);
tran (kme_cceip3_ob_out[64], \kme_cceip3_ob_out.tuser [0]);
tran (kme_cceip3_ob_out[63], \kme_cceip3_ob_out.tdata [63]);
tran (kme_cceip3_ob_out[62], \kme_cceip3_ob_out.tdata [62]);
tran (kme_cceip3_ob_out[61], \kme_cceip3_ob_out.tdata [61]);
tran (kme_cceip3_ob_out[60], \kme_cceip3_ob_out.tdata [60]);
tran (kme_cceip3_ob_out[59], \kme_cceip3_ob_out.tdata [59]);
tran (kme_cceip3_ob_out[58], \kme_cceip3_ob_out.tdata [58]);
tran (kme_cceip3_ob_out[57], \kme_cceip3_ob_out.tdata [57]);
tran (kme_cceip3_ob_out[56], \kme_cceip3_ob_out.tdata [56]);
tran (kme_cceip3_ob_out[55], \kme_cceip3_ob_out.tdata [55]);
tran (kme_cceip3_ob_out[54], \kme_cceip3_ob_out.tdata [54]);
tran (kme_cceip3_ob_out[53], \kme_cceip3_ob_out.tdata [53]);
tran (kme_cceip3_ob_out[52], \kme_cceip3_ob_out.tdata [52]);
tran (kme_cceip3_ob_out[51], \kme_cceip3_ob_out.tdata [51]);
tran (kme_cceip3_ob_out[50], \kme_cceip3_ob_out.tdata [50]);
tran (kme_cceip3_ob_out[49], \kme_cceip3_ob_out.tdata [49]);
tran (kme_cceip3_ob_out[48], \kme_cceip3_ob_out.tdata [48]);
tran (kme_cceip3_ob_out[47], \kme_cceip3_ob_out.tdata [47]);
tran (kme_cceip3_ob_out[46], \kme_cceip3_ob_out.tdata [46]);
tran (kme_cceip3_ob_out[45], \kme_cceip3_ob_out.tdata [45]);
tran (kme_cceip3_ob_out[44], \kme_cceip3_ob_out.tdata [44]);
tran (kme_cceip3_ob_out[43], \kme_cceip3_ob_out.tdata [43]);
tran (kme_cceip3_ob_out[42], \kme_cceip3_ob_out.tdata [42]);
tran (kme_cceip3_ob_out[41], \kme_cceip3_ob_out.tdata [41]);
tran (kme_cceip3_ob_out[40], \kme_cceip3_ob_out.tdata [40]);
tran (kme_cceip3_ob_out[39], \kme_cceip3_ob_out.tdata [39]);
tran (kme_cceip3_ob_out[38], \kme_cceip3_ob_out.tdata [38]);
tran (kme_cceip3_ob_out[37], \kme_cceip3_ob_out.tdata [37]);
tran (kme_cceip3_ob_out[36], \kme_cceip3_ob_out.tdata [36]);
tran (kme_cceip3_ob_out[35], \kme_cceip3_ob_out.tdata [35]);
tran (kme_cceip3_ob_out[34], \kme_cceip3_ob_out.tdata [34]);
tran (kme_cceip3_ob_out[33], \kme_cceip3_ob_out.tdata [33]);
tran (kme_cceip3_ob_out[32], \kme_cceip3_ob_out.tdata [32]);
tran (kme_cceip3_ob_out[31], \kme_cceip3_ob_out.tdata [31]);
tran (kme_cceip3_ob_out[30], \kme_cceip3_ob_out.tdata [30]);
tran (kme_cceip3_ob_out[29], \kme_cceip3_ob_out.tdata [29]);
tran (kme_cceip3_ob_out[28], \kme_cceip3_ob_out.tdata [28]);
tran (kme_cceip3_ob_out[27], \kme_cceip3_ob_out.tdata [27]);
tran (kme_cceip3_ob_out[26], \kme_cceip3_ob_out.tdata [26]);
tran (kme_cceip3_ob_out[25], \kme_cceip3_ob_out.tdata [25]);
tran (kme_cceip3_ob_out[24], \kme_cceip3_ob_out.tdata [24]);
tran (kme_cceip3_ob_out[23], \kme_cceip3_ob_out.tdata [23]);
tran (kme_cceip3_ob_out[22], \kme_cceip3_ob_out.tdata [22]);
tran (kme_cceip3_ob_out[21], \kme_cceip3_ob_out.tdata [21]);
tran (kme_cceip3_ob_out[20], \kme_cceip3_ob_out.tdata [20]);
tran (kme_cceip3_ob_out[19], \kme_cceip3_ob_out.tdata [19]);
tran (kme_cceip3_ob_out[18], \kme_cceip3_ob_out.tdata [18]);
tran (kme_cceip3_ob_out[17], \kme_cceip3_ob_out.tdata [17]);
tran (kme_cceip3_ob_out[16], \kme_cceip3_ob_out.tdata [16]);
tran (kme_cceip3_ob_out[15], \kme_cceip3_ob_out.tdata [15]);
tran (kme_cceip3_ob_out[14], \kme_cceip3_ob_out.tdata [14]);
tran (kme_cceip3_ob_out[13], \kme_cceip3_ob_out.tdata [13]);
tran (kme_cceip3_ob_out[12], \kme_cceip3_ob_out.tdata [12]);
tran (kme_cceip3_ob_out[11], \kme_cceip3_ob_out.tdata [11]);
tran (kme_cceip3_ob_out[10], \kme_cceip3_ob_out.tdata [10]);
tran (kme_cceip3_ob_out[9], \kme_cceip3_ob_out.tdata [9]);
tran (kme_cceip3_ob_out[8], \kme_cceip3_ob_out.tdata [8]);
tran (kme_cceip3_ob_out[7], \kme_cceip3_ob_out.tdata [7]);
tran (kme_cceip3_ob_out[6], \kme_cceip3_ob_out.tdata [6]);
tran (kme_cceip3_ob_out[5], \kme_cceip3_ob_out.tdata [5]);
tran (kme_cceip3_ob_out[4], \kme_cceip3_ob_out.tdata [4]);
tran (kme_cceip3_ob_out[3], \kme_cceip3_ob_out.tdata [3]);
tran (kme_cceip3_ob_out[2], \kme_cceip3_ob_out.tdata [2]);
tran (kme_cceip3_ob_out[1], \kme_cceip3_ob_out.tdata [1]);
tran (kme_cceip3_ob_out[0], \kme_cceip3_ob_out.tdata [0]);
tran (kme_cceip3_ob_in_mod[0], \kme_cceip3_ob_in_mod.tready );
tran (kme_cddip0_ob_out[82], \kme_cddip0_ob_out.tvalid );
tran (kme_cddip0_ob_out[81], \kme_cddip0_ob_out.tlast );
tran (kme_cddip0_ob_out[80], \kme_cddip0_ob_out.tid [0]);
tran (kme_cddip0_ob_out[79], \kme_cddip0_ob_out.tstrb [7]);
tran (kme_cddip0_ob_out[78], \kme_cddip0_ob_out.tstrb [6]);
tran (kme_cddip0_ob_out[77], \kme_cddip0_ob_out.tstrb [5]);
tran (kme_cddip0_ob_out[76], \kme_cddip0_ob_out.tstrb [4]);
tran (kme_cddip0_ob_out[75], \kme_cddip0_ob_out.tstrb [3]);
tran (kme_cddip0_ob_out[74], \kme_cddip0_ob_out.tstrb [2]);
tran (kme_cddip0_ob_out[73], \kme_cddip0_ob_out.tstrb [1]);
tran (kme_cddip0_ob_out[72], \kme_cddip0_ob_out.tstrb [0]);
tran (kme_cddip0_ob_out[71], \kme_cddip0_ob_out.tuser [7]);
tran (kme_cddip0_ob_out[70], \kme_cddip0_ob_out.tuser [6]);
tran (kme_cddip0_ob_out[69], \kme_cddip0_ob_out.tuser [5]);
tran (kme_cddip0_ob_out[68], \kme_cddip0_ob_out.tuser [4]);
tran (kme_cddip0_ob_out[67], \kme_cddip0_ob_out.tuser [3]);
tran (kme_cddip0_ob_out[66], \kme_cddip0_ob_out.tuser [2]);
tran (kme_cddip0_ob_out[65], \kme_cddip0_ob_out.tuser [1]);
tran (kme_cddip0_ob_out[64], \kme_cddip0_ob_out.tuser [0]);
tran (kme_cddip0_ob_out[63], \kme_cddip0_ob_out.tdata [63]);
tran (kme_cddip0_ob_out[62], \kme_cddip0_ob_out.tdata [62]);
tran (kme_cddip0_ob_out[61], \kme_cddip0_ob_out.tdata [61]);
tran (kme_cddip0_ob_out[60], \kme_cddip0_ob_out.tdata [60]);
tran (kme_cddip0_ob_out[59], \kme_cddip0_ob_out.tdata [59]);
tran (kme_cddip0_ob_out[58], \kme_cddip0_ob_out.tdata [58]);
tran (kme_cddip0_ob_out[57], \kme_cddip0_ob_out.tdata [57]);
tran (kme_cddip0_ob_out[56], \kme_cddip0_ob_out.tdata [56]);
tran (kme_cddip0_ob_out[55], \kme_cddip0_ob_out.tdata [55]);
tran (kme_cddip0_ob_out[54], \kme_cddip0_ob_out.tdata [54]);
tran (kme_cddip0_ob_out[53], \kme_cddip0_ob_out.tdata [53]);
tran (kme_cddip0_ob_out[52], \kme_cddip0_ob_out.tdata [52]);
tran (kme_cddip0_ob_out[51], \kme_cddip0_ob_out.tdata [51]);
tran (kme_cddip0_ob_out[50], \kme_cddip0_ob_out.tdata [50]);
tran (kme_cddip0_ob_out[49], \kme_cddip0_ob_out.tdata [49]);
tran (kme_cddip0_ob_out[48], \kme_cddip0_ob_out.tdata [48]);
tran (kme_cddip0_ob_out[47], \kme_cddip0_ob_out.tdata [47]);
tran (kme_cddip0_ob_out[46], \kme_cddip0_ob_out.tdata [46]);
tran (kme_cddip0_ob_out[45], \kme_cddip0_ob_out.tdata [45]);
tran (kme_cddip0_ob_out[44], \kme_cddip0_ob_out.tdata [44]);
tran (kme_cddip0_ob_out[43], \kme_cddip0_ob_out.tdata [43]);
tran (kme_cddip0_ob_out[42], \kme_cddip0_ob_out.tdata [42]);
tran (kme_cddip0_ob_out[41], \kme_cddip0_ob_out.tdata [41]);
tran (kme_cddip0_ob_out[40], \kme_cddip0_ob_out.tdata [40]);
tran (kme_cddip0_ob_out[39], \kme_cddip0_ob_out.tdata [39]);
tran (kme_cddip0_ob_out[38], \kme_cddip0_ob_out.tdata [38]);
tran (kme_cddip0_ob_out[37], \kme_cddip0_ob_out.tdata [37]);
tran (kme_cddip0_ob_out[36], \kme_cddip0_ob_out.tdata [36]);
tran (kme_cddip0_ob_out[35], \kme_cddip0_ob_out.tdata [35]);
tran (kme_cddip0_ob_out[34], \kme_cddip0_ob_out.tdata [34]);
tran (kme_cddip0_ob_out[33], \kme_cddip0_ob_out.tdata [33]);
tran (kme_cddip0_ob_out[32], \kme_cddip0_ob_out.tdata [32]);
tran (kme_cddip0_ob_out[31], \kme_cddip0_ob_out.tdata [31]);
tran (kme_cddip0_ob_out[30], \kme_cddip0_ob_out.tdata [30]);
tran (kme_cddip0_ob_out[29], \kme_cddip0_ob_out.tdata [29]);
tran (kme_cddip0_ob_out[28], \kme_cddip0_ob_out.tdata [28]);
tran (kme_cddip0_ob_out[27], \kme_cddip0_ob_out.tdata [27]);
tran (kme_cddip0_ob_out[26], \kme_cddip0_ob_out.tdata [26]);
tran (kme_cddip0_ob_out[25], \kme_cddip0_ob_out.tdata [25]);
tran (kme_cddip0_ob_out[24], \kme_cddip0_ob_out.tdata [24]);
tran (kme_cddip0_ob_out[23], \kme_cddip0_ob_out.tdata [23]);
tran (kme_cddip0_ob_out[22], \kme_cddip0_ob_out.tdata [22]);
tran (kme_cddip0_ob_out[21], \kme_cddip0_ob_out.tdata [21]);
tran (kme_cddip0_ob_out[20], \kme_cddip0_ob_out.tdata [20]);
tran (kme_cddip0_ob_out[19], \kme_cddip0_ob_out.tdata [19]);
tran (kme_cddip0_ob_out[18], \kme_cddip0_ob_out.tdata [18]);
tran (kme_cddip0_ob_out[17], \kme_cddip0_ob_out.tdata [17]);
tran (kme_cddip0_ob_out[16], \kme_cddip0_ob_out.tdata [16]);
tran (kme_cddip0_ob_out[15], \kme_cddip0_ob_out.tdata [15]);
tran (kme_cddip0_ob_out[14], \kme_cddip0_ob_out.tdata [14]);
tran (kme_cddip0_ob_out[13], \kme_cddip0_ob_out.tdata [13]);
tran (kme_cddip0_ob_out[12], \kme_cddip0_ob_out.tdata [12]);
tran (kme_cddip0_ob_out[11], \kme_cddip0_ob_out.tdata [11]);
tran (kme_cddip0_ob_out[10], \kme_cddip0_ob_out.tdata [10]);
tran (kme_cddip0_ob_out[9], \kme_cddip0_ob_out.tdata [9]);
tran (kme_cddip0_ob_out[8], \kme_cddip0_ob_out.tdata [8]);
tran (kme_cddip0_ob_out[7], \kme_cddip0_ob_out.tdata [7]);
tran (kme_cddip0_ob_out[6], \kme_cddip0_ob_out.tdata [6]);
tran (kme_cddip0_ob_out[5], \kme_cddip0_ob_out.tdata [5]);
tran (kme_cddip0_ob_out[4], \kme_cddip0_ob_out.tdata [4]);
tran (kme_cddip0_ob_out[3], \kme_cddip0_ob_out.tdata [3]);
tran (kme_cddip0_ob_out[2], \kme_cddip0_ob_out.tdata [2]);
tran (kme_cddip0_ob_out[1], \kme_cddip0_ob_out.tdata [1]);
tran (kme_cddip0_ob_out[0], \kme_cddip0_ob_out.tdata [0]);
tran (kme_cddip0_ob_in_mod[0], \kme_cddip0_ob_in_mod.tready );
tran (kme_cddip1_ob_out[82], \kme_cddip1_ob_out.tvalid );
tran (kme_cddip1_ob_out[81], \kme_cddip1_ob_out.tlast );
tran (kme_cddip1_ob_out[80], \kme_cddip1_ob_out.tid [0]);
tran (kme_cddip1_ob_out[79], \kme_cddip1_ob_out.tstrb [7]);
tran (kme_cddip1_ob_out[78], \kme_cddip1_ob_out.tstrb [6]);
tran (kme_cddip1_ob_out[77], \kme_cddip1_ob_out.tstrb [5]);
tran (kme_cddip1_ob_out[76], \kme_cddip1_ob_out.tstrb [4]);
tran (kme_cddip1_ob_out[75], \kme_cddip1_ob_out.tstrb [3]);
tran (kme_cddip1_ob_out[74], \kme_cddip1_ob_out.tstrb [2]);
tran (kme_cddip1_ob_out[73], \kme_cddip1_ob_out.tstrb [1]);
tran (kme_cddip1_ob_out[72], \kme_cddip1_ob_out.tstrb [0]);
tran (kme_cddip1_ob_out[71], \kme_cddip1_ob_out.tuser [7]);
tran (kme_cddip1_ob_out[70], \kme_cddip1_ob_out.tuser [6]);
tran (kme_cddip1_ob_out[69], \kme_cddip1_ob_out.tuser [5]);
tran (kme_cddip1_ob_out[68], \kme_cddip1_ob_out.tuser [4]);
tran (kme_cddip1_ob_out[67], \kme_cddip1_ob_out.tuser [3]);
tran (kme_cddip1_ob_out[66], \kme_cddip1_ob_out.tuser [2]);
tran (kme_cddip1_ob_out[65], \kme_cddip1_ob_out.tuser [1]);
tran (kme_cddip1_ob_out[64], \kme_cddip1_ob_out.tuser [0]);
tran (kme_cddip1_ob_out[63], \kme_cddip1_ob_out.tdata [63]);
tran (kme_cddip1_ob_out[62], \kme_cddip1_ob_out.tdata [62]);
tran (kme_cddip1_ob_out[61], \kme_cddip1_ob_out.tdata [61]);
tran (kme_cddip1_ob_out[60], \kme_cddip1_ob_out.tdata [60]);
tran (kme_cddip1_ob_out[59], \kme_cddip1_ob_out.tdata [59]);
tran (kme_cddip1_ob_out[58], \kme_cddip1_ob_out.tdata [58]);
tran (kme_cddip1_ob_out[57], \kme_cddip1_ob_out.tdata [57]);
tran (kme_cddip1_ob_out[56], \kme_cddip1_ob_out.tdata [56]);
tran (kme_cddip1_ob_out[55], \kme_cddip1_ob_out.tdata [55]);
tran (kme_cddip1_ob_out[54], \kme_cddip1_ob_out.tdata [54]);
tran (kme_cddip1_ob_out[53], \kme_cddip1_ob_out.tdata [53]);
tran (kme_cddip1_ob_out[52], \kme_cddip1_ob_out.tdata [52]);
tran (kme_cddip1_ob_out[51], \kme_cddip1_ob_out.tdata [51]);
tran (kme_cddip1_ob_out[50], \kme_cddip1_ob_out.tdata [50]);
tran (kme_cddip1_ob_out[49], \kme_cddip1_ob_out.tdata [49]);
tran (kme_cddip1_ob_out[48], \kme_cddip1_ob_out.tdata [48]);
tran (kme_cddip1_ob_out[47], \kme_cddip1_ob_out.tdata [47]);
tran (kme_cddip1_ob_out[46], \kme_cddip1_ob_out.tdata [46]);
tran (kme_cddip1_ob_out[45], \kme_cddip1_ob_out.tdata [45]);
tran (kme_cddip1_ob_out[44], \kme_cddip1_ob_out.tdata [44]);
tran (kme_cddip1_ob_out[43], \kme_cddip1_ob_out.tdata [43]);
tran (kme_cddip1_ob_out[42], \kme_cddip1_ob_out.tdata [42]);
tran (kme_cddip1_ob_out[41], \kme_cddip1_ob_out.tdata [41]);
tran (kme_cddip1_ob_out[40], \kme_cddip1_ob_out.tdata [40]);
tran (kme_cddip1_ob_out[39], \kme_cddip1_ob_out.tdata [39]);
tran (kme_cddip1_ob_out[38], \kme_cddip1_ob_out.tdata [38]);
tran (kme_cddip1_ob_out[37], \kme_cddip1_ob_out.tdata [37]);
tran (kme_cddip1_ob_out[36], \kme_cddip1_ob_out.tdata [36]);
tran (kme_cddip1_ob_out[35], \kme_cddip1_ob_out.tdata [35]);
tran (kme_cddip1_ob_out[34], \kme_cddip1_ob_out.tdata [34]);
tran (kme_cddip1_ob_out[33], \kme_cddip1_ob_out.tdata [33]);
tran (kme_cddip1_ob_out[32], \kme_cddip1_ob_out.tdata [32]);
tran (kme_cddip1_ob_out[31], \kme_cddip1_ob_out.tdata [31]);
tran (kme_cddip1_ob_out[30], \kme_cddip1_ob_out.tdata [30]);
tran (kme_cddip1_ob_out[29], \kme_cddip1_ob_out.tdata [29]);
tran (kme_cddip1_ob_out[28], \kme_cddip1_ob_out.tdata [28]);
tran (kme_cddip1_ob_out[27], \kme_cddip1_ob_out.tdata [27]);
tran (kme_cddip1_ob_out[26], \kme_cddip1_ob_out.tdata [26]);
tran (kme_cddip1_ob_out[25], \kme_cddip1_ob_out.tdata [25]);
tran (kme_cddip1_ob_out[24], \kme_cddip1_ob_out.tdata [24]);
tran (kme_cddip1_ob_out[23], \kme_cddip1_ob_out.tdata [23]);
tran (kme_cddip1_ob_out[22], \kme_cddip1_ob_out.tdata [22]);
tran (kme_cddip1_ob_out[21], \kme_cddip1_ob_out.tdata [21]);
tran (kme_cddip1_ob_out[20], \kme_cddip1_ob_out.tdata [20]);
tran (kme_cddip1_ob_out[19], \kme_cddip1_ob_out.tdata [19]);
tran (kme_cddip1_ob_out[18], \kme_cddip1_ob_out.tdata [18]);
tran (kme_cddip1_ob_out[17], \kme_cddip1_ob_out.tdata [17]);
tran (kme_cddip1_ob_out[16], \kme_cddip1_ob_out.tdata [16]);
tran (kme_cddip1_ob_out[15], \kme_cddip1_ob_out.tdata [15]);
tran (kme_cddip1_ob_out[14], \kme_cddip1_ob_out.tdata [14]);
tran (kme_cddip1_ob_out[13], \kme_cddip1_ob_out.tdata [13]);
tran (kme_cddip1_ob_out[12], \kme_cddip1_ob_out.tdata [12]);
tran (kme_cddip1_ob_out[11], \kme_cddip1_ob_out.tdata [11]);
tran (kme_cddip1_ob_out[10], \kme_cddip1_ob_out.tdata [10]);
tran (kme_cddip1_ob_out[9], \kme_cddip1_ob_out.tdata [9]);
tran (kme_cddip1_ob_out[8], \kme_cddip1_ob_out.tdata [8]);
tran (kme_cddip1_ob_out[7], \kme_cddip1_ob_out.tdata [7]);
tran (kme_cddip1_ob_out[6], \kme_cddip1_ob_out.tdata [6]);
tran (kme_cddip1_ob_out[5], \kme_cddip1_ob_out.tdata [5]);
tran (kme_cddip1_ob_out[4], \kme_cddip1_ob_out.tdata [4]);
tran (kme_cddip1_ob_out[3], \kme_cddip1_ob_out.tdata [3]);
tran (kme_cddip1_ob_out[2], \kme_cddip1_ob_out.tdata [2]);
tran (kme_cddip1_ob_out[1], \kme_cddip1_ob_out.tdata [1]);
tran (kme_cddip1_ob_out[0], \kme_cddip1_ob_out.tdata [0]);
tran (kme_cddip1_ob_in_mod[0], \kme_cddip1_ob_in_mod.tready );
tran (kme_cddip2_ob_out[82], \kme_cddip2_ob_out.tvalid );
tran (kme_cddip2_ob_out[81], \kme_cddip2_ob_out.tlast );
tran (kme_cddip2_ob_out[80], \kme_cddip2_ob_out.tid [0]);
tran (kme_cddip2_ob_out[79], \kme_cddip2_ob_out.tstrb [7]);
tran (kme_cddip2_ob_out[78], \kme_cddip2_ob_out.tstrb [6]);
tran (kme_cddip2_ob_out[77], \kme_cddip2_ob_out.tstrb [5]);
tran (kme_cddip2_ob_out[76], \kme_cddip2_ob_out.tstrb [4]);
tran (kme_cddip2_ob_out[75], \kme_cddip2_ob_out.tstrb [3]);
tran (kme_cddip2_ob_out[74], \kme_cddip2_ob_out.tstrb [2]);
tran (kme_cddip2_ob_out[73], \kme_cddip2_ob_out.tstrb [1]);
tran (kme_cddip2_ob_out[72], \kme_cddip2_ob_out.tstrb [0]);
tran (kme_cddip2_ob_out[71], \kme_cddip2_ob_out.tuser [7]);
tran (kme_cddip2_ob_out[70], \kme_cddip2_ob_out.tuser [6]);
tran (kme_cddip2_ob_out[69], \kme_cddip2_ob_out.tuser [5]);
tran (kme_cddip2_ob_out[68], \kme_cddip2_ob_out.tuser [4]);
tran (kme_cddip2_ob_out[67], \kme_cddip2_ob_out.tuser [3]);
tran (kme_cddip2_ob_out[66], \kme_cddip2_ob_out.tuser [2]);
tran (kme_cddip2_ob_out[65], \kme_cddip2_ob_out.tuser [1]);
tran (kme_cddip2_ob_out[64], \kme_cddip2_ob_out.tuser [0]);
tran (kme_cddip2_ob_out[63], \kme_cddip2_ob_out.tdata [63]);
tran (kme_cddip2_ob_out[62], \kme_cddip2_ob_out.tdata [62]);
tran (kme_cddip2_ob_out[61], \kme_cddip2_ob_out.tdata [61]);
tran (kme_cddip2_ob_out[60], \kme_cddip2_ob_out.tdata [60]);
tran (kme_cddip2_ob_out[59], \kme_cddip2_ob_out.tdata [59]);
tran (kme_cddip2_ob_out[58], \kme_cddip2_ob_out.tdata [58]);
tran (kme_cddip2_ob_out[57], \kme_cddip2_ob_out.tdata [57]);
tran (kme_cddip2_ob_out[56], \kme_cddip2_ob_out.tdata [56]);
tran (kme_cddip2_ob_out[55], \kme_cddip2_ob_out.tdata [55]);
tran (kme_cddip2_ob_out[54], \kme_cddip2_ob_out.tdata [54]);
tran (kme_cddip2_ob_out[53], \kme_cddip2_ob_out.tdata [53]);
tran (kme_cddip2_ob_out[52], \kme_cddip2_ob_out.tdata [52]);
tran (kme_cddip2_ob_out[51], \kme_cddip2_ob_out.tdata [51]);
tran (kme_cddip2_ob_out[50], \kme_cddip2_ob_out.tdata [50]);
tran (kme_cddip2_ob_out[49], \kme_cddip2_ob_out.tdata [49]);
tran (kme_cddip2_ob_out[48], \kme_cddip2_ob_out.tdata [48]);
tran (kme_cddip2_ob_out[47], \kme_cddip2_ob_out.tdata [47]);
tran (kme_cddip2_ob_out[46], \kme_cddip2_ob_out.tdata [46]);
tran (kme_cddip2_ob_out[45], \kme_cddip2_ob_out.tdata [45]);
tran (kme_cddip2_ob_out[44], \kme_cddip2_ob_out.tdata [44]);
tran (kme_cddip2_ob_out[43], \kme_cddip2_ob_out.tdata [43]);
tran (kme_cddip2_ob_out[42], \kme_cddip2_ob_out.tdata [42]);
tran (kme_cddip2_ob_out[41], \kme_cddip2_ob_out.tdata [41]);
tran (kme_cddip2_ob_out[40], \kme_cddip2_ob_out.tdata [40]);
tran (kme_cddip2_ob_out[39], \kme_cddip2_ob_out.tdata [39]);
tran (kme_cddip2_ob_out[38], \kme_cddip2_ob_out.tdata [38]);
tran (kme_cddip2_ob_out[37], \kme_cddip2_ob_out.tdata [37]);
tran (kme_cddip2_ob_out[36], \kme_cddip2_ob_out.tdata [36]);
tran (kme_cddip2_ob_out[35], \kme_cddip2_ob_out.tdata [35]);
tran (kme_cddip2_ob_out[34], \kme_cddip2_ob_out.tdata [34]);
tran (kme_cddip2_ob_out[33], \kme_cddip2_ob_out.tdata [33]);
tran (kme_cddip2_ob_out[32], \kme_cddip2_ob_out.tdata [32]);
tran (kme_cddip2_ob_out[31], \kme_cddip2_ob_out.tdata [31]);
tran (kme_cddip2_ob_out[30], \kme_cddip2_ob_out.tdata [30]);
tran (kme_cddip2_ob_out[29], \kme_cddip2_ob_out.tdata [29]);
tran (kme_cddip2_ob_out[28], \kme_cddip2_ob_out.tdata [28]);
tran (kme_cddip2_ob_out[27], \kme_cddip2_ob_out.tdata [27]);
tran (kme_cddip2_ob_out[26], \kme_cddip2_ob_out.tdata [26]);
tran (kme_cddip2_ob_out[25], \kme_cddip2_ob_out.tdata [25]);
tran (kme_cddip2_ob_out[24], \kme_cddip2_ob_out.tdata [24]);
tran (kme_cddip2_ob_out[23], \kme_cddip2_ob_out.tdata [23]);
tran (kme_cddip2_ob_out[22], \kme_cddip2_ob_out.tdata [22]);
tran (kme_cddip2_ob_out[21], \kme_cddip2_ob_out.tdata [21]);
tran (kme_cddip2_ob_out[20], \kme_cddip2_ob_out.tdata [20]);
tran (kme_cddip2_ob_out[19], \kme_cddip2_ob_out.tdata [19]);
tran (kme_cddip2_ob_out[18], \kme_cddip2_ob_out.tdata [18]);
tran (kme_cddip2_ob_out[17], \kme_cddip2_ob_out.tdata [17]);
tran (kme_cddip2_ob_out[16], \kme_cddip2_ob_out.tdata [16]);
tran (kme_cddip2_ob_out[15], \kme_cddip2_ob_out.tdata [15]);
tran (kme_cddip2_ob_out[14], \kme_cddip2_ob_out.tdata [14]);
tran (kme_cddip2_ob_out[13], \kme_cddip2_ob_out.tdata [13]);
tran (kme_cddip2_ob_out[12], \kme_cddip2_ob_out.tdata [12]);
tran (kme_cddip2_ob_out[11], \kme_cddip2_ob_out.tdata [11]);
tran (kme_cddip2_ob_out[10], \kme_cddip2_ob_out.tdata [10]);
tran (kme_cddip2_ob_out[9], \kme_cddip2_ob_out.tdata [9]);
tran (kme_cddip2_ob_out[8], \kme_cddip2_ob_out.tdata [8]);
tran (kme_cddip2_ob_out[7], \kme_cddip2_ob_out.tdata [7]);
tran (kme_cddip2_ob_out[6], \kme_cddip2_ob_out.tdata [6]);
tran (kme_cddip2_ob_out[5], \kme_cddip2_ob_out.tdata [5]);
tran (kme_cddip2_ob_out[4], \kme_cddip2_ob_out.tdata [4]);
tran (kme_cddip2_ob_out[3], \kme_cddip2_ob_out.tdata [3]);
tran (kme_cddip2_ob_out[2], \kme_cddip2_ob_out.tdata [2]);
tran (kme_cddip2_ob_out[1], \kme_cddip2_ob_out.tdata [1]);
tran (kme_cddip2_ob_out[0], \kme_cddip2_ob_out.tdata [0]);
tran (kme_cddip2_ob_in_mod[0], \kme_cddip2_ob_in_mod.tready );
tran (kme_cddip3_ob_out[82], \kme_cddip3_ob_out.tvalid );
tran (kme_cddip3_ob_out[81], \kme_cddip3_ob_out.tlast );
tran (kme_cddip3_ob_out[80], \kme_cddip3_ob_out.tid [0]);
tran (kme_cddip3_ob_out[79], \kme_cddip3_ob_out.tstrb [7]);
tran (kme_cddip3_ob_out[78], \kme_cddip3_ob_out.tstrb [6]);
tran (kme_cddip3_ob_out[77], \kme_cddip3_ob_out.tstrb [5]);
tran (kme_cddip3_ob_out[76], \kme_cddip3_ob_out.tstrb [4]);
tran (kme_cddip3_ob_out[75], \kme_cddip3_ob_out.tstrb [3]);
tran (kme_cddip3_ob_out[74], \kme_cddip3_ob_out.tstrb [2]);
tran (kme_cddip3_ob_out[73], \kme_cddip3_ob_out.tstrb [1]);
tran (kme_cddip3_ob_out[72], \kme_cddip3_ob_out.tstrb [0]);
tran (kme_cddip3_ob_out[71], \kme_cddip3_ob_out.tuser [7]);
tran (kme_cddip3_ob_out[70], \kme_cddip3_ob_out.tuser [6]);
tran (kme_cddip3_ob_out[69], \kme_cddip3_ob_out.tuser [5]);
tran (kme_cddip3_ob_out[68], \kme_cddip3_ob_out.tuser [4]);
tran (kme_cddip3_ob_out[67], \kme_cddip3_ob_out.tuser [3]);
tran (kme_cddip3_ob_out[66], \kme_cddip3_ob_out.tuser [2]);
tran (kme_cddip3_ob_out[65], \kme_cddip3_ob_out.tuser [1]);
tran (kme_cddip3_ob_out[64], \kme_cddip3_ob_out.tuser [0]);
tran (kme_cddip3_ob_out[63], \kme_cddip3_ob_out.tdata [63]);
tran (kme_cddip3_ob_out[62], \kme_cddip3_ob_out.tdata [62]);
tran (kme_cddip3_ob_out[61], \kme_cddip3_ob_out.tdata [61]);
tran (kme_cddip3_ob_out[60], \kme_cddip3_ob_out.tdata [60]);
tran (kme_cddip3_ob_out[59], \kme_cddip3_ob_out.tdata [59]);
tran (kme_cddip3_ob_out[58], \kme_cddip3_ob_out.tdata [58]);
tran (kme_cddip3_ob_out[57], \kme_cddip3_ob_out.tdata [57]);
tran (kme_cddip3_ob_out[56], \kme_cddip3_ob_out.tdata [56]);
tran (kme_cddip3_ob_out[55], \kme_cddip3_ob_out.tdata [55]);
tran (kme_cddip3_ob_out[54], \kme_cddip3_ob_out.tdata [54]);
tran (kme_cddip3_ob_out[53], \kme_cddip3_ob_out.tdata [53]);
tran (kme_cddip3_ob_out[52], \kme_cddip3_ob_out.tdata [52]);
tran (kme_cddip3_ob_out[51], \kme_cddip3_ob_out.tdata [51]);
tran (kme_cddip3_ob_out[50], \kme_cddip3_ob_out.tdata [50]);
tran (kme_cddip3_ob_out[49], \kme_cddip3_ob_out.tdata [49]);
tran (kme_cddip3_ob_out[48], \kme_cddip3_ob_out.tdata [48]);
tran (kme_cddip3_ob_out[47], \kme_cddip3_ob_out.tdata [47]);
tran (kme_cddip3_ob_out[46], \kme_cddip3_ob_out.tdata [46]);
tran (kme_cddip3_ob_out[45], \kme_cddip3_ob_out.tdata [45]);
tran (kme_cddip3_ob_out[44], \kme_cddip3_ob_out.tdata [44]);
tran (kme_cddip3_ob_out[43], \kme_cddip3_ob_out.tdata [43]);
tran (kme_cddip3_ob_out[42], \kme_cddip3_ob_out.tdata [42]);
tran (kme_cddip3_ob_out[41], \kme_cddip3_ob_out.tdata [41]);
tran (kme_cddip3_ob_out[40], \kme_cddip3_ob_out.tdata [40]);
tran (kme_cddip3_ob_out[39], \kme_cddip3_ob_out.tdata [39]);
tran (kme_cddip3_ob_out[38], \kme_cddip3_ob_out.tdata [38]);
tran (kme_cddip3_ob_out[37], \kme_cddip3_ob_out.tdata [37]);
tran (kme_cddip3_ob_out[36], \kme_cddip3_ob_out.tdata [36]);
tran (kme_cddip3_ob_out[35], \kme_cddip3_ob_out.tdata [35]);
tran (kme_cddip3_ob_out[34], \kme_cddip3_ob_out.tdata [34]);
tran (kme_cddip3_ob_out[33], \kme_cddip3_ob_out.tdata [33]);
tran (kme_cddip3_ob_out[32], \kme_cddip3_ob_out.tdata [32]);
tran (kme_cddip3_ob_out[31], \kme_cddip3_ob_out.tdata [31]);
tran (kme_cddip3_ob_out[30], \kme_cddip3_ob_out.tdata [30]);
tran (kme_cddip3_ob_out[29], \kme_cddip3_ob_out.tdata [29]);
tran (kme_cddip3_ob_out[28], \kme_cddip3_ob_out.tdata [28]);
tran (kme_cddip3_ob_out[27], \kme_cddip3_ob_out.tdata [27]);
tran (kme_cddip3_ob_out[26], \kme_cddip3_ob_out.tdata [26]);
tran (kme_cddip3_ob_out[25], \kme_cddip3_ob_out.tdata [25]);
tran (kme_cddip3_ob_out[24], \kme_cddip3_ob_out.tdata [24]);
tran (kme_cddip3_ob_out[23], \kme_cddip3_ob_out.tdata [23]);
tran (kme_cddip3_ob_out[22], \kme_cddip3_ob_out.tdata [22]);
tran (kme_cddip3_ob_out[21], \kme_cddip3_ob_out.tdata [21]);
tran (kme_cddip3_ob_out[20], \kme_cddip3_ob_out.tdata [20]);
tran (kme_cddip3_ob_out[19], \kme_cddip3_ob_out.tdata [19]);
tran (kme_cddip3_ob_out[18], \kme_cddip3_ob_out.tdata [18]);
tran (kme_cddip3_ob_out[17], \kme_cddip3_ob_out.tdata [17]);
tran (kme_cddip3_ob_out[16], \kme_cddip3_ob_out.tdata [16]);
tran (kme_cddip3_ob_out[15], \kme_cddip3_ob_out.tdata [15]);
tran (kme_cddip3_ob_out[14], \kme_cddip3_ob_out.tdata [14]);
tran (kme_cddip3_ob_out[13], \kme_cddip3_ob_out.tdata [13]);
tran (kme_cddip3_ob_out[12], \kme_cddip3_ob_out.tdata [12]);
tran (kme_cddip3_ob_out[11], \kme_cddip3_ob_out.tdata [11]);
tran (kme_cddip3_ob_out[10], \kme_cddip3_ob_out.tdata [10]);
tran (kme_cddip3_ob_out[9], \kme_cddip3_ob_out.tdata [9]);
tran (kme_cddip3_ob_out[8], \kme_cddip3_ob_out.tdata [8]);
tran (kme_cddip3_ob_out[7], \kme_cddip3_ob_out.tdata [7]);
tran (kme_cddip3_ob_out[6], \kme_cddip3_ob_out.tdata [6]);
tran (kme_cddip3_ob_out[5], \kme_cddip3_ob_out.tdata [5]);
tran (kme_cddip3_ob_out[4], \kme_cddip3_ob_out.tdata [4]);
tran (kme_cddip3_ob_out[3], \kme_cddip3_ob_out.tdata [3]);
tran (kme_cddip3_ob_out[2], \kme_cddip3_ob_out.tdata [2]);
tran (kme_cddip3_ob_out[1], \kme_cddip3_ob_out.tdata [1]);
tran (kme_cddip3_ob_out[0], \kme_cddip3_ob_out.tdata [0]);
tran (kme_cddip3_ob_in_mod[0], \kme_cddip3_ob_in_mod.tready );
tran (kim_dout[37], \kim_dout.valid [0]);
tran (kim_dout[36], \kim_dout.label_index [2]);
tran (kim_dout[35], \kim_dout.label_index [1]);
tran (kim_dout[34], \kim_dout.label_index [0]);
tran (kim_dout[33], \kim_dout.ckv_length [1]);
tran (kim_dout[32], \kim_dout.ckv_length [0]);
tran (kim_dout[31], \kim_dout.ckv_pointer [14]);
tran (kim_dout[30], \kim_dout.ckv_pointer [13]);
tran (kim_dout[29], \kim_dout.ckv_pointer [12]);
tran (kim_dout[28], \kim_dout.ckv_pointer [11]);
tran (kim_dout[27], \kim_dout.ckv_pointer [10]);
tran (kim_dout[26], \kim_dout.ckv_pointer [9]);
tran (kim_dout[25], \kim_dout.ckv_pointer [8]);
tran (kim_dout[24], \kim_dout.ckv_pointer [7]);
tran (kim_dout[23], \kim_dout.ckv_pointer [6]);
tran (kim_dout[22], \kim_dout.ckv_pointer [5]);
tran (kim_dout[21], \kim_dout.ckv_pointer [4]);
tran (kim_dout[20], \kim_dout.ckv_pointer [3]);
tran (kim_dout[19], \kim_dout.ckv_pointer [2]);
tran (kim_dout[18], \kim_dout.ckv_pointer [1]);
tran (kim_dout[17], \kim_dout.ckv_pointer [0]);
tran (kim_dout[16], \kim_dout.pf_num [3]);
tran (kim_dout[15], \kim_dout.pf_num [2]);
tran (kim_dout[14], \kim_dout.pf_num [1]);
tran (kim_dout[13], \kim_dout.pf_num [0]);
tran (kim_dout[12], \kim_dout.vf_num [11]);
tran (kim_dout[11], \kim_dout.vf_num [10]);
tran (kim_dout[10], \kim_dout.vf_num [9]);
tran (kim_dout[9], \kim_dout.vf_num [8]);
tran (kim_dout[8], \kim_dout.vf_num [7]);
tran (kim_dout[7], \kim_dout.vf_num [6]);
tran (kim_dout[6], \kim_dout.vf_num [5]);
tran (kim_dout[5], \kim_dout.vf_num [4]);
tran (kim_dout[4], \kim_dout.vf_num [3]);
tran (kim_dout[3], \kim_dout.vf_num [2]);
tran (kim_dout[2], \kim_dout.vf_num [1]);
tran (kim_dout[1], \kim_dout.vf_num [0]);
tran (kim_dout[0], \kim_dout.vf_valid [0]);
tran (\labels[0][0] , \labels[0].delimiter[0] );
tran (\labels[0][1] , \labels[0].delimiter[1] );
tran (\labels[0][2] , \labels[0].delimiter[2] );
tran (\labels[0][3] , \labels[0].delimiter[3] );
tran (\labels[0][4] , \labels[0].delimiter[4] );
tran (\labels[0][5] , \labels[0].delimiter[5] );
tran (\labels[0][6] , \labels[0].delimiter[6] );
tran (\labels[0][7] , \labels[0].delimiter[7] );
tran (\labels[0][8] , \labels[0].delimiter_valid[0] );
tran (\labels[0][9] , \labels[0].label[0] );
tran (\labels[0][10] , \labels[0].label[1] );
tran (\labels[0][11] , \labels[0].label[2] );
tran (\labels[0][12] , \labels[0].label[3] );
tran (\labels[0][13] , \labels[0].label[4] );
tran (\labels[0][14] , \labels[0].label[5] );
tran (\labels[0][15] , \labels[0].label[6] );
tran (\labels[0][16] , \labels[0].label[7] );
tran (\labels[0][17] , \labels[0].label[8] );
tran (\labels[0][18] , \labels[0].label[9] );
tran (\labels[0][19] , \labels[0].label[10] );
tran (\labels[0][20] , \labels[0].label[11] );
tran (\labels[0][21] , \labels[0].label[12] );
tran (\labels[0][22] , \labels[0].label[13] );
tran (\labels[0][23] , \labels[0].label[14] );
tran (\labels[0][24] , \labels[0].label[15] );
tran (\labels[0][25] , \labels[0].label[16] );
tran (\labels[0][26] , \labels[0].label[17] );
tran (\labels[0][27] , \labels[0].label[18] );
tran (\labels[0][28] , \labels[0].label[19] );
tran (\labels[0][29] , \labels[0].label[20] );
tran (\labels[0][30] , \labels[0].label[21] );
tran (\labels[0][31] , \labels[0].label[22] );
tran (\labels[0][32] , \labels[0].label[23] );
tran (\labels[0][33] , \labels[0].label[24] );
tran (\labels[0][34] , \labels[0].label[25] );
tran (\labels[0][35] , \labels[0].label[26] );
tran (\labels[0][36] , \labels[0].label[27] );
tran (\labels[0][37] , \labels[0].label[28] );
tran (\labels[0][38] , \labels[0].label[29] );
tran (\labels[0][39] , \labels[0].label[30] );
tran (\labels[0][40] , \labels[0].label[31] );
tran (\labels[0][41] , \labels[0].label[32] );
tran (\labels[0][42] , \labels[0].label[33] );
tran (\labels[0][43] , \labels[0].label[34] );
tran (\labels[0][44] , \labels[0].label[35] );
tran (\labels[0][45] , \labels[0].label[36] );
tran (\labels[0][46] , \labels[0].label[37] );
tran (\labels[0][47] , \labels[0].label[38] );
tran (\labels[0][48] , \labels[0].label[39] );
tran (\labels[0][49] , \labels[0].label[40] );
tran (\labels[0][50] , \labels[0].label[41] );
tran (\labels[0][51] , \labels[0].label[42] );
tran (\labels[0][52] , \labels[0].label[43] );
tran (\labels[0][53] , \labels[0].label[44] );
tran (\labels[0][54] , \labels[0].label[45] );
tran (\labels[0][55] , \labels[0].label[46] );
tran (\labels[0][56] , \labels[0].label[47] );
tran (\labels[0][57] , \labels[0].label[48] );
tran (\labels[0][58] , \labels[0].label[49] );
tran (\labels[0][59] , \labels[0].label[50] );
tran (\labels[0][60] , \labels[0].label[51] );
tran (\labels[0][61] , \labels[0].label[52] );
tran (\labels[0][62] , \labels[0].label[53] );
tran (\labels[0][63] , \labels[0].label[54] );
tran (\labels[0][64] , \labels[0].label[55] );
tran (\labels[0][65] , \labels[0].label[56] );
tran (\labels[0][66] , \labels[0].label[57] );
tran (\labels[0][67] , \labels[0].label[58] );
tran (\labels[0][68] , \labels[0].label[59] );
tran (\labels[0][69] , \labels[0].label[60] );
tran (\labels[0][70] , \labels[0].label[61] );
tran (\labels[0][71] , \labels[0].label[62] );
tran (\labels[0][72] , \labels[0].label[63] );
tran (\labels[0][73] , \labels[0].label[64] );
tran (\labels[0][74] , \labels[0].label[65] );
tran (\labels[0][75] , \labels[0].label[66] );
tran (\labels[0][76] , \labels[0].label[67] );
tran (\labels[0][77] , \labels[0].label[68] );
tran (\labels[0][78] , \labels[0].label[69] );
tran (\labels[0][79] , \labels[0].label[70] );
tran (\labels[0][80] , \labels[0].label[71] );
tran (\labels[0][81] , \labels[0].label[72] );
tran (\labels[0][82] , \labels[0].label[73] );
tran (\labels[0][83] , \labels[0].label[74] );
tran (\labels[0][84] , \labels[0].label[75] );
tran (\labels[0][85] , \labels[0].label[76] );
tran (\labels[0][86] , \labels[0].label[77] );
tran (\labels[0][87] , \labels[0].label[78] );
tran (\labels[0][88] , \labels[0].label[79] );
tran (\labels[0][89] , \labels[0].label[80] );
tran (\labels[0][90] , \labels[0].label[81] );
tran (\labels[0][91] , \labels[0].label[82] );
tran (\labels[0][92] , \labels[0].label[83] );
tran (\labels[0][93] , \labels[0].label[84] );
tran (\labels[0][94] , \labels[0].label[85] );
tran (\labels[0][95] , \labels[0].label[86] );
tran (\labels[0][96] , \labels[0].label[87] );
tran (\labels[0][97] , \labels[0].label[88] );
tran (\labels[0][98] , \labels[0].label[89] );
tran (\labels[0][99] , \labels[0].label[90] );
tran (\labels[0][100] , \labels[0].label[91] );
tran (\labels[0][101] , \labels[0].label[92] );
tran (\labels[0][102] , \labels[0].label[93] );
tran (\labels[0][103] , \labels[0].label[94] );
tran (\labels[0][104] , \labels[0].label[95] );
tran (\labels[0][105] , \labels[0].label[96] );
tran (\labels[0][106] , \labels[0].label[97] );
tran (\labels[0][107] , \labels[0].label[98] );
tran (\labels[0][108] , \labels[0].label[99] );
tran (\labels[0][109] , \labels[0].label[100] );
tran (\labels[0][110] , \labels[0].label[101] );
tran (\labels[0][111] , \labels[0].label[102] );
tran (\labels[0][112] , \labels[0].label[103] );
tran (\labels[0][113] , \labels[0].label[104] );
tran (\labels[0][114] , \labels[0].label[105] );
tran (\labels[0][115] , \labels[0].label[106] );
tran (\labels[0][116] , \labels[0].label[107] );
tran (\labels[0][117] , \labels[0].label[108] );
tran (\labels[0][118] , \labels[0].label[109] );
tran (\labels[0][119] , \labels[0].label[110] );
tran (\labels[0][120] , \labels[0].label[111] );
tran (\labels[0][121] , \labels[0].label[112] );
tran (\labels[0][122] , \labels[0].label[113] );
tran (\labels[0][123] , \labels[0].label[114] );
tran (\labels[0][124] , \labels[0].label[115] );
tran (\labels[0][125] , \labels[0].label[116] );
tran (\labels[0][126] , \labels[0].label[117] );
tran (\labels[0][127] , \labels[0].label[118] );
tran (\labels[0][128] , \labels[0].label[119] );
tran (\labels[0][129] , \labels[0].label[120] );
tran (\labels[0][130] , \labels[0].label[121] );
tran (\labels[0][131] , \labels[0].label[122] );
tran (\labels[0][132] , \labels[0].label[123] );
tran (\labels[0][133] , \labels[0].label[124] );
tran (\labels[0][134] , \labels[0].label[125] );
tran (\labels[0][135] , \labels[0].label[126] );
tran (\labels[0][136] , \labels[0].label[127] );
tran (\labels[0][137] , \labels[0].label[128] );
tran (\labels[0][138] , \labels[0].label[129] );
tran (\labels[0][139] , \labels[0].label[130] );
tran (\labels[0][140] , \labels[0].label[131] );
tran (\labels[0][141] , \labels[0].label[132] );
tran (\labels[0][142] , \labels[0].label[133] );
tran (\labels[0][143] , \labels[0].label[134] );
tran (\labels[0][144] , \labels[0].label[135] );
tran (\labels[0][145] , \labels[0].label[136] );
tran (\labels[0][146] , \labels[0].label[137] );
tran (\labels[0][147] , \labels[0].label[138] );
tran (\labels[0][148] , \labels[0].label[139] );
tran (\labels[0][149] , \labels[0].label[140] );
tran (\labels[0][150] , \labels[0].label[141] );
tran (\labels[0][151] , \labels[0].label[142] );
tran (\labels[0][152] , \labels[0].label[143] );
tran (\labels[0][153] , \labels[0].label[144] );
tran (\labels[0][154] , \labels[0].label[145] );
tran (\labels[0][155] , \labels[0].label[146] );
tran (\labels[0][156] , \labels[0].label[147] );
tran (\labels[0][157] , \labels[0].label[148] );
tran (\labels[0][158] , \labels[0].label[149] );
tran (\labels[0][159] , \labels[0].label[150] );
tran (\labels[0][160] , \labels[0].label[151] );
tran (\labels[0][161] , \labels[0].label[152] );
tran (\labels[0][162] , \labels[0].label[153] );
tran (\labels[0][163] , \labels[0].label[154] );
tran (\labels[0][164] , \labels[0].label[155] );
tran (\labels[0][165] , \labels[0].label[156] );
tran (\labels[0][166] , \labels[0].label[157] );
tran (\labels[0][167] , \labels[0].label[158] );
tran (\labels[0][168] , \labels[0].label[159] );
tran (\labels[0][169] , \labels[0].label[160] );
tran (\labels[0][170] , \labels[0].label[161] );
tran (\labels[0][171] , \labels[0].label[162] );
tran (\labels[0][172] , \labels[0].label[163] );
tran (\labels[0][173] , \labels[0].label[164] );
tran (\labels[0][174] , \labels[0].label[165] );
tran (\labels[0][175] , \labels[0].label[166] );
tran (\labels[0][176] , \labels[0].label[167] );
tran (\labels[0][177] , \labels[0].label[168] );
tran (\labels[0][178] , \labels[0].label[169] );
tran (\labels[0][179] , \labels[0].label[170] );
tran (\labels[0][180] , \labels[0].label[171] );
tran (\labels[0][181] , \labels[0].label[172] );
tran (\labels[0][182] , \labels[0].label[173] );
tran (\labels[0][183] , \labels[0].label[174] );
tran (\labels[0][184] , \labels[0].label[175] );
tran (\labels[0][185] , \labels[0].label[176] );
tran (\labels[0][186] , \labels[0].label[177] );
tran (\labels[0][187] , \labels[0].label[178] );
tran (\labels[0][188] , \labels[0].label[179] );
tran (\labels[0][189] , \labels[0].label[180] );
tran (\labels[0][190] , \labels[0].label[181] );
tran (\labels[0][191] , \labels[0].label[182] );
tran (\labels[0][192] , \labels[0].label[183] );
tran (\labels[0][193] , \labels[0].label[184] );
tran (\labels[0][194] , \labels[0].label[185] );
tran (\labels[0][195] , \labels[0].label[186] );
tran (\labels[0][196] , \labels[0].label[187] );
tran (\labels[0][197] , \labels[0].label[188] );
tran (\labels[0][198] , \labels[0].label[189] );
tran (\labels[0][199] , \labels[0].label[190] );
tran (\labels[0][200] , \labels[0].label[191] );
tran (\labels[0][201] , \labels[0].label[192] );
tran (\labels[0][202] , \labels[0].label[193] );
tran (\labels[0][203] , \labels[0].label[194] );
tran (\labels[0][204] , \labels[0].label[195] );
tran (\labels[0][205] , \labels[0].label[196] );
tran (\labels[0][206] , \labels[0].label[197] );
tran (\labels[0][207] , \labels[0].label[198] );
tran (\labels[0][208] , \labels[0].label[199] );
tran (\labels[0][209] , \labels[0].label[200] );
tran (\labels[0][210] , \labels[0].label[201] );
tran (\labels[0][211] , \labels[0].label[202] );
tran (\labels[0][212] , \labels[0].label[203] );
tran (\labels[0][213] , \labels[0].label[204] );
tran (\labels[0][214] , \labels[0].label[205] );
tran (\labels[0][215] , \labels[0].label[206] );
tran (\labels[0][216] , \labels[0].label[207] );
tran (\labels[0][217] , \labels[0].label[208] );
tran (\labels[0][218] , \labels[0].label[209] );
tran (\labels[0][219] , \labels[0].label[210] );
tran (\labels[0][220] , \labels[0].label[211] );
tran (\labels[0][221] , \labels[0].label[212] );
tran (\labels[0][222] , \labels[0].label[213] );
tran (\labels[0][223] , \labels[0].label[214] );
tran (\labels[0][224] , \labels[0].label[215] );
tran (\labels[0][225] , \labels[0].label[216] );
tran (\labels[0][226] , \labels[0].label[217] );
tran (\labels[0][227] , \labels[0].label[218] );
tran (\labels[0][228] , \labels[0].label[219] );
tran (\labels[0][229] , \labels[0].label[220] );
tran (\labels[0][230] , \labels[0].label[221] );
tran (\labels[0][231] , \labels[0].label[222] );
tran (\labels[0][232] , \labels[0].label[223] );
tran (\labels[0][233] , \labels[0].label[224] );
tran (\labels[0][234] , \labels[0].label[225] );
tran (\labels[0][235] , \labels[0].label[226] );
tran (\labels[0][236] , \labels[0].label[227] );
tran (\labels[0][237] , \labels[0].label[228] );
tran (\labels[0][238] , \labels[0].label[229] );
tran (\labels[0][239] , \labels[0].label[230] );
tran (\labels[0][240] , \labels[0].label[231] );
tran (\labels[0][241] , \labels[0].label[232] );
tran (\labels[0][242] , \labels[0].label[233] );
tran (\labels[0][243] , \labels[0].label[234] );
tran (\labels[0][244] , \labels[0].label[235] );
tran (\labels[0][245] , \labels[0].label[236] );
tran (\labels[0][246] , \labels[0].label[237] );
tran (\labels[0][247] , \labels[0].label[238] );
tran (\labels[0][248] , \labels[0].label[239] );
tran (\labels[0][249] , \labels[0].label[240] );
tran (\labels[0][250] , \labels[0].label[241] );
tran (\labels[0][251] , \labels[0].label[242] );
tran (\labels[0][252] , \labels[0].label[243] );
tran (\labels[0][253] , \labels[0].label[244] );
tran (\labels[0][254] , \labels[0].label[245] );
tran (\labels[0][255] , \labels[0].label[246] );
tran (\labels[0][256] , \labels[0].label[247] );
tran (\labels[0][257] , \labels[0].label[248] );
tran (\labels[0][258] , \labels[0].label[249] );
tran (\labels[0][259] , \labels[0].label[250] );
tran (\labels[0][260] , \labels[0].label[251] );
tran (\labels[0][261] , \labels[0].label[252] );
tran (\labels[0][262] , \labels[0].label[253] );
tran (\labels[0][263] , \labels[0].label[254] );
tran (\labels[0][264] , \labels[0].label[255] );
tran (\labels[0][265] , \labels[0].label_size[0] );
tran (\labels[0][266] , \labels[0].label_size[1] );
tran (\labels[0][267] , \labels[0].label_size[2] );
tran (\labels[0][268] , \labels[0].label_size[3] );
tran (\labels[0][269] , \labels[0].label_size[4] );
tran (\labels[0][270] , \labels[0].label_size[5] );
tran (\labels[0][271] , \labels[0].guid_size[0] );
tran (\labels[1][0] , \labels[1].delimiter[0] );
tran (\labels[1][1] , \labels[1].delimiter[1] );
tran (\labels[1][2] , \labels[1].delimiter[2] );
tran (\labels[1][3] , \labels[1].delimiter[3] );
tran (\labels[1][4] , \labels[1].delimiter[4] );
tran (\labels[1][5] , \labels[1].delimiter[5] );
tran (\labels[1][6] , \labels[1].delimiter[6] );
tran (\labels[1][7] , \labels[1].delimiter[7] );
tran (\labels[1][8] , \labels[1].delimiter_valid[0] );
tran (\labels[1][9] , \labels[1].label[0] );
tran (\labels[1][10] , \labels[1].label[1] );
tran (\labels[1][11] , \labels[1].label[2] );
tran (\labels[1][12] , \labels[1].label[3] );
tran (\labels[1][13] , \labels[1].label[4] );
tran (\labels[1][14] , \labels[1].label[5] );
tran (\labels[1][15] , \labels[1].label[6] );
tran (\labels[1][16] , \labels[1].label[7] );
tran (\labels[1][17] , \labels[1].label[8] );
tran (\labels[1][18] , \labels[1].label[9] );
tran (\labels[1][19] , \labels[1].label[10] );
tran (\labels[1][20] , \labels[1].label[11] );
tran (\labels[1][21] , \labels[1].label[12] );
tran (\labels[1][22] , \labels[1].label[13] );
tran (\labels[1][23] , \labels[1].label[14] );
tran (\labels[1][24] , \labels[1].label[15] );
tran (\labels[1][25] , \labels[1].label[16] );
tran (\labels[1][26] , \labels[1].label[17] );
tran (\labels[1][27] , \labels[1].label[18] );
tran (\labels[1][28] , \labels[1].label[19] );
tran (\labels[1][29] , \labels[1].label[20] );
tran (\labels[1][30] , \labels[1].label[21] );
tran (\labels[1][31] , \labels[1].label[22] );
tran (\labels[1][32] , \labels[1].label[23] );
tran (\labels[1][33] , \labels[1].label[24] );
tran (\labels[1][34] , \labels[1].label[25] );
tran (\labels[1][35] , \labels[1].label[26] );
tran (\labels[1][36] , \labels[1].label[27] );
tran (\labels[1][37] , \labels[1].label[28] );
tran (\labels[1][38] , \labels[1].label[29] );
tran (\labels[1][39] , \labels[1].label[30] );
tran (\labels[1][40] , \labels[1].label[31] );
tran (\labels[1][41] , \labels[1].label[32] );
tran (\labels[1][42] , \labels[1].label[33] );
tran (\labels[1][43] , \labels[1].label[34] );
tran (\labels[1][44] , \labels[1].label[35] );
tran (\labels[1][45] , \labels[1].label[36] );
tran (\labels[1][46] , \labels[1].label[37] );
tran (\labels[1][47] , \labels[1].label[38] );
tran (\labels[1][48] , \labels[1].label[39] );
tran (\labels[1][49] , \labels[1].label[40] );
tran (\labels[1][50] , \labels[1].label[41] );
tran (\labels[1][51] , \labels[1].label[42] );
tran (\labels[1][52] , \labels[1].label[43] );
tran (\labels[1][53] , \labels[1].label[44] );
tran (\labels[1][54] , \labels[1].label[45] );
tran (\labels[1][55] , \labels[1].label[46] );
tran (\labels[1][56] , \labels[1].label[47] );
tran (\labels[1][57] , \labels[1].label[48] );
tran (\labels[1][58] , \labels[1].label[49] );
tran (\labels[1][59] , \labels[1].label[50] );
tran (\labels[1][60] , \labels[1].label[51] );
tran (\labels[1][61] , \labels[1].label[52] );
tran (\labels[1][62] , \labels[1].label[53] );
tran (\labels[1][63] , \labels[1].label[54] );
tran (\labels[1][64] , \labels[1].label[55] );
tran (\labels[1][65] , \labels[1].label[56] );
tran (\labels[1][66] , \labels[1].label[57] );
tran (\labels[1][67] , \labels[1].label[58] );
tran (\labels[1][68] , \labels[1].label[59] );
tran (\labels[1][69] , \labels[1].label[60] );
tran (\labels[1][70] , \labels[1].label[61] );
tran (\labels[1][71] , \labels[1].label[62] );
tran (\labels[1][72] , \labels[1].label[63] );
tran (\labels[1][73] , \labels[1].label[64] );
tran (\labels[1][74] , \labels[1].label[65] );
tran (\labels[1][75] , \labels[1].label[66] );
tran (\labels[1][76] , \labels[1].label[67] );
tran (\labels[1][77] , \labels[1].label[68] );
tran (\labels[1][78] , \labels[1].label[69] );
tran (\labels[1][79] , \labels[1].label[70] );
tran (\labels[1][80] , \labels[1].label[71] );
tran (\labels[1][81] , \labels[1].label[72] );
tran (\labels[1][82] , \labels[1].label[73] );
tran (\labels[1][83] , \labels[1].label[74] );
tran (\labels[1][84] , \labels[1].label[75] );
tran (\labels[1][85] , \labels[1].label[76] );
tran (\labels[1][86] , \labels[1].label[77] );
tran (\labels[1][87] , \labels[1].label[78] );
tran (\labels[1][88] , \labels[1].label[79] );
tran (\labels[1][89] , \labels[1].label[80] );
tran (\labels[1][90] , \labels[1].label[81] );
tran (\labels[1][91] , \labels[1].label[82] );
tran (\labels[1][92] , \labels[1].label[83] );
tran (\labels[1][93] , \labels[1].label[84] );
tran (\labels[1][94] , \labels[1].label[85] );
tran (\labels[1][95] , \labels[1].label[86] );
tran (\labels[1][96] , \labels[1].label[87] );
tran (\labels[1][97] , \labels[1].label[88] );
tran (\labels[1][98] , \labels[1].label[89] );
tran (\labels[1][99] , \labels[1].label[90] );
tran (\labels[1][100] , \labels[1].label[91] );
tran (\labels[1][101] , \labels[1].label[92] );
tran (\labels[1][102] , \labels[1].label[93] );
tran (\labels[1][103] , \labels[1].label[94] );
tran (\labels[1][104] , \labels[1].label[95] );
tran (\labels[1][105] , \labels[1].label[96] );
tran (\labels[1][106] , \labels[1].label[97] );
tran (\labels[1][107] , \labels[1].label[98] );
tran (\labels[1][108] , \labels[1].label[99] );
tran (\labels[1][109] , \labels[1].label[100] );
tran (\labels[1][110] , \labels[1].label[101] );
tran (\labels[1][111] , \labels[1].label[102] );
tran (\labels[1][112] , \labels[1].label[103] );
tran (\labels[1][113] , \labels[1].label[104] );
tran (\labels[1][114] , \labels[1].label[105] );
tran (\labels[1][115] , \labels[1].label[106] );
tran (\labels[1][116] , \labels[1].label[107] );
tran (\labels[1][117] , \labels[1].label[108] );
tran (\labels[1][118] , \labels[1].label[109] );
tran (\labels[1][119] , \labels[1].label[110] );
tran (\labels[1][120] , \labels[1].label[111] );
tran (\labels[1][121] , \labels[1].label[112] );
tran (\labels[1][122] , \labels[1].label[113] );
tran (\labels[1][123] , \labels[1].label[114] );
tran (\labels[1][124] , \labels[1].label[115] );
tran (\labels[1][125] , \labels[1].label[116] );
tran (\labels[1][126] , \labels[1].label[117] );
tran (\labels[1][127] , \labels[1].label[118] );
tran (\labels[1][128] , \labels[1].label[119] );
tran (\labels[1][129] , \labels[1].label[120] );
tran (\labels[1][130] , \labels[1].label[121] );
tran (\labels[1][131] , \labels[1].label[122] );
tran (\labels[1][132] , \labels[1].label[123] );
tran (\labels[1][133] , \labels[1].label[124] );
tran (\labels[1][134] , \labels[1].label[125] );
tran (\labels[1][135] , \labels[1].label[126] );
tran (\labels[1][136] , \labels[1].label[127] );
tran (\labels[1][137] , \labels[1].label[128] );
tran (\labels[1][138] , \labels[1].label[129] );
tran (\labels[1][139] , \labels[1].label[130] );
tran (\labels[1][140] , \labels[1].label[131] );
tran (\labels[1][141] , \labels[1].label[132] );
tran (\labels[1][142] , \labels[1].label[133] );
tran (\labels[1][143] , \labels[1].label[134] );
tran (\labels[1][144] , \labels[1].label[135] );
tran (\labels[1][145] , \labels[1].label[136] );
tran (\labels[1][146] , \labels[1].label[137] );
tran (\labels[1][147] , \labels[1].label[138] );
tran (\labels[1][148] , \labels[1].label[139] );
tran (\labels[1][149] , \labels[1].label[140] );
tran (\labels[1][150] , \labels[1].label[141] );
tran (\labels[1][151] , \labels[1].label[142] );
tran (\labels[1][152] , \labels[1].label[143] );
tran (\labels[1][153] , \labels[1].label[144] );
tran (\labels[1][154] , \labels[1].label[145] );
tran (\labels[1][155] , \labels[1].label[146] );
tran (\labels[1][156] , \labels[1].label[147] );
tran (\labels[1][157] , \labels[1].label[148] );
tran (\labels[1][158] , \labels[1].label[149] );
tran (\labels[1][159] , \labels[1].label[150] );
tran (\labels[1][160] , \labels[1].label[151] );
tran (\labels[1][161] , \labels[1].label[152] );
tran (\labels[1][162] , \labels[1].label[153] );
tran (\labels[1][163] , \labels[1].label[154] );
tran (\labels[1][164] , \labels[1].label[155] );
tran (\labels[1][165] , \labels[1].label[156] );
tran (\labels[1][166] , \labels[1].label[157] );
tran (\labels[1][167] , \labels[1].label[158] );
tran (\labels[1][168] , \labels[1].label[159] );
tran (\labels[1][169] , \labels[1].label[160] );
tran (\labels[1][170] , \labels[1].label[161] );
tran (\labels[1][171] , \labels[1].label[162] );
tran (\labels[1][172] , \labels[1].label[163] );
tran (\labels[1][173] , \labels[1].label[164] );
tran (\labels[1][174] , \labels[1].label[165] );
tran (\labels[1][175] , \labels[1].label[166] );
tran (\labels[1][176] , \labels[1].label[167] );
tran (\labels[1][177] , \labels[1].label[168] );
tran (\labels[1][178] , \labels[1].label[169] );
tran (\labels[1][179] , \labels[1].label[170] );
tran (\labels[1][180] , \labels[1].label[171] );
tran (\labels[1][181] , \labels[1].label[172] );
tran (\labels[1][182] , \labels[1].label[173] );
tran (\labels[1][183] , \labels[1].label[174] );
tran (\labels[1][184] , \labels[1].label[175] );
tran (\labels[1][185] , \labels[1].label[176] );
tran (\labels[1][186] , \labels[1].label[177] );
tran (\labels[1][187] , \labels[1].label[178] );
tran (\labels[1][188] , \labels[1].label[179] );
tran (\labels[1][189] , \labels[1].label[180] );
tran (\labels[1][190] , \labels[1].label[181] );
tran (\labels[1][191] , \labels[1].label[182] );
tran (\labels[1][192] , \labels[1].label[183] );
tran (\labels[1][193] , \labels[1].label[184] );
tran (\labels[1][194] , \labels[1].label[185] );
tran (\labels[1][195] , \labels[1].label[186] );
tran (\labels[1][196] , \labels[1].label[187] );
tran (\labels[1][197] , \labels[1].label[188] );
tran (\labels[1][198] , \labels[1].label[189] );
tran (\labels[1][199] , \labels[1].label[190] );
tran (\labels[1][200] , \labels[1].label[191] );
tran (\labels[1][201] , \labels[1].label[192] );
tran (\labels[1][202] , \labels[1].label[193] );
tran (\labels[1][203] , \labels[1].label[194] );
tran (\labels[1][204] , \labels[1].label[195] );
tran (\labels[1][205] , \labels[1].label[196] );
tran (\labels[1][206] , \labels[1].label[197] );
tran (\labels[1][207] , \labels[1].label[198] );
tran (\labels[1][208] , \labels[1].label[199] );
tran (\labels[1][209] , \labels[1].label[200] );
tran (\labels[1][210] , \labels[1].label[201] );
tran (\labels[1][211] , \labels[1].label[202] );
tran (\labels[1][212] , \labels[1].label[203] );
tran (\labels[1][213] , \labels[1].label[204] );
tran (\labels[1][214] , \labels[1].label[205] );
tran (\labels[1][215] , \labels[1].label[206] );
tran (\labels[1][216] , \labels[1].label[207] );
tran (\labels[1][217] , \labels[1].label[208] );
tran (\labels[1][218] , \labels[1].label[209] );
tran (\labels[1][219] , \labels[1].label[210] );
tran (\labels[1][220] , \labels[1].label[211] );
tran (\labels[1][221] , \labels[1].label[212] );
tran (\labels[1][222] , \labels[1].label[213] );
tran (\labels[1][223] , \labels[1].label[214] );
tran (\labels[1][224] , \labels[1].label[215] );
tran (\labels[1][225] , \labels[1].label[216] );
tran (\labels[1][226] , \labels[1].label[217] );
tran (\labels[1][227] , \labels[1].label[218] );
tran (\labels[1][228] , \labels[1].label[219] );
tran (\labels[1][229] , \labels[1].label[220] );
tran (\labels[1][230] , \labels[1].label[221] );
tran (\labels[1][231] , \labels[1].label[222] );
tran (\labels[1][232] , \labels[1].label[223] );
tran (\labels[1][233] , \labels[1].label[224] );
tran (\labels[1][234] , \labels[1].label[225] );
tran (\labels[1][235] , \labels[1].label[226] );
tran (\labels[1][236] , \labels[1].label[227] );
tran (\labels[1][237] , \labels[1].label[228] );
tran (\labels[1][238] , \labels[1].label[229] );
tran (\labels[1][239] , \labels[1].label[230] );
tran (\labels[1][240] , \labels[1].label[231] );
tran (\labels[1][241] , \labels[1].label[232] );
tran (\labels[1][242] , \labels[1].label[233] );
tran (\labels[1][243] , \labels[1].label[234] );
tran (\labels[1][244] , \labels[1].label[235] );
tran (\labels[1][245] , \labels[1].label[236] );
tran (\labels[1][246] , \labels[1].label[237] );
tran (\labels[1][247] , \labels[1].label[238] );
tran (\labels[1][248] , \labels[1].label[239] );
tran (\labels[1][249] , \labels[1].label[240] );
tran (\labels[1][250] , \labels[1].label[241] );
tran (\labels[1][251] , \labels[1].label[242] );
tran (\labels[1][252] , \labels[1].label[243] );
tran (\labels[1][253] , \labels[1].label[244] );
tran (\labels[1][254] , \labels[1].label[245] );
tran (\labels[1][255] , \labels[1].label[246] );
tran (\labels[1][256] , \labels[1].label[247] );
tran (\labels[1][257] , \labels[1].label[248] );
tran (\labels[1][258] , \labels[1].label[249] );
tran (\labels[1][259] , \labels[1].label[250] );
tran (\labels[1][260] , \labels[1].label[251] );
tran (\labels[1][261] , \labels[1].label[252] );
tran (\labels[1][262] , \labels[1].label[253] );
tran (\labels[1][263] , \labels[1].label[254] );
tran (\labels[1][264] , \labels[1].label[255] );
tran (\labels[1][265] , \labels[1].label_size[0] );
tran (\labels[1][266] , \labels[1].label_size[1] );
tran (\labels[1][267] , \labels[1].label_size[2] );
tran (\labels[1][268] , \labels[1].label_size[3] );
tran (\labels[1][269] , \labels[1].label_size[4] );
tran (\labels[1][270] , \labels[1].label_size[5] );
tran (\labels[1][271] , \labels[1].guid_size[0] );
tran (\labels[2][0] , \labels[2].delimiter[0] );
tran (\labels[2][1] , \labels[2].delimiter[1] );
tran (\labels[2][2] , \labels[2].delimiter[2] );
tran (\labels[2][3] , \labels[2].delimiter[3] );
tran (\labels[2][4] , \labels[2].delimiter[4] );
tran (\labels[2][5] , \labels[2].delimiter[5] );
tran (\labels[2][6] , \labels[2].delimiter[6] );
tran (\labels[2][7] , \labels[2].delimiter[7] );
tran (\labels[2][8] , \labels[2].delimiter_valid[0] );
tran (\labels[2][9] , \labels[2].label[0] );
tran (\labels[2][10] , \labels[2].label[1] );
tran (\labels[2][11] , \labels[2].label[2] );
tran (\labels[2][12] , \labels[2].label[3] );
tran (\labels[2][13] , \labels[2].label[4] );
tran (\labels[2][14] , \labels[2].label[5] );
tran (\labels[2][15] , \labels[2].label[6] );
tran (\labels[2][16] , \labels[2].label[7] );
tran (\labels[2][17] , \labels[2].label[8] );
tran (\labels[2][18] , \labels[2].label[9] );
tran (\labels[2][19] , \labels[2].label[10] );
tran (\labels[2][20] , \labels[2].label[11] );
tran (\labels[2][21] , \labels[2].label[12] );
tran (\labels[2][22] , \labels[2].label[13] );
tran (\labels[2][23] , \labels[2].label[14] );
tran (\labels[2][24] , \labels[2].label[15] );
tran (\labels[2][25] , \labels[2].label[16] );
tran (\labels[2][26] , \labels[2].label[17] );
tran (\labels[2][27] , \labels[2].label[18] );
tran (\labels[2][28] , \labels[2].label[19] );
tran (\labels[2][29] , \labels[2].label[20] );
tran (\labels[2][30] , \labels[2].label[21] );
tran (\labels[2][31] , \labels[2].label[22] );
tran (\labels[2][32] , \labels[2].label[23] );
tran (\labels[2][33] , \labels[2].label[24] );
tran (\labels[2][34] , \labels[2].label[25] );
tran (\labels[2][35] , \labels[2].label[26] );
tran (\labels[2][36] , \labels[2].label[27] );
tran (\labels[2][37] , \labels[2].label[28] );
tran (\labels[2][38] , \labels[2].label[29] );
tran (\labels[2][39] , \labels[2].label[30] );
tran (\labels[2][40] , \labels[2].label[31] );
tran (\labels[2][41] , \labels[2].label[32] );
tran (\labels[2][42] , \labels[2].label[33] );
tran (\labels[2][43] , \labels[2].label[34] );
tran (\labels[2][44] , \labels[2].label[35] );
tran (\labels[2][45] , \labels[2].label[36] );
tran (\labels[2][46] , \labels[2].label[37] );
tran (\labels[2][47] , \labels[2].label[38] );
tran (\labels[2][48] , \labels[2].label[39] );
tran (\labels[2][49] , \labels[2].label[40] );
tran (\labels[2][50] , \labels[2].label[41] );
tran (\labels[2][51] , \labels[2].label[42] );
tran (\labels[2][52] , \labels[2].label[43] );
tran (\labels[2][53] , \labels[2].label[44] );
tran (\labels[2][54] , \labels[2].label[45] );
tran (\labels[2][55] , \labels[2].label[46] );
tran (\labels[2][56] , \labels[2].label[47] );
tran (\labels[2][57] , \labels[2].label[48] );
tran (\labels[2][58] , \labels[2].label[49] );
tran (\labels[2][59] , \labels[2].label[50] );
tran (\labels[2][60] , \labels[2].label[51] );
tran (\labels[2][61] , \labels[2].label[52] );
tran (\labels[2][62] , \labels[2].label[53] );
tran (\labels[2][63] , \labels[2].label[54] );
tran (\labels[2][64] , \labels[2].label[55] );
tran (\labels[2][65] , \labels[2].label[56] );
tran (\labels[2][66] , \labels[2].label[57] );
tran (\labels[2][67] , \labels[2].label[58] );
tran (\labels[2][68] , \labels[2].label[59] );
tran (\labels[2][69] , \labels[2].label[60] );
tran (\labels[2][70] , \labels[2].label[61] );
tran (\labels[2][71] , \labels[2].label[62] );
tran (\labels[2][72] , \labels[2].label[63] );
tran (\labels[2][73] , \labels[2].label[64] );
tran (\labels[2][74] , \labels[2].label[65] );
tran (\labels[2][75] , \labels[2].label[66] );
tran (\labels[2][76] , \labels[2].label[67] );
tran (\labels[2][77] , \labels[2].label[68] );
tran (\labels[2][78] , \labels[2].label[69] );
tran (\labels[2][79] , \labels[2].label[70] );
tran (\labels[2][80] , \labels[2].label[71] );
tran (\labels[2][81] , \labels[2].label[72] );
tran (\labels[2][82] , \labels[2].label[73] );
tran (\labels[2][83] , \labels[2].label[74] );
tran (\labels[2][84] , \labels[2].label[75] );
tran (\labels[2][85] , \labels[2].label[76] );
tran (\labels[2][86] , \labels[2].label[77] );
tran (\labels[2][87] , \labels[2].label[78] );
tran (\labels[2][88] , \labels[2].label[79] );
tran (\labels[2][89] , \labels[2].label[80] );
tran (\labels[2][90] , \labels[2].label[81] );
tran (\labels[2][91] , \labels[2].label[82] );
tran (\labels[2][92] , \labels[2].label[83] );
tran (\labels[2][93] , \labels[2].label[84] );
tran (\labels[2][94] , \labels[2].label[85] );
tran (\labels[2][95] , \labels[2].label[86] );
tran (\labels[2][96] , \labels[2].label[87] );
tran (\labels[2][97] , \labels[2].label[88] );
tran (\labels[2][98] , \labels[2].label[89] );
tran (\labels[2][99] , \labels[2].label[90] );
tran (\labels[2][100] , \labels[2].label[91] );
tran (\labels[2][101] , \labels[2].label[92] );
tran (\labels[2][102] , \labels[2].label[93] );
tran (\labels[2][103] , \labels[2].label[94] );
tran (\labels[2][104] , \labels[2].label[95] );
tran (\labels[2][105] , \labels[2].label[96] );
tran (\labels[2][106] , \labels[2].label[97] );
tran (\labels[2][107] , \labels[2].label[98] );
tran (\labels[2][108] , \labels[2].label[99] );
tran (\labels[2][109] , \labels[2].label[100] );
tran (\labels[2][110] , \labels[2].label[101] );
tran (\labels[2][111] , \labels[2].label[102] );
tran (\labels[2][112] , \labels[2].label[103] );
tran (\labels[2][113] , \labels[2].label[104] );
tran (\labels[2][114] , \labels[2].label[105] );
tran (\labels[2][115] , \labels[2].label[106] );
tran (\labels[2][116] , \labels[2].label[107] );
tran (\labels[2][117] , \labels[2].label[108] );
tran (\labels[2][118] , \labels[2].label[109] );
tran (\labels[2][119] , \labels[2].label[110] );
tran (\labels[2][120] , \labels[2].label[111] );
tran (\labels[2][121] , \labels[2].label[112] );
tran (\labels[2][122] , \labels[2].label[113] );
tran (\labels[2][123] , \labels[2].label[114] );
tran (\labels[2][124] , \labels[2].label[115] );
tran (\labels[2][125] , \labels[2].label[116] );
tran (\labels[2][126] , \labels[2].label[117] );
tran (\labels[2][127] , \labels[2].label[118] );
tran (\labels[2][128] , \labels[2].label[119] );
tran (\labels[2][129] , \labels[2].label[120] );
tran (\labels[2][130] , \labels[2].label[121] );
tran (\labels[2][131] , \labels[2].label[122] );
tran (\labels[2][132] , \labels[2].label[123] );
tran (\labels[2][133] , \labels[2].label[124] );
tran (\labels[2][134] , \labels[2].label[125] );
tran (\labels[2][135] , \labels[2].label[126] );
tran (\labels[2][136] , \labels[2].label[127] );
tran (\labels[2][137] , \labels[2].label[128] );
tran (\labels[2][138] , \labels[2].label[129] );
tran (\labels[2][139] , \labels[2].label[130] );
tran (\labels[2][140] , \labels[2].label[131] );
tran (\labels[2][141] , \labels[2].label[132] );
tran (\labels[2][142] , \labels[2].label[133] );
tran (\labels[2][143] , \labels[2].label[134] );
tran (\labels[2][144] , \labels[2].label[135] );
tran (\labels[2][145] , \labels[2].label[136] );
tran (\labels[2][146] , \labels[2].label[137] );
tran (\labels[2][147] , \labels[2].label[138] );
tran (\labels[2][148] , \labels[2].label[139] );
tran (\labels[2][149] , \labels[2].label[140] );
tran (\labels[2][150] , \labels[2].label[141] );
tran (\labels[2][151] , \labels[2].label[142] );
tran (\labels[2][152] , \labels[2].label[143] );
tran (\labels[2][153] , \labels[2].label[144] );
tran (\labels[2][154] , \labels[2].label[145] );
tran (\labels[2][155] , \labels[2].label[146] );
tran (\labels[2][156] , \labels[2].label[147] );
tran (\labels[2][157] , \labels[2].label[148] );
tran (\labels[2][158] , \labels[2].label[149] );
tran (\labels[2][159] , \labels[2].label[150] );
tran (\labels[2][160] , \labels[2].label[151] );
tran (\labels[2][161] , \labels[2].label[152] );
tran (\labels[2][162] , \labels[2].label[153] );
tran (\labels[2][163] , \labels[2].label[154] );
tran (\labels[2][164] , \labels[2].label[155] );
tran (\labels[2][165] , \labels[2].label[156] );
tran (\labels[2][166] , \labels[2].label[157] );
tran (\labels[2][167] , \labels[2].label[158] );
tran (\labels[2][168] , \labels[2].label[159] );
tran (\labels[2][169] , \labels[2].label[160] );
tran (\labels[2][170] , \labels[2].label[161] );
tran (\labels[2][171] , \labels[2].label[162] );
tran (\labels[2][172] , \labels[2].label[163] );
tran (\labels[2][173] , \labels[2].label[164] );
tran (\labels[2][174] , \labels[2].label[165] );
tran (\labels[2][175] , \labels[2].label[166] );
tran (\labels[2][176] , \labels[2].label[167] );
tran (\labels[2][177] , \labels[2].label[168] );
tran (\labels[2][178] , \labels[2].label[169] );
tran (\labels[2][179] , \labels[2].label[170] );
tran (\labels[2][180] , \labels[2].label[171] );
tran (\labels[2][181] , \labels[2].label[172] );
tran (\labels[2][182] , \labels[2].label[173] );
tran (\labels[2][183] , \labels[2].label[174] );
tran (\labels[2][184] , \labels[2].label[175] );
tran (\labels[2][185] , \labels[2].label[176] );
tran (\labels[2][186] , \labels[2].label[177] );
tran (\labels[2][187] , \labels[2].label[178] );
tran (\labels[2][188] , \labels[2].label[179] );
tran (\labels[2][189] , \labels[2].label[180] );
tran (\labels[2][190] , \labels[2].label[181] );
tran (\labels[2][191] , \labels[2].label[182] );
tran (\labels[2][192] , \labels[2].label[183] );
tran (\labels[2][193] , \labels[2].label[184] );
tran (\labels[2][194] , \labels[2].label[185] );
tran (\labels[2][195] , \labels[2].label[186] );
tran (\labels[2][196] , \labels[2].label[187] );
tran (\labels[2][197] , \labels[2].label[188] );
tran (\labels[2][198] , \labels[2].label[189] );
tran (\labels[2][199] , \labels[2].label[190] );
tran (\labels[2][200] , \labels[2].label[191] );
tran (\labels[2][201] , \labels[2].label[192] );
tran (\labels[2][202] , \labels[2].label[193] );
tran (\labels[2][203] , \labels[2].label[194] );
tran (\labels[2][204] , \labels[2].label[195] );
tran (\labels[2][205] , \labels[2].label[196] );
tran (\labels[2][206] , \labels[2].label[197] );
tran (\labels[2][207] , \labels[2].label[198] );
tran (\labels[2][208] , \labels[2].label[199] );
tran (\labels[2][209] , \labels[2].label[200] );
tran (\labels[2][210] , \labels[2].label[201] );
tran (\labels[2][211] , \labels[2].label[202] );
tran (\labels[2][212] , \labels[2].label[203] );
tran (\labels[2][213] , \labels[2].label[204] );
tran (\labels[2][214] , \labels[2].label[205] );
tran (\labels[2][215] , \labels[2].label[206] );
tran (\labels[2][216] , \labels[2].label[207] );
tran (\labels[2][217] , \labels[2].label[208] );
tran (\labels[2][218] , \labels[2].label[209] );
tran (\labels[2][219] , \labels[2].label[210] );
tran (\labels[2][220] , \labels[2].label[211] );
tran (\labels[2][221] , \labels[2].label[212] );
tran (\labels[2][222] , \labels[2].label[213] );
tran (\labels[2][223] , \labels[2].label[214] );
tran (\labels[2][224] , \labels[2].label[215] );
tran (\labels[2][225] , \labels[2].label[216] );
tran (\labels[2][226] , \labels[2].label[217] );
tran (\labels[2][227] , \labels[2].label[218] );
tran (\labels[2][228] , \labels[2].label[219] );
tran (\labels[2][229] , \labels[2].label[220] );
tran (\labels[2][230] , \labels[2].label[221] );
tran (\labels[2][231] , \labels[2].label[222] );
tran (\labels[2][232] , \labels[2].label[223] );
tran (\labels[2][233] , \labels[2].label[224] );
tran (\labels[2][234] , \labels[2].label[225] );
tran (\labels[2][235] , \labels[2].label[226] );
tran (\labels[2][236] , \labels[2].label[227] );
tran (\labels[2][237] , \labels[2].label[228] );
tran (\labels[2][238] , \labels[2].label[229] );
tran (\labels[2][239] , \labels[2].label[230] );
tran (\labels[2][240] , \labels[2].label[231] );
tran (\labels[2][241] , \labels[2].label[232] );
tran (\labels[2][242] , \labels[2].label[233] );
tran (\labels[2][243] , \labels[2].label[234] );
tran (\labels[2][244] , \labels[2].label[235] );
tran (\labels[2][245] , \labels[2].label[236] );
tran (\labels[2][246] , \labels[2].label[237] );
tran (\labels[2][247] , \labels[2].label[238] );
tran (\labels[2][248] , \labels[2].label[239] );
tran (\labels[2][249] , \labels[2].label[240] );
tran (\labels[2][250] , \labels[2].label[241] );
tran (\labels[2][251] , \labels[2].label[242] );
tran (\labels[2][252] , \labels[2].label[243] );
tran (\labels[2][253] , \labels[2].label[244] );
tran (\labels[2][254] , \labels[2].label[245] );
tran (\labels[2][255] , \labels[2].label[246] );
tran (\labels[2][256] , \labels[2].label[247] );
tran (\labels[2][257] , \labels[2].label[248] );
tran (\labels[2][258] , \labels[2].label[249] );
tran (\labels[2][259] , \labels[2].label[250] );
tran (\labels[2][260] , \labels[2].label[251] );
tran (\labels[2][261] , \labels[2].label[252] );
tran (\labels[2][262] , \labels[2].label[253] );
tran (\labels[2][263] , \labels[2].label[254] );
tran (\labels[2][264] , \labels[2].label[255] );
tran (\labels[2][265] , \labels[2].label_size[0] );
tran (\labels[2][266] , \labels[2].label_size[1] );
tran (\labels[2][267] , \labels[2].label_size[2] );
tran (\labels[2][268] , \labels[2].label_size[3] );
tran (\labels[2][269] , \labels[2].label_size[4] );
tran (\labels[2][270] , \labels[2].label_size[5] );
tran (\labels[2][271] , \labels[2].guid_size[0] );
tran (\labels[3][0] , \labels[3].delimiter[0] );
tran (\labels[3][1] , \labels[3].delimiter[1] );
tran (\labels[3][2] , \labels[3].delimiter[2] );
tran (\labels[3][3] , \labels[3].delimiter[3] );
tran (\labels[3][4] , \labels[3].delimiter[4] );
tran (\labels[3][5] , \labels[3].delimiter[5] );
tran (\labels[3][6] , \labels[3].delimiter[6] );
tran (\labels[3][7] , \labels[3].delimiter[7] );
tran (\labels[3][8] , \labels[3].delimiter_valid[0] );
tran (\labels[3][9] , \labels[3].label[0] );
tran (\labels[3][10] , \labels[3].label[1] );
tran (\labels[3][11] , \labels[3].label[2] );
tran (\labels[3][12] , \labels[3].label[3] );
tran (\labels[3][13] , \labels[3].label[4] );
tran (\labels[3][14] , \labels[3].label[5] );
tran (\labels[3][15] , \labels[3].label[6] );
tran (\labels[3][16] , \labels[3].label[7] );
tran (\labels[3][17] , \labels[3].label[8] );
tran (\labels[3][18] , \labels[3].label[9] );
tran (\labels[3][19] , \labels[3].label[10] );
tran (\labels[3][20] , \labels[3].label[11] );
tran (\labels[3][21] , \labels[3].label[12] );
tran (\labels[3][22] , \labels[3].label[13] );
tran (\labels[3][23] , \labels[3].label[14] );
tran (\labels[3][24] , \labels[3].label[15] );
tran (\labels[3][25] , \labels[3].label[16] );
tran (\labels[3][26] , \labels[3].label[17] );
tran (\labels[3][27] , \labels[3].label[18] );
tran (\labels[3][28] , \labels[3].label[19] );
tran (\labels[3][29] , \labels[3].label[20] );
tran (\labels[3][30] , \labels[3].label[21] );
tran (\labels[3][31] , \labels[3].label[22] );
tran (\labels[3][32] , \labels[3].label[23] );
tran (\labels[3][33] , \labels[3].label[24] );
tran (\labels[3][34] , \labels[3].label[25] );
tran (\labels[3][35] , \labels[3].label[26] );
tran (\labels[3][36] , \labels[3].label[27] );
tran (\labels[3][37] , \labels[3].label[28] );
tran (\labels[3][38] , \labels[3].label[29] );
tran (\labels[3][39] , \labels[3].label[30] );
tran (\labels[3][40] , \labels[3].label[31] );
tran (\labels[3][41] , \labels[3].label[32] );
tran (\labels[3][42] , \labels[3].label[33] );
tran (\labels[3][43] , \labels[3].label[34] );
tran (\labels[3][44] , \labels[3].label[35] );
tran (\labels[3][45] , \labels[3].label[36] );
tran (\labels[3][46] , \labels[3].label[37] );
tran (\labels[3][47] , \labels[3].label[38] );
tran (\labels[3][48] , \labels[3].label[39] );
tran (\labels[3][49] , \labels[3].label[40] );
tran (\labels[3][50] , \labels[3].label[41] );
tran (\labels[3][51] , \labels[3].label[42] );
tran (\labels[3][52] , \labels[3].label[43] );
tran (\labels[3][53] , \labels[3].label[44] );
tran (\labels[3][54] , \labels[3].label[45] );
tran (\labels[3][55] , \labels[3].label[46] );
tran (\labels[3][56] , \labels[3].label[47] );
tran (\labels[3][57] , \labels[3].label[48] );
tran (\labels[3][58] , \labels[3].label[49] );
tran (\labels[3][59] , \labels[3].label[50] );
tran (\labels[3][60] , \labels[3].label[51] );
tran (\labels[3][61] , \labels[3].label[52] );
tran (\labels[3][62] , \labels[3].label[53] );
tran (\labels[3][63] , \labels[3].label[54] );
tran (\labels[3][64] , \labels[3].label[55] );
tran (\labels[3][65] , \labels[3].label[56] );
tran (\labels[3][66] , \labels[3].label[57] );
tran (\labels[3][67] , \labels[3].label[58] );
tran (\labels[3][68] , \labels[3].label[59] );
tran (\labels[3][69] , \labels[3].label[60] );
tran (\labels[3][70] , \labels[3].label[61] );
tran (\labels[3][71] , \labels[3].label[62] );
tran (\labels[3][72] , \labels[3].label[63] );
tran (\labels[3][73] , \labels[3].label[64] );
tran (\labels[3][74] , \labels[3].label[65] );
tran (\labels[3][75] , \labels[3].label[66] );
tran (\labels[3][76] , \labels[3].label[67] );
tran (\labels[3][77] , \labels[3].label[68] );
tran (\labels[3][78] , \labels[3].label[69] );
tran (\labels[3][79] , \labels[3].label[70] );
tran (\labels[3][80] , \labels[3].label[71] );
tran (\labels[3][81] , \labels[3].label[72] );
tran (\labels[3][82] , \labels[3].label[73] );
tran (\labels[3][83] , \labels[3].label[74] );
tran (\labels[3][84] , \labels[3].label[75] );
tran (\labels[3][85] , \labels[3].label[76] );
tran (\labels[3][86] , \labels[3].label[77] );
tran (\labels[3][87] , \labels[3].label[78] );
tran (\labels[3][88] , \labels[3].label[79] );
tran (\labels[3][89] , \labels[3].label[80] );
tran (\labels[3][90] , \labels[3].label[81] );
tran (\labels[3][91] , \labels[3].label[82] );
tran (\labels[3][92] , \labels[3].label[83] );
tran (\labels[3][93] , \labels[3].label[84] );
tran (\labels[3][94] , \labels[3].label[85] );
tran (\labels[3][95] , \labels[3].label[86] );
tran (\labels[3][96] , \labels[3].label[87] );
tran (\labels[3][97] , \labels[3].label[88] );
tran (\labels[3][98] , \labels[3].label[89] );
tran (\labels[3][99] , \labels[3].label[90] );
tran (\labels[3][100] , \labels[3].label[91] );
tran (\labels[3][101] , \labels[3].label[92] );
tran (\labels[3][102] , \labels[3].label[93] );
tran (\labels[3][103] , \labels[3].label[94] );
tran (\labels[3][104] , \labels[3].label[95] );
tran (\labels[3][105] , \labels[3].label[96] );
tran (\labels[3][106] , \labels[3].label[97] );
tran (\labels[3][107] , \labels[3].label[98] );
tran (\labels[3][108] , \labels[3].label[99] );
tran (\labels[3][109] , \labels[3].label[100] );
tran (\labels[3][110] , \labels[3].label[101] );
tran (\labels[3][111] , \labels[3].label[102] );
tran (\labels[3][112] , \labels[3].label[103] );
tran (\labels[3][113] , \labels[3].label[104] );
tran (\labels[3][114] , \labels[3].label[105] );
tran (\labels[3][115] , \labels[3].label[106] );
tran (\labels[3][116] , \labels[3].label[107] );
tran (\labels[3][117] , \labels[3].label[108] );
tran (\labels[3][118] , \labels[3].label[109] );
tran (\labels[3][119] , \labels[3].label[110] );
tran (\labels[3][120] , \labels[3].label[111] );
tran (\labels[3][121] , \labels[3].label[112] );
tran (\labels[3][122] , \labels[3].label[113] );
tran (\labels[3][123] , \labels[3].label[114] );
tran (\labels[3][124] , \labels[3].label[115] );
tran (\labels[3][125] , \labels[3].label[116] );
tran (\labels[3][126] , \labels[3].label[117] );
tran (\labels[3][127] , \labels[3].label[118] );
tran (\labels[3][128] , \labels[3].label[119] );
tran (\labels[3][129] , \labels[3].label[120] );
tran (\labels[3][130] , \labels[3].label[121] );
tran (\labels[3][131] , \labels[3].label[122] );
tran (\labels[3][132] , \labels[3].label[123] );
tran (\labels[3][133] , \labels[3].label[124] );
tran (\labels[3][134] , \labels[3].label[125] );
tran (\labels[3][135] , \labels[3].label[126] );
tran (\labels[3][136] , \labels[3].label[127] );
tran (\labels[3][137] , \labels[3].label[128] );
tran (\labels[3][138] , \labels[3].label[129] );
tran (\labels[3][139] , \labels[3].label[130] );
tran (\labels[3][140] , \labels[3].label[131] );
tran (\labels[3][141] , \labels[3].label[132] );
tran (\labels[3][142] , \labels[3].label[133] );
tran (\labels[3][143] , \labels[3].label[134] );
tran (\labels[3][144] , \labels[3].label[135] );
tran (\labels[3][145] , \labels[3].label[136] );
tran (\labels[3][146] , \labels[3].label[137] );
tran (\labels[3][147] , \labels[3].label[138] );
tran (\labels[3][148] , \labels[3].label[139] );
tran (\labels[3][149] , \labels[3].label[140] );
tran (\labels[3][150] , \labels[3].label[141] );
tran (\labels[3][151] , \labels[3].label[142] );
tran (\labels[3][152] , \labels[3].label[143] );
tran (\labels[3][153] , \labels[3].label[144] );
tran (\labels[3][154] , \labels[3].label[145] );
tran (\labels[3][155] , \labels[3].label[146] );
tran (\labels[3][156] , \labels[3].label[147] );
tran (\labels[3][157] , \labels[3].label[148] );
tran (\labels[3][158] , \labels[3].label[149] );
tran (\labels[3][159] , \labels[3].label[150] );
tran (\labels[3][160] , \labels[3].label[151] );
tran (\labels[3][161] , \labels[3].label[152] );
tran (\labels[3][162] , \labels[3].label[153] );
tran (\labels[3][163] , \labels[3].label[154] );
tran (\labels[3][164] , \labels[3].label[155] );
tran (\labels[3][165] , \labels[3].label[156] );
tran (\labels[3][166] , \labels[3].label[157] );
tran (\labels[3][167] , \labels[3].label[158] );
tran (\labels[3][168] , \labels[3].label[159] );
tran (\labels[3][169] , \labels[3].label[160] );
tran (\labels[3][170] , \labels[3].label[161] );
tran (\labels[3][171] , \labels[3].label[162] );
tran (\labels[3][172] , \labels[3].label[163] );
tran (\labels[3][173] , \labels[3].label[164] );
tran (\labels[3][174] , \labels[3].label[165] );
tran (\labels[3][175] , \labels[3].label[166] );
tran (\labels[3][176] , \labels[3].label[167] );
tran (\labels[3][177] , \labels[3].label[168] );
tran (\labels[3][178] , \labels[3].label[169] );
tran (\labels[3][179] , \labels[3].label[170] );
tran (\labels[3][180] , \labels[3].label[171] );
tran (\labels[3][181] , \labels[3].label[172] );
tran (\labels[3][182] , \labels[3].label[173] );
tran (\labels[3][183] , \labels[3].label[174] );
tran (\labels[3][184] , \labels[3].label[175] );
tran (\labels[3][185] , \labels[3].label[176] );
tran (\labels[3][186] , \labels[3].label[177] );
tran (\labels[3][187] , \labels[3].label[178] );
tran (\labels[3][188] , \labels[3].label[179] );
tran (\labels[3][189] , \labels[3].label[180] );
tran (\labels[3][190] , \labels[3].label[181] );
tran (\labels[3][191] , \labels[3].label[182] );
tran (\labels[3][192] , \labels[3].label[183] );
tran (\labels[3][193] , \labels[3].label[184] );
tran (\labels[3][194] , \labels[3].label[185] );
tran (\labels[3][195] , \labels[3].label[186] );
tran (\labels[3][196] , \labels[3].label[187] );
tran (\labels[3][197] , \labels[3].label[188] );
tran (\labels[3][198] , \labels[3].label[189] );
tran (\labels[3][199] , \labels[3].label[190] );
tran (\labels[3][200] , \labels[3].label[191] );
tran (\labels[3][201] , \labels[3].label[192] );
tran (\labels[3][202] , \labels[3].label[193] );
tran (\labels[3][203] , \labels[3].label[194] );
tran (\labels[3][204] , \labels[3].label[195] );
tran (\labels[3][205] , \labels[3].label[196] );
tran (\labels[3][206] , \labels[3].label[197] );
tran (\labels[3][207] , \labels[3].label[198] );
tran (\labels[3][208] , \labels[3].label[199] );
tran (\labels[3][209] , \labels[3].label[200] );
tran (\labels[3][210] , \labels[3].label[201] );
tran (\labels[3][211] , \labels[3].label[202] );
tran (\labels[3][212] , \labels[3].label[203] );
tran (\labels[3][213] , \labels[3].label[204] );
tran (\labels[3][214] , \labels[3].label[205] );
tran (\labels[3][215] , \labels[3].label[206] );
tran (\labels[3][216] , \labels[3].label[207] );
tran (\labels[3][217] , \labels[3].label[208] );
tran (\labels[3][218] , \labels[3].label[209] );
tran (\labels[3][219] , \labels[3].label[210] );
tran (\labels[3][220] , \labels[3].label[211] );
tran (\labels[3][221] , \labels[3].label[212] );
tran (\labels[3][222] , \labels[3].label[213] );
tran (\labels[3][223] , \labels[3].label[214] );
tran (\labels[3][224] , \labels[3].label[215] );
tran (\labels[3][225] , \labels[3].label[216] );
tran (\labels[3][226] , \labels[3].label[217] );
tran (\labels[3][227] , \labels[3].label[218] );
tran (\labels[3][228] , \labels[3].label[219] );
tran (\labels[3][229] , \labels[3].label[220] );
tran (\labels[3][230] , \labels[3].label[221] );
tran (\labels[3][231] , \labels[3].label[222] );
tran (\labels[3][232] , \labels[3].label[223] );
tran (\labels[3][233] , \labels[3].label[224] );
tran (\labels[3][234] , \labels[3].label[225] );
tran (\labels[3][235] , \labels[3].label[226] );
tran (\labels[3][236] , \labels[3].label[227] );
tran (\labels[3][237] , \labels[3].label[228] );
tran (\labels[3][238] , \labels[3].label[229] );
tran (\labels[3][239] , \labels[3].label[230] );
tran (\labels[3][240] , \labels[3].label[231] );
tran (\labels[3][241] , \labels[3].label[232] );
tran (\labels[3][242] , \labels[3].label[233] );
tran (\labels[3][243] , \labels[3].label[234] );
tran (\labels[3][244] , \labels[3].label[235] );
tran (\labels[3][245] , \labels[3].label[236] );
tran (\labels[3][246] , \labels[3].label[237] );
tran (\labels[3][247] , \labels[3].label[238] );
tran (\labels[3][248] , \labels[3].label[239] );
tran (\labels[3][249] , \labels[3].label[240] );
tran (\labels[3][250] , \labels[3].label[241] );
tran (\labels[3][251] , \labels[3].label[242] );
tran (\labels[3][252] , \labels[3].label[243] );
tran (\labels[3][253] , \labels[3].label[244] );
tran (\labels[3][254] , \labels[3].label[245] );
tran (\labels[3][255] , \labels[3].label[246] );
tran (\labels[3][256] , \labels[3].label[247] );
tran (\labels[3][257] , \labels[3].label[248] );
tran (\labels[3][258] , \labels[3].label[249] );
tran (\labels[3][259] , \labels[3].label[250] );
tran (\labels[3][260] , \labels[3].label[251] );
tran (\labels[3][261] , \labels[3].label[252] );
tran (\labels[3][262] , \labels[3].label[253] );
tran (\labels[3][263] , \labels[3].label[254] );
tran (\labels[3][264] , \labels[3].label[255] );
tran (\labels[3][265] , \labels[3].label_size[0] );
tran (\labels[3][266] , \labels[3].label_size[1] );
tran (\labels[3][267] , \labels[3].label_size[2] );
tran (\labels[3][268] , \labels[3].label_size[3] );
tran (\labels[3][269] , \labels[3].label_size[4] );
tran (\labels[3][270] , \labels[3].label_size[5] );
tran (\labels[3][271] , \labels[3].guid_size[0] );
tran (\labels[4][0] , \labels[4].delimiter[0] );
tran (\labels[4][1] , \labels[4].delimiter[1] );
tran (\labels[4][2] , \labels[4].delimiter[2] );
tran (\labels[4][3] , \labels[4].delimiter[3] );
tran (\labels[4][4] , \labels[4].delimiter[4] );
tran (\labels[4][5] , \labels[4].delimiter[5] );
tran (\labels[4][6] , \labels[4].delimiter[6] );
tran (\labels[4][7] , \labels[4].delimiter[7] );
tran (\labels[4][8] , \labels[4].delimiter_valid[0] );
tran (\labels[4][9] , \labels[4].label[0] );
tran (\labels[4][10] , \labels[4].label[1] );
tran (\labels[4][11] , \labels[4].label[2] );
tran (\labels[4][12] , \labels[4].label[3] );
tran (\labels[4][13] , \labels[4].label[4] );
tran (\labels[4][14] , \labels[4].label[5] );
tran (\labels[4][15] , \labels[4].label[6] );
tran (\labels[4][16] , \labels[4].label[7] );
tran (\labels[4][17] , \labels[4].label[8] );
tran (\labels[4][18] , \labels[4].label[9] );
tran (\labels[4][19] , \labels[4].label[10] );
tran (\labels[4][20] , \labels[4].label[11] );
tran (\labels[4][21] , \labels[4].label[12] );
tran (\labels[4][22] , \labels[4].label[13] );
tran (\labels[4][23] , \labels[4].label[14] );
tran (\labels[4][24] , \labels[4].label[15] );
tran (\labels[4][25] , \labels[4].label[16] );
tran (\labels[4][26] , \labels[4].label[17] );
tran (\labels[4][27] , \labels[4].label[18] );
tran (\labels[4][28] , \labels[4].label[19] );
tran (\labels[4][29] , \labels[4].label[20] );
tran (\labels[4][30] , \labels[4].label[21] );
tran (\labels[4][31] , \labels[4].label[22] );
tran (\labels[4][32] , \labels[4].label[23] );
tran (\labels[4][33] , \labels[4].label[24] );
tran (\labels[4][34] , \labels[4].label[25] );
tran (\labels[4][35] , \labels[4].label[26] );
tran (\labels[4][36] , \labels[4].label[27] );
tran (\labels[4][37] , \labels[4].label[28] );
tran (\labels[4][38] , \labels[4].label[29] );
tran (\labels[4][39] , \labels[4].label[30] );
tran (\labels[4][40] , \labels[4].label[31] );
tran (\labels[4][41] , \labels[4].label[32] );
tran (\labels[4][42] , \labels[4].label[33] );
tran (\labels[4][43] , \labels[4].label[34] );
tran (\labels[4][44] , \labels[4].label[35] );
tran (\labels[4][45] , \labels[4].label[36] );
tran (\labels[4][46] , \labels[4].label[37] );
tran (\labels[4][47] , \labels[4].label[38] );
tran (\labels[4][48] , \labels[4].label[39] );
tran (\labels[4][49] , \labels[4].label[40] );
tran (\labels[4][50] , \labels[4].label[41] );
tran (\labels[4][51] , \labels[4].label[42] );
tran (\labels[4][52] , \labels[4].label[43] );
tran (\labels[4][53] , \labels[4].label[44] );
tran (\labels[4][54] , \labels[4].label[45] );
tran (\labels[4][55] , \labels[4].label[46] );
tran (\labels[4][56] , \labels[4].label[47] );
tran (\labels[4][57] , \labels[4].label[48] );
tran (\labels[4][58] , \labels[4].label[49] );
tran (\labels[4][59] , \labels[4].label[50] );
tran (\labels[4][60] , \labels[4].label[51] );
tran (\labels[4][61] , \labels[4].label[52] );
tran (\labels[4][62] , \labels[4].label[53] );
tran (\labels[4][63] , \labels[4].label[54] );
tran (\labels[4][64] , \labels[4].label[55] );
tran (\labels[4][65] , \labels[4].label[56] );
tran (\labels[4][66] , \labels[4].label[57] );
tran (\labels[4][67] , \labels[4].label[58] );
tran (\labels[4][68] , \labels[4].label[59] );
tran (\labels[4][69] , \labels[4].label[60] );
tran (\labels[4][70] , \labels[4].label[61] );
tran (\labels[4][71] , \labels[4].label[62] );
tran (\labels[4][72] , \labels[4].label[63] );
tran (\labels[4][73] , \labels[4].label[64] );
tran (\labels[4][74] , \labels[4].label[65] );
tran (\labels[4][75] , \labels[4].label[66] );
tran (\labels[4][76] , \labels[4].label[67] );
tran (\labels[4][77] , \labels[4].label[68] );
tran (\labels[4][78] , \labels[4].label[69] );
tran (\labels[4][79] , \labels[4].label[70] );
tran (\labels[4][80] , \labels[4].label[71] );
tran (\labels[4][81] , \labels[4].label[72] );
tran (\labels[4][82] , \labels[4].label[73] );
tran (\labels[4][83] , \labels[4].label[74] );
tran (\labels[4][84] , \labels[4].label[75] );
tran (\labels[4][85] , \labels[4].label[76] );
tran (\labels[4][86] , \labels[4].label[77] );
tran (\labels[4][87] , \labels[4].label[78] );
tran (\labels[4][88] , \labels[4].label[79] );
tran (\labels[4][89] , \labels[4].label[80] );
tran (\labels[4][90] , \labels[4].label[81] );
tran (\labels[4][91] , \labels[4].label[82] );
tran (\labels[4][92] , \labels[4].label[83] );
tran (\labels[4][93] , \labels[4].label[84] );
tran (\labels[4][94] , \labels[4].label[85] );
tran (\labels[4][95] , \labels[4].label[86] );
tran (\labels[4][96] , \labels[4].label[87] );
tran (\labels[4][97] , \labels[4].label[88] );
tran (\labels[4][98] , \labels[4].label[89] );
tran (\labels[4][99] , \labels[4].label[90] );
tran (\labels[4][100] , \labels[4].label[91] );
tran (\labels[4][101] , \labels[4].label[92] );
tran (\labels[4][102] , \labels[4].label[93] );
tran (\labels[4][103] , \labels[4].label[94] );
tran (\labels[4][104] , \labels[4].label[95] );
tran (\labels[4][105] , \labels[4].label[96] );
tran (\labels[4][106] , \labels[4].label[97] );
tran (\labels[4][107] , \labels[4].label[98] );
tran (\labels[4][108] , \labels[4].label[99] );
tran (\labels[4][109] , \labels[4].label[100] );
tran (\labels[4][110] , \labels[4].label[101] );
tran (\labels[4][111] , \labels[4].label[102] );
tran (\labels[4][112] , \labels[4].label[103] );
tran (\labels[4][113] , \labels[4].label[104] );
tran (\labels[4][114] , \labels[4].label[105] );
tran (\labels[4][115] , \labels[4].label[106] );
tran (\labels[4][116] , \labels[4].label[107] );
tran (\labels[4][117] , \labels[4].label[108] );
tran (\labels[4][118] , \labels[4].label[109] );
tran (\labels[4][119] , \labels[4].label[110] );
tran (\labels[4][120] , \labels[4].label[111] );
tran (\labels[4][121] , \labels[4].label[112] );
tran (\labels[4][122] , \labels[4].label[113] );
tran (\labels[4][123] , \labels[4].label[114] );
tran (\labels[4][124] , \labels[4].label[115] );
tran (\labels[4][125] , \labels[4].label[116] );
tran (\labels[4][126] , \labels[4].label[117] );
tran (\labels[4][127] , \labels[4].label[118] );
tran (\labels[4][128] , \labels[4].label[119] );
tran (\labels[4][129] , \labels[4].label[120] );
tran (\labels[4][130] , \labels[4].label[121] );
tran (\labels[4][131] , \labels[4].label[122] );
tran (\labels[4][132] , \labels[4].label[123] );
tran (\labels[4][133] , \labels[4].label[124] );
tran (\labels[4][134] , \labels[4].label[125] );
tran (\labels[4][135] , \labels[4].label[126] );
tran (\labels[4][136] , \labels[4].label[127] );
tran (\labels[4][137] , \labels[4].label[128] );
tran (\labels[4][138] , \labels[4].label[129] );
tran (\labels[4][139] , \labels[4].label[130] );
tran (\labels[4][140] , \labels[4].label[131] );
tran (\labels[4][141] , \labels[4].label[132] );
tran (\labels[4][142] , \labels[4].label[133] );
tran (\labels[4][143] , \labels[4].label[134] );
tran (\labels[4][144] , \labels[4].label[135] );
tran (\labels[4][145] , \labels[4].label[136] );
tran (\labels[4][146] , \labels[4].label[137] );
tran (\labels[4][147] , \labels[4].label[138] );
tran (\labels[4][148] , \labels[4].label[139] );
tran (\labels[4][149] , \labels[4].label[140] );
tran (\labels[4][150] , \labels[4].label[141] );
tran (\labels[4][151] , \labels[4].label[142] );
tran (\labels[4][152] , \labels[4].label[143] );
tran (\labels[4][153] , \labels[4].label[144] );
tran (\labels[4][154] , \labels[4].label[145] );
tran (\labels[4][155] , \labels[4].label[146] );
tran (\labels[4][156] , \labels[4].label[147] );
tran (\labels[4][157] , \labels[4].label[148] );
tran (\labels[4][158] , \labels[4].label[149] );
tran (\labels[4][159] , \labels[4].label[150] );
tran (\labels[4][160] , \labels[4].label[151] );
tran (\labels[4][161] , \labels[4].label[152] );
tran (\labels[4][162] , \labels[4].label[153] );
tran (\labels[4][163] , \labels[4].label[154] );
tran (\labels[4][164] , \labels[4].label[155] );
tran (\labels[4][165] , \labels[4].label[156] );
tran (\labels[4][166] , \labels[4].label[157] );
tran (\labels[4][167] , \labels[4].label[158] );
tran (\labels[4][168] , \labels[4].label[159] );
tran (\labels[4][169] , \labels[4].label[160] );
tran (\labels[4][170] , \labels[4].label[161] );
tran (\labels[4][171] , \labels[4].label[162] );
tran (\labels[4][172] , \labels[4].label[163] );
tran (\labels[4][173] , \labels[4].label[164] );
tran (\labels[4][174] , \labels[4].label[165] );
tran (\labels[4][175] , \labels[4].label[166] );
tran (\labels[4][176] , \labels[4].label[167] );
tran (\labels[4][177] , \labels[4].label[168] );
tran (\labels[4][178] , \labels[4].label[169] );
tran (\labels[4][179] , \labels[4].label[170] );
tran (\labels[4][180] , \labels[4].label[171] );
tran (\labels[4][181] , \labels[4].label[172] );
tran (\labels[4][182] , \labels[4].label[173] );
tran (\labels[4][183] , \labels[4].label[174] );
tran (\labels[4][184] , \labels[4].label[175] );
tran (\labels[4][185] , \labels[4].label[176] );
tran (\labels[4][186] , \labels[4].label[177] );
tran (\labels[4][187] , \labels[4].label[178] );
tran (\labels[4][188] , \labels[4].label[179] );
tran (\labels[4][189] , \labels[4].label[180] );
tran (\labels[4][190] , \labels[4].label[181] );
tran (\labels[4][191] , \labels[4].label[182] );
tran (\labels[4][192] , \labels[4].label[183] );
tran (\labels[4][193] , \labels[4].label[184] );
tran (\labels[4][194] , \labels[4].label[185] );
tran (\labels[4][195] , \labels[4].label[186] );
tran (\labels[4][196] , \labels[4].label[187] );
tran (\labels[4][197] , \labels[4].label[188] );
tran (\labels[4][198] , \labels[4].label[189] );
tran (\labels[4][199] , \labels[4].label[190] );
tran (\labels[4][200] , \labels[4].label[191] );
tran (\labels[4][201] , \labels[4].label[192] );
tran (\labels[4][202] , \labels[4].label[193] );
tran (\labels[4][203] , \labels[4].label[194] );
tran (\labels[4][204] , \labels[4].label[195] );
tran (\labels[4][205] , \labels[4].label[196] );
tran (\labels[4][206] , \labels[4].label[197] );
tran (\labels[4][207] , \labels[4].label[198] );
tran (\labels[4][208] , \labels[4].label[199] );
tran (\labels[4][209] , \labels[4].label[200] );
tran (\labels[4][210] , \labels[4].label[201] );
tran (\labels[4][211] , \labels[4].label[202] );
tran (\labels[4][212] , \labels[4].label[203] );
tran (\labels[4][213] , \labels[4].label[204] );
tran (\labels[4][214] , \labels[4].label[205] );
tran (\labels[4][215] , \labels[4].label[206] );
tran (\labels[4][216] , \labels[4].label[207] );
tran (\labels[4][217] , \labels[4].label[208] );
tran (\labels[4][218] , \labels[4].label[209] );
tran (\labels[4][219] , \labels[4].label[210] );
tran (\labels[4][220] , \labels[4].label[211] );
tran (\labels[4][221] , \labels[4].label[212] );
tran (\labels[4][222] , \labels[4].label[213] );
tran (\labels[4][223] , \labels[4].label[214] );
tran (\labels[4][224] , \labels[4].label[215] );
tran (\labels[4][225] , \labels[4].label[216] );
tran (\labels[4][226] , \labels[4].label[217] );
tran (\labels[4][227] , \labels[4].label[218] );
tran (\labels[4][228] , \labels[4].label[219] );
tran (\labels[4][229] , \labels[4].label[220] );
tran (\labels[4][230] , \labels[4].label[221] );
tran (\labels[4][231] , \labels[4].label[222] );
tran (\labels[4][232] , \labels[4].label[223] );
tran (\labels[4][233] , \labels[4].label[224] );
tran (\labels[4][234] , \labels[4].label[225] );
tran (\labels[4][235] , \labels[4].label[226] );
tran (\labels[4][236] , \labels[4].label[227] );
tran (\labels[4][237] , \labels[4].label[228] );
tran (\labels[4][238] , \labels[4].label[229] );
tran (\labels[4][239] , \labels[4].label[230] );
tran (\labels[4][240] , \labels[4].label[231] );
tran (\labels[4][241] , \labels[4].label[232] );
tran (\labels[4][242] , \labels[4].label[233] );
tran (\labels[4][243] , \labels[4].label[234] );
tran (\labels[4][244] , \labels[4].label[235] );
tran (\labels[4][245] , \labels[4].label[236] );
tran (\labels[4][246] , \labels[4].label[237] );
tran (\labels[4][247] , \labels[4].label[238] );
tran (\labels[4][248] , \labels[4].label[239] );
tran (\labels[4][249] , \labels[4].label[240] );
tran (\labels[4][250] , \labels[4].label[241] );
tran (\labels[4][251] , \labels[4].label[242] );
tran (\labels[4][252] , \labels[4].label[243] );
tran (\labels[4][253] , \labels[4].label[244] );
tran (\labels[4][254] , \labels[4].label[245] );
tran (\labels[4][255] , \labels[4].label[246] );
tran (\labels[4][256] , \labels[4].label[247] );
tran (\labels[4][257] , \labels[4].label[248] );
tran (\labels[4][258] , \labels[4].label[249] );
tran (\labels[4][259] , \labels[4].label[250] );
tran (\labels[4][260] , \labels[4].label[251] );
tran (\labels[4][261] , \labels[4].label[252] );
tran (\labels[4][262] , \labels[4].label[253] );
tran (\labels[4][263] , \labels[4].label[254] );
tran (\labels[4][264] , \labels[4].label[255] );
tran (\labels[4][265] , \labels[4].label_size[0] );
tran (\labels[4][266] , \labels[4].label_size[1] );
tran (\labels[4][267] , \labels[4].label_size[2] );
tran (\labels[4][268] , \labels[4].label_size[3] );
tran (\labels[4][269] , \labels[4].label_size[4] );
tran (\labels[4][270] , \labels[4].label_size[5] );
tran (\labels[4][271] , \labels[4].guid_size[0] );
tran (\labels[5][0] , \labels[5].delimiter[0] );
tran (\labels[5][1] , \labels[5].delimiter[1] );
tran (\labels[5][2] , \labels[5].delimiter[2] );
tran (\labels[5][3] , \labels[5].delimiter[3] );
tran (\labels[5][4] , \labels[5].delimiter[4] );
tran (\labels[5][5] , \labels[5].delimiter[5] );
tran (\labels[5][6] , \labels[5].delimiter[6] );
tran (\labels[5][7] , \labels[5].delimiter[7] );
tran (\labels[5][8] , \labels[5].delimiter_valid[0] );
tran (\labels[5][9] , \labels[5].label[0] );
tran (\labels[5][10] , \labels[5].label[1] );
tran (\labels[5][11] , \labels[5].label[2] );
tran (\labels[5][12] , \labels[5].label[3] );
tran (\labels[5][13] , \labels[5].label[4] );
tran (\labels[5][14] , \labels[5].label[5] );
tran (\labels[5][15] , \labels[5].label[6] );
tran (\labels[5][16] , \labels[5].label[7] );
tran (\labels[5][17] , \labels[5].label[8] );
tran (\labels[5][18] , \labels[5].label[9] );
tran (\labels[5][19] , \labels[5].label[10] );
tran (\labels[5][20] , \labels[5].label[11] );
tran (\labels[5][21] , \labels[5].label[12] );
tran (\labels[5][22] , \labels[5].label[13] );
tran (\labels[5][23] , \labels[5].label[14] );
tran (\labels[5][24] , \labels[5].label[15] );
tran (\labels[5][25] , \labels[5].label[16] );
tran (\labels[5][26] , \labels[5].label[17] );
tran (\labels[5][27] , \labels[5].label[18] );
tran (\labels[5][28] , \labels[5].label[19] );
tran (\labels[5][29] , \labels[5].label[20] );
tran (\labels[5][30] , \labels[5].label[21] );
tran (\labels[5][31] , \labels[5].label[22] );
tran (\labels[5][32] , \labels[5].label[23] );
tran (\labels[5][33] , \labels[5].label[24] );
tran (\labels[5][34] , \labels[5].label[25] );
tran (\labels[5][35] , \labels[5].label[26] );
tran (\labels[5][36] , \labels[5].label[27] );
tran (\labels[5][37] , \labels[5].label[28] );
tran (\labels[5][38] , \labels[5].label[29] );
tran (\labels[5][39] , \labels[5].label[30] );
tran (\labels[5][40] , \labels[5].label[31] );
tran (\labels[5][41] , \labels[5].label[32] );
tran (\labels[5][42] , \labels[5].label[33] );
tran (\labels[5][43] , \labels[5].label[34] );
tran (\labels[5][44] , \labels[5].label[35] );
tran (\labels[5][45] , \labels[5].label[36] );
tran (\labels[5][46] , \labels[5].label[37] );
tran (\labels[5][47] , \labels[5].label[38] );
tran (\labels[5][48] , \labels[5].label[39] );
tran (\labels[5][49] , \labels[5].label[40] );
tran (\labels[5][50] , \labels[5].label[41] );
tran (\labels[5][51] , \labels[5].label[42] );
tran (\labels[5][52] , \labels[5].label[43] );
tran (\labels[5][53] , \labels[5].label[44] );
tran (\labels[5][54] , \labels[5].label[45] );
tran (\labels[5][55] , \labels[5].label[46] );
tran (\labels[5][56] , \labels[5].label[47] );
tran (\labels[5][57] , \labels[5].label[48] );
tran (\labels[5][58] , \labels[5].label[49] );
tran (\labels[5][59] , \labels[5].label[50] );
tran (\labels[5][60] , \labels[5].label[51] );
tran (\labels[5][61] , \labels[5].label[52] );
tran (\labels[5][62] , \labels[5].label[53] );
tran (\labels[5][63] , \labels[5].label[54] );
tran (\labels[5][64] , \labels[5].label[55] );
tran (\labels[5][65] , \labels[5].label[56] );
tran (\labels[5][66] , \labels[5].label[57] );
tran (\labels[5][67] , \labels[5].label[58] );
tran (\labels[5][68] , \labels[5].label[59] );
tran (\labels[5][69] , \labels[5].label[60] );
tran (\labels[5][70] , \labels[5].label[61] );
tran (\labels[5][71] , \labels[5].label[62] );
tran (\labels[5][72] , \labels[5].label[63] );
tran (\labels[5][73] , \labels[5].label[64] );
tran (\labels[5][74] , \labels[5].label[65] );
tran (\labels[5][75] , \labels[5].label[66] );
tran (\labels[5][76] , \labels[5].label[67] );
tran (\labels[5][77] , \labels[5].label[68] );
tran (\labels[5][78] , \labels[5].label[69] );
tran (\labels[5][79] , \labels[5].label[70] );
tran (\labels[5][80] , \labels[5].label[71] );
tran (\labels[5][81] , \labels[5].label[72] );
tran (\labels[5][82] , \labels[5].label[73] );
tran (\labels[5][83] , \labels[5].label[74] );
tran (\labels[5][84] , \labels[5].label[75] );
tran (\labels[5][85] , \labels[5].label[76] );
tran (\labels[5][86] , \labels[5].label[77] );
tran (\labels[5][87] , \labels[5].label[78] );
tran (\labels[5][88] , \labels[5].label[79] );
tran (\labels[5][89] , \labels[5].label[80] );
tran (\labels[5][90] , \labels[5].label[81] );
tran (\labels[5][91] , \labels[5].label[82] );
tran (\labels[5][92] , \labels[5].label[83] );
tran (\labels[5][93] , \labels[5].label[84] );
tran (\labels[5][94] , \labels[5].label[85] );
tran (\labels[5][95] , \labels[5].label[86] );
tran (\labels[5][96] , \labels[5].label[87] );
tran (\labels[5][97] , \labels[5].label[88] );
tran (\labels[5][98] , \labels[5].label[89] );
tran (\labels[5][99] , \labels[5].label[90] );
tran (\labels[5][100] , \labels[5].label[91] );
tran (\labels[5][101] , \labels[5].label[92] );
tran (\labels[5][102] , \labels[5].label[93] );
tran (\labels[5][103] , \labels[5].label[94] );
tran (\labels[5][104] , \labels[5].label[95] );
tran (\labels[5][105] , \labels[5].label[96] );
tran (\labels[5][106] , \labels[5].label[97] );
tran (\labels[5][107] , \labels[5].label[98] );
tran (\labels[5][108] , \labels[5].label[99] );
tran (\labels[5][109] , \labels[5].label[100] );
tran (\labels[5][110] , \labels[5].label[101] );
tran (\labels[5][111] , \labels[5].label[102] );
tran (\labels[5][112] , \labels[5].label[103] );
tran (\labels[5][113] , \labels[5].label[104] );
tran (\labels[5][114] , \labels[5].label[105] );
tran (\labels[5][115] , \labels[5].label[106] );
tran (\labels[5][116] , \labels[5].label[107] );
tran (\labels[5][117] , \labels[5].label[108] );
tran (\labels[5][118] , \labels[5].label[109] );
tran (\labels[5][119] , \labels[5].label[110] );
tran (\labels[5][120] , \labels[5].label[111] );
tran (\labels[5][121] , \labels[5].label[112] );
tran (\labels[5][122] , \labels[5].label[113] );
tran (\labels[5][123] , \labels[5].label[114] );
tran (\labels[5][124] , \labels[5].label[115] );
tran (\labels[5][125] , \labels[5].label[116] );
tran (\labels[5][126] , \labels[5].label[117] );
tran (\labels[5][127] , \labels[5].label[118] );
tran (\labels[5][128] , \labels[5].label[119] );
tran (\labels[5][129] , \labels[5].label[120] );
tran (\labels[5][130] , \labels[5].label[121] );
tran (\labels[5][131] , \labels[5].label[122] );
tran (\labels[5][132] , \labels[5].label[123] );
tran (\labels[5][133] , \labels[5].label[124] );
tran (\labels[5][134] , \labels[5].label[125] );
tran (\labels[5][135] , \labels[5].label[126] );
tran (\labels[5][136] , \labels[5].label[127] );
tran (\labels[5][137] , \labels[5].label[128] );
tran (\labels[5][138] , \labels[5].label[129] );
tran (\labels[5][139] , \labels[5].label[130] );
tran (\labels[5][140] , \labels[5].label[131] );
tran (\labels[5][141] , \labels[5].label[132] );
tran (\labels[5][142] , \labels[5].label[133] );
tran (\labels[5][143] , \labels[5].label[134] );
tran (\labels[5][144] , \labels[5].label[135] );
tran (\labels[5][145] , \labels[5].label[136] );
tran (\labels[5][146] , \labels[5].label[137] );
tran (\labels[5][147] , \labels[5].label[138] );
tran (\labels[5][148] , \labels[5].label[139] );
tran (\labels[5][149] , \labels[5].label[140] );
tran (\labels[5][150] , \labels[5].label[141] );
tran (\labels[5][151] , \labels[5].label[142] );
tran (\labels[5][152] , \labels[5].label[143] );
tran (\labels[5][153] , \labels[5].label[144] );
tran (\labels[5][154] , \labels[5].label[145] );
tran (\labels[5][155] , \labels[5].label[146] );
tran (\labels[5][156] , \labels[5].label[147] );
tran (\labels[5][157] , \labels[5].label[148] );
tran (\labels[5][158] , \labels[5].label[149] );
tran (\labels[5][159] , \labels[5].label[150] );
tran (\labels[5][160] , \labels[5].label[151] );
tran (\labels[5][161] , \labels[5].label[152] );
tran (\labels[5][162] , \labels[5].label[153] );
tran (\labels[5][163] , \labels[5].label[154] );
tran (\labels[5][164] , \labels[5].label[155] );
tran (\labels[5][165] , \labels[5].label[156] );
tran (\labels[5][166] , \labels[5].label[157] );
tran (\labels[5][167] , \labels[5].label[158] );
tran (\labels[5][168] , \labels[5].label[159] );
tran (\labels[5][169] , \labels[5].label[160] );
tran (\labels[5][170] , \labels[5].label[161] );
tran (\labels[5][171] , \labels[5].label[162] );
tran (\labels[5][172] , \labels[5].label[163] );
tran (\labels[5][173] , \labels[5].label[164] );
tran (\labels[5][174] , \labels[5].label[165] );
tran (\labels[5][175] , \labels[5].label[166] );
tran (\labels[5][176] , \labels[5].label[167] );
tran (\labels[5][177] , \labels[5].label[168] );
tran (\labels[5][178] , \labels[5].label[169] );
tran (\labels[5][179] , \labels[5].label[170] );
tran (\labels[5][180] , \labels[5].label[171] );
tran (\labels[5][181] , \labels[5].label[172] );
tran (\labels[5][182] , \labels[5].label[173] );
tran (\labels[5][183] , \labels[5].label[174] );
tran (\labels[5][184] , \labels[5].label[175] );
tran (\labels[5][185] , \labels[5].label[176] );
tran (\labels[5][186] , \labels[5].label[177] );
tran (\labels[5][187] , \labels[5].label[178] );
tran (\labels[5][188] , \labels[5].label[179] );
tran (\labels[5][189] , \labels[5].label[180] );
tran (\labels[5][190] , \labels[5].label[181] );
tran (\labels[5][191] , \labels[5].label[182] );
tran (\labels[5][192] , \labels[5].label[183] );
tran (\labels[5][193] , \labels[5].label[184] );
tran (\labels[5][194] , \labels[5].label[185] );
tran (\labels[5][195] , \labels[5].label[186] );
tran (\labels[5][196] , \labels[5].label[187] );
tran (\labels[5][197] , \labels[5].label[188] );
tran (\labels[5][198] , \labels[5].label[189] );
tran (\labels[5][199] , \labels[5].label[190] );
tran (\labels[5][200] , \labels[5].label[191] );
tran (\labels[5][201] , \labels[5].label[192] );
tran (\labels[5][202] , \labels[5].label[193] );
tran (\labels[5][203] , \labels[5].label[194] );
tran (\labels[5][204] , \labels[5].label[195] );
tran (\labels[5][205] , \labels[5].label[196] );
tran (\labels[5][206] , \labels[5].label[197] );
tran (\labels[5][207] , \labels[5].label[198] );
tran (\labels[5][208] , \labels[5].label[199] );
tran (\labels[5][209] , \labels[5].label[200] );
tran (\labels[5][210] , \labels[5].label[201] );
tran (\labels[5][211] , \labels[5].label[202] );
tran (\labels[5][212] , \labels[5].label[203] );
tran (\labels[5][213] , \labels[5].label[204] );
tran (\labels[5][214] , \labels[5].label[205] );
tran (\labels[5][215] , \labels[5].label[206] );
tran (\labels[5][216] , \labels[5].label[207] );
tran (\labels[5][217] , \labels[5].label[208] );
tran (\labels[5][218] , \labels[5].label[209] );
tran (\labels[5][219] , \labels[5].label[210] );
tran (\labels[5][220] , \labels[5].label[211] );
tran (\labels[5][221] , \labels[5].label[212] );
tran (\labels[5][222] , \labels[5].label[213] );
tran (\labels[5][223] , \labels[5].label[214] );
tran (\labels[5][224] , \labels[5].label[215] );
tran (\labels[5][225] , \labels[5].label[216] );
tran (\labels[5][226] , \labels[5].label[217] );
tran (\labels[5][227] , \labels[5].label[218] );
tran (\labels[5][228] , \labels[5].label[219] );
tran (\labels[5][229] , \labels[5].label[220] );
tran (\labels[5][230] , \labels[5].label[221] );
tran (\labels[5][231] , \labels[5].label[222] );
tran (\labels[5][232] , \labels[5].label[223] );
tran (\labels[5][233] , \labels[5].label[224] );
tran (\labels[5][234] , \labels[5].label[225] );
tran (\labels[5][235] , \labels[5].label[226] );
tran (\labels[5][236] , \labels[5].label[227] );
tran (\labels[5][237] , \labels[5].label[228] );
tran (\labels[5][238] , \labels[5].label[229] );
tran (\labels[5][239] , \labels[5].label[230] );
tran (\labels[5][240] , \labels[5].label[231] );
tran (\labels[5][241] , \labels[5].label[232] );
tran (\labels[5][242] , \labels[5].label[233] );
tran (\labels[5][243] , \labels[5].label[234] );
tran (\labels[5][244] , \labels[5].label[235] );
tran (\labels[5][245] , \labels[5].label[236] );
tran (\labels[5][246] , \labels[5].label[237] );
tran (\labels[5][247] , \labels[5].label[238] );
tran (\labels[5][248] , \labels[5].label[239] );
tran (\labels[5][249] , \labels[5].label[240] );
tran (\labels[5][250] , \labels[5].label[241] );
tran (\labels[5][251] , \labels[5].label[242] );
tran (\labels[5][252] , \labels[5].label[243] );
tran (\labels[5][253] , \labels[5].label[244] );
tran (\labels[5][254] , \labels[5].label[245] );
tran (\labels[5][255] , \labels[5].label[246] );
tran (\labels[5][256] , \labels[5].label[247] );
tran (\labels[5][257] , \labels[5].label[248] );
tran (\labels[5][258] , \labels[5].label[249] );
tran (\labels[5][259] , \labels[5].label[250] );
tran (\labels[5][260] , \labels[5].label[251] );
tran (\labels[5][261] , \labels[5].label[252] );
tran (\labels[5][262] , \labels[5].label[253] );
tran (\labels[5][263] , \labels[5].label[254] );
tran (\labels[5][264] , \labels[5].label[255] );
tran (\labels[5][265] , \labels[5].label_size[0] );
tran (\labels[5][266] , \labels[5].label_size[1] );
tran (\labels[5][267] , \labels[5].label_size[2] );
tran (\labels[5][268] , \labels[5].label_size[3] );
tran (\labels[5][269] , \labels[5].label_size[4] );
tran (\labels[5][270] , \labels[5].label_size[5] );
tran (\labels[5][271] , \labels[5].guid_size[0] );
tran (\labels[6][0] , \labels[6].delimiter[0] );
tran (\labels[6][1] , \labels[6].delimiter[1] );
tran (\labels[6][2] , \labels[6].delimiter[2] );
tran (\labels[6][3] , \labels[6].delimiter[3] );
tran (\labels[6][4] , \labels[6].delimiter[4] );
tran (\labels[6][5] , \labels[6].delimiter[5] );
tran (\labels[6][6] , \labels[6].delimiter[6] );
tran (\labels[6][7] , \labels[6].delimiter[7] );
tran (\labels[6][8] , \labels[6].delimiter_valid[0] );
tran (\labels[6][9] , \labels[6].label[0] );
tran (\labels[6][10] , \labels[6].label[1] );
tran (\labels[6][11] , \labels[6].label[2] );
tran (\labels[6][12] , \labels[6].label[3] );
tran (\labels[6][13] , \labels[6].label[4] );
tran (\labels[6][14] , \labels[6].label[5] );
tran (\labels[6][15] , \labels[6].label[6] );
tran (\labels[6][16] , \labels[6].label[7] );
tran (\labels[6][17] , \labels[6].label[8] );
tran (\labels[6][18] , \labels[6].label[9] );
tran (\labels[6][19] , \labels[6].label[10] );
tran (\labels[6][20] , \labels[6].label[11] );
tran (\labels[6][21] , \labels[6].label[12] );
tran (\labels[6][22] , \labels[6].label[13] );
tran (\labels[6][23] , \labels[6].label[14] );
tran (\labels[6][24] , \labels[6].label[15] );
tran (\labels[6][25] , \labels[6].label[16] );
tran (\labels[6][26] , \labels[6].label[17] );
tran (\labels[6][27] , \labels[6].label[18] );
tran (\labels[6][28] , \labels[6].label[19] );
tran (\labels[6][29] , \labels[6].label[20] );
tran (\labels[6][30] , \labels[6].label[21] );
tran (\labels[6][31] , \labels[6].label[22] );
tran (\labels[6][32] , \labels[6].label[23] );
tran (\labels[6][33] , \labels[6].label[24] );
tran (\labels[6][34] , \labels[6].label[25] );
tran (\labels[6][35] , \labels[6].label[26] );
tran (\labels[6][36] , \labels[6].label[27] );
tran (\labels[6][37] , \labels[6].label[28] );
tran (\labels[6][38] , \labels[6].label[29] );
tran (\labels[6][39] , \labels[6].label[30] );
tran (\labels[6][40] , \labels[6].label[31] );
tran (\labels[6][41] , \labels[6].label[32] );
tran (\labels[6][42] , \labels[6].label[33] );
tran (\labels[6][43] , \labels[6].label[34] );
tran (\labels[6][44] , \labels[6].label[35] );
tran (\labels[6][45] , \labels[6].label[36] );
tran (\labels[6][46] , \labels[6].label[37] );
tran (\labels[6][47] , \labels[6].label[38] );
tran (\labels[6][48] , \labels[6].label[39] );
tran (\labels[6][49] , \labels[6].label[40] );
tran (\labels[6][50] , \labels[6].label[41] );
tran (\labels[6][51] , \labels[6].label[42] );
tran (\labels[6][52] , \labels[6].label[43] );
tran (\labels[6][53] , \labels[6].label[44] );
tran (\labels[6][54] , \labels[6].label[45] );
tran (\labels[6][55] , \labels[6].label[46] );
tran (\labels[6][56] , \labels[6].label[47] );
tran (\labels[6][57] , \labels[6].label[48] );
tran (\labels[6][58] , \labels[6].label[49] );
tran (\labels[6][59] , \labels[6].label[50] );
tran (\labels[6][60] , \labels[6].label[51] );
tran (\labels[6][61] , \labels[6].label[52] );
tran (\labels[6][62] , \labels[6].label[53] );
tran (\labels[6][63] , \labels[6].label[54] );
tran (\labels[6][64] , \labels[6].label[55] );
tran (\labels[6][65] , \labels[6].label[56] );
tran (\labels[6][66] , \labels[6].label[57] );
tran (\labels[6][67] , \labels[6].label[58] );
tran (\labels[6][68] , \labels[6].label[59] );
tran (\labels[6][69] , \labels[6].label[60] );
tran (\labels[6][70] , \labels[6].label[61] );
tran (\labels[6][71] , \labels[6].label[62] );
tran (\labels[6][72] , \labels[6].label[63] );
tran (\labels[6][73] , \labels[6].label[64] );
tran (\labels[6][74] , \labels[6].label[65] );
tran (\labels[6][75] , \labels[6].label[66] );
tran (\labels[6][76] , \labels[6].label[67] );
tran (\labels[6][77] , \labels[6].label[68] );
tran (\labels[6][78] , \labels[6].label[69] );
tran (\labels[6][79] , \labels[6].label[70] );
tran (\labels[6][80] , \labels[6].label[71] );
tran (\labels[6][81] , \labels[6].label[72] );
tran (\labels[6][82] , \labels[6].label[73] );
tran (\labels[6][83] , \labels[6].label[74] );
tran (\labels[6][84] , \labels[6].label[75] );
tran (\labels[6][85] , \labels[6].label[76] );
tran (\labels[6][86] , \labels[6].label[77] );
tran (\labels[6][87] , \labels[6].label[78] );
tran (\labels[6][88] , \labels[6].label[79] );
tran (\labels[6][89] , \labels[6].label[80] );
tran (\labels[6][90] , \labels[6].label[81] );
tran (\labels[6][91] , \labels[6].label[82] );
tran (\labels[6][92] , \labels[6].label[83] );
tran (\labels[6][93] , \labels[6].label[84] );
tran (\labels[6][94] , \labels[6].label[85] );
tran (\labels[6][95] , \labels[6].label[86] );
tran (\labels[6][96] , \labels[6].label[87] );
tran (\labels[6][97] , \labels[6].label[88] );
tran (\labels[6][98] , \labels[6].label[89] );
tran (\labels[6][99] , \labels[6].label[90] );
tran (\labels[6][100] , \labels[6].label[91] );
tran (\labels[6][101] , \labels[6].label[92] );
tran (\labels[6][102] , \labels[6].label[93] );
tran (\labels[6][103] , \labels[6].label[94] );
tran (\labels[6][104] , \labels[6].label[95] );
tran (\labels[6][105] , \labels[6].label[96] );
tran (\labels[6][106] , \labels[6].label[97] );
tran (\labels[6][107] , \labels[6].label[98] );
tran (\labels[6][108] , \labels[6].label[99] );
tran (\labels[6][109] , \labels[6].label[100] );
tran (\labels[6][110] , \labels[6].label[101] );
tran (\labels[6][111] , \labels[6].label[102] );
tran (\labels[6][112] , \labels[6].label[103] );
tran (\labels[6][113] , \labels[6].label[104] );
tran (\labels[6][114] , \labels[6].label[105] );
tran (\labels[6][115] , \labels[6].label[106] );
tran (\labels[6][116] , \labels[6].label[107] );
tran (\labels[6][117] , \labels[6].label[108] );
tran (\labels[6][118] , \labels[6].label[109] );
tran (\labels[6][119] , \labels[6].label[110] );
tran (\labels[6][120] , \labels[6].label[111] );
tran (\labels[6][121] , \labels[6].label[112] );
tran (\labels[6][122] , \labels[6].label[113] );
tran (\labels[6][123] , \labels[6].label[114] );
tran (\labels[6][124] , \labels[6].label[115] );
tran (\labels[6][125] , \labels[6].label[116] );
tran (\labels[6][126] , \labels[6].label[117] );
tran (\labels[6][127] , \labels[6].label[118] );
tran (\labels[6][128] , \labels[6].label[119] );
tran (\labels[6][129] , \labels[6].label[120] );
tran (\labels[6][130] , \labels[6].label[121] );
tran (\labels[6][131] , \labels[6].label[122] );
tran (\labels[6][132] , \labels[6].label[123] );
tran (\labels[6][133] , \labels[6].label[124] );
tran (\labels[6][134] , \labels[6].label[125] );
tran (\labels[6][135] , \labels[6].label[126] );
tran (\labels[6][136] , \labels[6].label[127] );
tran (\labels[6][137] , \labels[6].label[128] );
tran (\labels[6][138] , \labels[6].label[129] );
tran (\labels[6][139] , \labels[6].label[130] );
tran (\labels[6][140] , \labels[6].label[131] );
tran (\labels[6][141] , \labels[6].label[132] );
tran (\labels[6][142] , \labels[6].label[133] );
tran (\labels[6][143] , \labels[6].label[134] );
tran (\labels[6][144] , \labels[6].label[135] );
tran (\labels[6][145] , \labels[6].label[136] );
tran (\labels[6][146] , \labels[6].label[137] );
tran (\labels[6][147] , \labels[6].label[138] );
tran (\labels[6][148] , \labels[6].label[139] );
tran (\labels[6][149] , \labels[6].label[140] );
tran (\labels[6][150] , \labels[6].label[141] );
tran (\labels[6][151] , \labels[6].label[142] );
tran (\labels[6][152] , \labels[6].label[143] );
tran (\labels[6][153] , \labels[6].label[144] );
tran (\labels[6][154] , \labels[6].label[145] );
tran (\labels[6][155] , \labels[6].label[146] );
tran (\labels[6][156] , \labels[6].label[147] );
tran (\labels[6][157] , \labels[6].label[148] );
tran (\labels[6][158] , \labels[6].label[149] );
tran (\labels[6][159] , \labels[6].label[150] );
tran (\labels[6][160] , \labels[6].label[151] );
tran (\labels[6][161] , \labels[6].label[152] );
tran (\labels[6][162] , \labels[6].label[153] );
tran (\labels[6][163] , \labels[6].label[154] );
tran (\labels[6][164] , \labels[6].label[155] );
tran (\labels[6][165] , \labels[6].label[156] );
tran (\labels[6][166] , \labels[6].label[157] );
tran (\labels[6][167] , \labels[6].label[158] );
tran (\labels[6][168] , \labels[6].label[159] );
tran (\labels[6][169] , \labels[6].label[160] );
tran (\labels[6][170] , \labels[6].label[161] );
tran (\labels[6][171] , \labels[6].label[162] );
tran (\labels[6][172] , \labels[6].label[163] );
tran (\labels[6][173] , \labels[6].label[164] );
tran (\labels[6][174] , \labels[6].label[165] );
tran (\labels[6][175] , \labels[6].label[166] );
tran (\labels[6][176] , \labels[6].label[167] );
tran (\labels[6][177] , \labels[6].label[168] );
tran (\labels[6][178] , \labels[6].label[169] );
tran (\labels[6][179] , \labels[6].label[170] );
tran (\labels[6][180] , \labels[6].label[171] );
tran (\labels[6][181] , \labels[6].label[172] );
tran (\labels[6][182] , \labels[6].label[173] );
tran (\labels[6][183] , \labels[6].label[174] );
tran (\labels[6][184] , \labels[6].label[175] );
tran (\labels[6][185] , \labels[6].label[176] );
tran (\labels[6][186] , \labels[6].label[177] );
tran (\labels[6][187] , \labels[6].label[178] );
tran (\labels[6][188] , \labels[6].label[179] );
tran (\labels[6][189] , \labels[6].label[180] );
tran (\labels[6][190] , \labels[6].label[181] );
tran (\labels[6][191] , \labels[6].label[182] );
tran (\labels[6][192] , \labels[6].label[183] );
tran (\labels[6][193] , \labels[6].label[184] );
tran (\labels[6][194] , \labels[6].label[185] );
tran (\labels[6][195] , \labels[6].label[186] );
tran (\labels[6][196] , \labels[6].label[187] );
tran (\labels[6][197] , \labels[6].label[188] );
tran (\labels[6][198] , \labels[6].label[189] );
tran (\labels[6][199] , \labels[6].label[190] );
tran (\labels[6][200] , \labels[6].label[191] );
tran (\labels[6][201] , \labels[6].label[192] );
tran (\labels[6][202] , \labels[6].label[193] );
tran (\labels[6][203] , \labels[6].label[194] );
tran (\labels[6][204] , \labels[6].label[195] );
tran (\labels[6][205] , \labels[6].label[196] );
tran (\labels[6][206] , \labels[6].label[197] );
tran (\labels[6][207] , \labels[6].label[198] );
tran (\labels[6][208] , \labels[6].label[199] );
tran (\labels[6][209] , \labels[6].label[200] );
tran (\labels[6][210] , \labels[6].label[201] );
tran (\labels[6][211] , \labels[6].label[202] );
tran (\labels[6][212] , \labels[6].label[203] );
tran (\labels[6][213] , \labels[6].label[204] );
tran (\labels[6][214] , \labels[6].label[205] );
tran (\labels[6][215] , \labels[6].label[206] );
tran (\labels[6][216] , \labels[6].label[207] );
tran (\labels[6][217] , \labels[6].label[208] );
tran (\labels[6][218] , \labels[6].label[209] );
tran (\labels[6][219] , \labels[6].label[210] );
tran (\labels[6][220] , \labels[6].label[211] );
tran (\labels[6][221] , \labels[6].label[212] );
tran (\labels[6][222] , \labels[6].label[213] );
tran (\labels[6][223] , \labels[6].label[214] );
tran (\labels[6][224] , \labels[6].label[215] );
tran (\labels[6][225] , \labels[6].label[216] );
tran (\labels[6][226] , \labels[6].label[217] );
tran (\labels[6][227] , \labels[6].label[218] );
tran (\labels[6][228] , \labels[6].label[219] );
tran (\labels[6][229] , \labels[6].label[220] );
tran (\labels[6][230] , \labels[6].label[221] );
tran (\labels[6][231] , \labels[6].label[222] );
tran (\labels[6][232] , \labels[6].label[223] );
tran (\labels[6][233] , \labels[6].label[224] );
tran (\labels[6][234] , \labels[6].label[225] );
tran (\labels[6][235] , \labels[6].label[226] );
tran (\labels[6][236] , \labels[6].label[227] );
tran (\labels[6][237] , \labels[6].label[228] );
tran (\labels[6][238] , \labels[6].label[229] );
tran (\labels[6][239] , \labels[6].label[230] );
tran (\labels[6][240] , \labels[6].label[231] );
tran (\labels[6][241] , \labels[6].label[232] );
tran (\labels[6][242] , \labels[6].label[233] );
tran (\labels[6][243] , \labels[6].label[234] );
tran (\labels[6][244] , \labels[6].label[235] );
tran (\labels[6][245] , \labels[6].label[236] );
tran (\labels[6][246] , \labels[6].label[237] );
tran (\labels[6][247] , \labels[6].label[238] );
tran (\labels[6][248] , \labels[6].label[239] );
tran (\labels[6][249] , \labels[6].label[240] );
tran (\labels[6][250] , \labels[6].label[241] );
tran (\labels[6][251] , \labels[6].label[242] );
tran (\labels[6][252] , \labels[6].label[243] );
tran (\labels[6][253] , \labels[6].label[244] );
tran (\labels[6][254] , \labels[6].label[245] );
tran (\labels[6][255] , \labels[6].label[246] );
tran (\labels[6][256] , \labels[6].label[247] );
tran (\labels[6][257] , \labels[6].label[248] );
tran (\labels[6][258] , \labels[6].label[249] );
tran (\labels[6][259] , \labels[6].label[250] );
tran (\labels[6][260] , \labels[6].label[251] );
tran (\labels[6][261] , \labels[6].label[252] );
tran (\labels[6][262] , \labels[6].label[253] );
tran (\labels[6][263] , \labels[6].label[254] );
tran (\labels[6][264] , \labels[6].label[255] );
tran (\labels[6][265] , \labels[6].label_size[0] );
tran (\labels[6][266] , \labels[6].label_size[1] );
tran (\labels[6][267] , \labels[6].label_size[2] );
tran (\labels[6][268] , \labels[6].label_size[3] );
tran (\labels[6][269] , \labels[6].label_size[4] );
tran (\labels[6][270] , \labels[6].label_size[5] );
tran (\labels[6][271] , \labels[6].guid_size[0] );
tran (\labels[7][0] , \labels[7].delimiter[0] );
tran (\labels[7][1] , \labels[7].delimiter[1] );
tran (\labels[7][2] , \labels[7].delimiter[2] );
tran (\labels[7][3] , \labels[7].delimiter[3] );
tran (\labels[7][4] , \labels[7].delimiter[4] );
tran (\labels[7][5] , \labels[7].delimiter[5] );
tran (\labels[7][6] , \labels[7].delimiter[6] );
tran (\labels[7][7] , \labels[7].delimiter[7] );
tran (\labels[7][8] , \labels[7].delimiter_valid[0] );
tran (\labels[7][9] , \labels[7].label[0] );
tran (\labels[7][10] , \labels[7].label[1] );
tran (\labels[7][11] , \labels[7].label[2] );
tran (\labels[7][12] , \labels[7].label[3] );
tran (\labels[7][13] , \labels[7].label[4] );
tran (\labels[7][14] , \labels[7].label[5] );
tran (\labels[7][15] , \labels[7].label[6] );
tran (\labels[7][16] , \labels[7].label[7] );
tran (\labels[7][17] , \labels[7].label[8] );
tran (\labels[7][18] , \labels[7].label[9] );
tran (\labels[7][19] , \labels[7].label[10] );
tran (\labels[7][20] , \labels[7].label[11] );
tran (\labels[7][21] , \labels[7].label[12] );
tran (\labels[7][22] , \labels[7].label[13] );
tran (\labels[7][23] , \labels[7].label[14] );
tran (\labels[7][24] , \labels[7].label[15] );
tran (\labels[7][25] , \labels[7].label[16] );
tran (\labels[7][26] , \labels[7].label[17] );
tran (\labels[7][27] , \labels[7].label[18] );
tran (\labels[7][28] , \labels[7].label[19] );
tran (\labels[7][29] , \labels[7].label[20] );
tran (\labels[7][30] , \labels[7].label[21] );
tran (\labels[7][31] , \labels[7].label[22] );
tran (\labels[7][32] , \labels[7].label[23] );
tran (\labels[7][33] , \labels[7].label[24] );
tran (\labels[7][34] , \labels[7].label[25] );
tran (\labels[7][35] , \labels[7].label[26] );
tran (\labels[7][36] , \labels[7].label[27] );
tran (\labels[7][37] , \labels[7].label[28] );
tran (\labels[7][38] , \labels[7].label[29] );
tran (\labels[7][39] , \labels[7].label[30] );
tran (\labels[7][40] , \labels[7].label[31] );
tran (\labels[7][41] , \labels[7].label[32] );
tran (\labels[7][42] , \labels[7].label[33] );
tran (\labels[7][43] , \labels[7].label[34] );
tran (\labels[7][44] , \labels[7].label[35] );
tran (\labels[7][45] , \labels[7].label[36] );
tran (\labels[7][46] , \labels[7].label[37] );
tran (\labels[7][47] , \labels[7].label[38] );
tran (\labels[7][48] , \labels[7].label[39] );
tran (\labels[7][49] , \labels[7].label[40] );
tran (\labels[7][50] , \labels[7].label[41] );
tran (\labels[7][51] , \labels[7].label[42] );
tran (\labels[7][52] , \labels[7].label[43] );
tran (\labels[7][53] , \labels[7].label[44] );
tran (\labels[7][54] , \labels[7].label[45] );
tran (\labels[7][55] , \labels[7].label[46] );
tran (\labels[7][56] , \labels[7].label[47] );
tran (\labels[7][57] , \labels[7].label[48] );
tran (\labels[7][58] , \labels[7].label[49] );
tran (\labels[7][59] , \labels[7].label[50] );
tran (\labels[7][60] , \labels[7].label[51] );
tran (\labels[7][61] , \labels[7].label[52] );
tran (\labels[7][62] , \labels[7].label[53] );
tran (\labels[7][63] , \labels[7].label[54] );
tran (\labels[7][64] , \labels[7].label[55] );
tran (\labels[7][65] , \labels[7].label[56] );
tran (\labels[7][66] , \labels[7].label[57] );
tran (\labels[7][67] , \labels[7].label[58] );
tran (\labels[7][68] , \labels[7].label[59] );
tran (\labels[7][69] , \labels[7].label[60] );
tran (\labels[7][70] , \labels[7].label[61] );
tran (\labels[7][71] , \labels[7].label[62] );
tran (\labels[7][72] , \labels[7].label[63] );
tran (\labels[7][73] , \labels[7].label[64] );
tran (\labels[7][74] , \labels[7].label[65] );
tran (\labels[7][75] , \labels[7].label[66] );
tran (\labels[7][76] , \labels[7].label[67] );
tran (\labels[7][77] , \labels[7].label[68] );
tran (\labels[7][78] , \labels[7].label[69] );
tran (\labels[7][79] , \labels[7].label[70] );
tran (\labels[7][80] , \labels[7].label[71] );
tran (\labels[7][81] , \labels[7].label[72] );
tran (\labels[7][82] , \labels[7].label[73] );
tran (\labels[7][83] , \labels[7].label[74] );
tran (\labels[7][84] , \labels[7].label[75] );
tran (\labels[7][85] , \labels[7].label[76] );
tran (\labels[7][86] , \labels[7].label[77] );
tran (\labels[7][87] , \labels[7].label[78] );
tran (\labels[7][88] , \labels[7].label[79] );
tran (\labels[7][89] , \labels[7].label[80] );
tran (\labels[7][90] , \labels[7].label[81] );
tran (\labels[7][91] , \labels[7].label[82] );
tran (\labels[7][92] , \labels[7].label[83] );
tran (\labels[7][93] , \labels[7].label[84] );
tran (\labels[7][94] , \labels[7].label[85] );
tran (\labels[7][95] , \labels[7].label[86] );
tran (\labels[7][96] , \labels[7].label[87] );
tran (\labels[7][97] , \labels[7].label[88] );
tran (\labels[7][98] , \labels[7].label[89] );
tran (\labels[7][99] , \labels[7].label[90] );
tran (\labels[7][100] , \labels[7].label[91] );
tran (\labels[7][101] , \labels[7].label[92] );
tran (\labels[7][102] , \labels[7].label[93] );
tran (\labels[7][103] , \labels[7].label[94] );
tran (\labels[7][104] , \labels[7].label[95] );
tran (\labels[7][105] , \labels[7].label[96] );
tran (\labels[7][106] , \labels[7].label[97] );
tran (\labels[7][107] , \labels[7].label[98] );
tran (\labels[7][108] , \labels[7].label[99] );
tran (\labels[7][109] , \labels[7].label[100] );
tran (\labels[7][110] , \labels[7].label[101] );
tran (\labels[7][111] , \labels[7].label[102] );
tran (\labels[7][112] , \labels[7].label[103] );
tran (\labels[7][113] , \labels[7].label[104] );
tran (\labels[7][114] , \labels[7].label[105] );
tran (\labels[7][115] , \labels[7].label[106] );
tran (\labels[7][116] , \labels[7].label[107] );
tran (\labels[7][117] , \labels[7].label[108] );
tran (\labels[7][118] , \labels[7].label[109] );
tran (\labels[7][119] , \labels[7].label[110] );
tran (\labels[7][120] , \labels[7].label[111] );
tran (\labels[7][121] , \labels[7].label[112] );
tran (\labels[7][122] , \labels[7].label[113] );
tran (\labels[7][123] , \labels[7].label[114] );
tran (\labels[7][124] , \labels[7].label[115] );
tran (\labels[7][125] , \labels[7].label[116] );
tran (\labels[7][126] , \labels[7].label[117] );
tran (\labels[7][127] , \labels[7].label[118] );
tran (\labels[7][128] , \labels[7].label[119] );
tran (\labels[7][129] , \labels[7].label[120] );
tran (\labels[7][130] , \labels[7].label[121] );
tran (\labels[7][131] , \labels[7].label[122] );
tran (\labels[7][132] , \labels[7].label[123] );
tran (\labels[7][133] , \labels[7].label[124] );
tran (\labels[7][134] , \labels[7].label[125] );
tran (\labels[7][135] , \labels[7].label[126] );
tran (\labels[7][136] , \labels[7].label[127] );
tran (\labels[7][137] , \labels[7].label[128] );
tran (\labels[7][138] , \labels[7].label[129] );
tran (\labels[7][139] , \labels[7].label[130] );
tran (\labels[7][140] , \labels[7].label[131] );
tran (\labels[7][141] , \labels[7].label[132] );
tran (\labels[7][142] , \labels[7].label[133] );
tran (\labels[7][143] , \labels[7].label[134] );
tran (\labels[7][144] , \labels[7].label[135] );
tran (\labels[7][145] , \labels[7].label[136] );
tran (\labels[7][146] , \labels[7].label[137] );
tran (\labels[7][147] , \labels[7].label[138] );
tran (\labels[7][148] , \labels[7].label[139] );
tran (\labels[7][149] , \labels[7].label[140] );
tran (\labels[7][150] , \labels[7].label[141] );
tran (\labels[7][151] , \labels[7].label[142] );
tran (\labels[7][152] , \labels[7].label[143] );
tran (\labels[7][153] , \labels[7].label[144] );
tran (\labels[7][154] , \labels[7].label[145] );
tran (\labels[7][155] , \labels[7].label[146] );
tran (\labels[7][156] , \labels[7].label[147] );
tran (\labels[7][157] , \labels[7].label[148] );
tran (\labels[7][158] , \labels[7].label[149] );
tran (\labels[7][159] , \labels[7].label[150] );
tran (\labels[7][160] , \labels[7].label[151] );
tran (\labels[7][161] , \labels[7].label[152] );
tran (\labels[7][162] , \labels[7].label[153] );
tran (\labels[7][163] , \labels[7].label[154] );
tran (\labels[7][164] , \labels[7].label[155] );
tran (\labels[7][165] , \labels[7].label[156] );
tran (\labels[7][166] , \labels[7].label[157] );
tran (\labels[7][167] , \labels[7].label[158] );
tran (\labels[7][168] , \labels[7].label[159] );
tran (\labels[7][169] , \labels[7].label[160] );
tran (\labels[7][170] , \labels[7].label[161] );
tran (\labels[7][171] , \labels[7].label[162] );
tran (\labels[7][172] , \labels[7].label[163] );
tran (\labels[7][173] , \labels[7].label[164] );
tran (\labels[7][174] , \labels[7].label[165] );
tran (\labels[7][175] , \labels[7].label[166] );
tran (\labels[7][176] , \labels[7].label[167] );
tran (\labels[7][177] , \labels[7].label[168] );
tran (\labels[7][178] , \labels[7].label[169] );
tran (\labels[7][179] , \labels[7].label[170] );
tran (\labels[7][180] , \labels[7].label[171] );
tran (\labels[7][181] , \labels[7].label[172] );
tran (\labels[7][182] , \labels[7].label[173] );
tran (\labels[7][183] , \labels[7].label[174] );
tran (\labels[7][184] , \labels[7].label[175] );
tran (\labels[7][185] , \labels[7].label[176] );
tran (\labels[7][186] , \labels[7].label[177] );
tran (\labels[7][187] , \labels[7].label[178] );
tran (\labels[7][188] , \labels[7].label[179] );
tran (\labels[7][189] , \labels[7].label[180] );
tran (\labels[7][190] , \labels[7].label[181] );
tran (\labels[7][191] , \labels[7].label[182] );
tran (\labels[7][192] , \labels[7].label[183] );
tran (\labels[7][193] , \labels[7].label[184] );
tran (\labels[7][194] , \labels[7].label[185] );
tran (\labels[7][195] , \labels[7].label[186] );
tran (\labels[7][196] , \labels[7].label[187] );
tran (\labels[7][197] , \labels[7].label[188] );
tran (\labels[7][198] , \labels[7].label[189] );
tran (\labels[7][199] , \labels[7].label[190] );
tran (\labels[7][200] , \labels[7].label[191] );
tran (\labels[7][201] , \labels[7].label[192] );
tran (\labels[7][202] , \labels[7].label[193] );
tran (\labels[7][203] , \labels[7].label[194] );
tran (\labels[7][204] , \labels[7].label[195] );
tran (\labels[7][205] , \labels[7].label[196] );
tran (\labels[7][206] , \labels[7].label[197] );
tran (\labels[7][207] , \labels[7].label[198] );
tran (\labels[7][208] , \labels[7].label[199] );
tran (\labels[7][209] , \labels[7].label[200] );
tran (\labels[7][210] , \labels[7].label[201] );
tran (\labels[7][211] , \labels[7].label[202] );
tran (\labels[7][212] , \labels[7].label[203] );
tran (\labels[7][213] , \labels[7].label[204] );
tran (\labels[7][214] , \labels[7].label[205] );
tran (\labels[7][215] , \labels[7].label[206] );
tran (\labels[7][216] , \labels[7].label[207] );
tran (\labels[7][217] , \labels[7].label[208] );
tran (\labels[7][218] , \labels[7].label[209] );
tran (\labels[7][219] , \labels[7].label[210] );
tran (\labels[7][220] , \labels[7].label[211] );
tran (\labels[7][221] , \labels[7].label[212] );
tran (\labels[7][222] , \labels[7].label[213] );
tran (\labels[7][223] , \labels[7].label[214] );
tran (\labels[7][224] , \labels[7].label[215] );
tran (\labels[7][225] , \labels[7].label[216] );
tran (\labels[7][226] , \labels[7].label[217] );
tran (\labels[7][227] , \labels[7].label[218] );
tran (\labels[7][228] , \labels[7].label[219] );
tran (\labels[7][229] , \labels[7].label[220] );
tran (\labels[7][230] , \labels[7].label[221] );
tran (\labels[7][231] , \labels[7].label[222] );
tran (\labels[7][232] , \labels[7].label[223] );
tran (\labels[7][233] , \labels[7].label[224] );
tran (\labels[7][234] , \labels[7].label[225] );
tran (\labels[7][235] , \labels[7].label[226] );
tran (\labels[7][236] , \labels[7].label[227] );
tran (\labels[7][237] , \labels[7].label[228] );
tran (\labels[7][238] , \labels[7].label[229] );
tran (\labels[7][239] , \labels[7].label[230] );
tran (\labels[7][240] , \labels[7].label[231] );
tran (\labels[7][241] , \labels[7].label[232] );
tran (\labels[7][242] , \labels[7].label[233] );
tran (\labels[7][243] , \labels[7].label[234] );
tran (\labels[7][244] , \labels[7].label[235] );
tran (\labels[7][245] , \labels[7].label[236] );
tran (\labels[7][246] , \labels[7].label[237] );
tran (\labels[7][247] , \labels[7].label[238] );
tran (\labels[7][248] , \labels[7].label[239] );
tran (\labels[7][249] , \labels[7].label[240] );
tran (\labels[7][250] , \labels[7].label[241] );
tran (\labels[7][251] , \labels[7].label[242] );
tran (\labels[7][252] , \labels[7].label[243] );
tran (\labels[7][253] , \labels[7].label[244] );
tran (\labels[7][254] , \labels[7].label[245] );
tran (\labels[7][255] , \labels[7].label[246] );
tran (\labels[7][256] , \labels[7].label[247] );
tran (\labels[7][257] , \labels[7].label[248] );
tran (\labels[7][258] , \labels[7].label[249] );
tran (\labels[7][259] , \labels[7].label[250] );
tran (\labels[7][260] , \labels[7].label[251] );
tran (\labels[7][261] , \labels[7].label[252] );
tran (\labels[7][262] , \labels[7].label[253] );
tran (\labels[7][263] , \labels[7].label[254] );
tran (\labels[7][264] , \labels[7].label[255] );
tran (\labels[7][265] , \labels[7].label_size[0] );
tran (\labels[7][266] , \labels[7].label_size[1] );
tran (\labels[7][267] , \labels[7].label_size[2] );
tran (\labels[7][268] , \labels[7].label_size[3] );
tran (\labels[7][269] , \labels[7].label_size[4] );
tran (\labels[7][270] , \labels[7].label_size[5] );
tran (\labels[7][271] , \labels[7].guid_size[0] );
tran (tready_override[8], \tready_override.r.part0 [8]);
tran (tready_override[8], \tready_override.f.txc_tready_override );
tran (tready_override[7], \tready_override.r.part0 [7]);
tran (tready_override[7], \tready_override.f.engine_7_tready_override );
tran (tready_override[6], \tready_override.r.part0 [6]);
tran (tready_override[6], \tready_override.f.engine_6_tready_override );
tran (tready_override[5], \tready_override.r.part0 [5]);
tran (tready_override[5], \tready_override.f.engine_5_tready_override );
tran (tready_override[4], \tready_override.r.part0 [4]);
tran (tready_override[4], \tready_override.f.engine_4_tready_override );
tran (tready_override[3], \tready_override.r.part0 [3]);
tran (tready_override[3], \tready_override.f.engine_3_tready_override );
tran (tready_override[2], \tready_override.r.part0 [2]);
tran (tready_override[2], \tready_override.f.engine_2_tready_override );
tran (tready_override[1], \tready_override.r.part0 [1]);
tran (tready_override[1], \tready_override.f.engine_1_tready_override );
tran (tready_override[0], \tready_override.r.part0 [0]);
tran (tready_override[0], \tready_override.f.engine_0_tready_override );
tran (cceip_encrypt_kop_fifo_override[6], \cceip_encrypt_kop_fifo_override.r.part0 [6]);
tran (cceip_encrypt_kop_fifo_override[6], \cceip_encrypt_kop_fifo_override.f.gcm_status_data_fifo );
tran (cceip_encrypt_kop_fifo_override[5], \cceip_encrypt_kop_fifo_override.r.part0 [5]);
tran (cceip_encrypt_kop_fifo_override[5], \cceip_encrypt_kop_fifo_override.f.tlv_sb_data_fifo );
tran (cceip_encrypt_kop_fifo_override[4], \cceip_encrypt_kop_fifo_override.r.part0 [4]);
tran (cceip_encrypt_kop_fifo_override[4], \cceip_encrypt_kop_fifo_override.f.kdf_cmd_fifo );
tran (cceip_encrypt_kop_fifo_override[3], \cceip_encrypt_kop_fifo_override.r.part0 [3]);
tran (cceip_encrypt_kop_fifo_override[3], \cceip_encrypt_kop_fifo_override.f.kdfstream_cmd_fifo );
tran (cceip_encrypt_kop_fifo_override[2], \cceip_encrypt_kop_fifo_override.r.part0 [2]);
tran (cceip_encrypt_kop_fifo_override[2], \cceip_encrypt_kop_fifo_override.f.keyfilter_cmd_fifo );
tran (cceip_encrypt_kop_fifo_override[1], \cceip_encrypt_kop_fifo_override.r.part0 [1]);
tran (cceip_encrypt_kop_fifo_override[1], \cceip_encrypt_kop_fifo_override.f.gcm_tag_data_fifo );
tran (cceip_encrypt_kop_fifo_override[0], \cceip_encrypt_kop_fifo_override.r.part0 [0]);
tran (cceip_encrypt_kop_fifo_override[0], \cceip_encrypt_kop_fifo_override.f.gcm_cmd_fifo );
tran (cceip_validate_kop_fifo_override[6], \cceip_validate_kop_fifo_override.r.part0 [6]);
tran (cceip_validate_kop_fifo_override[6], \cceip_validate_kop_fifo_override.f.gcm_status_data_fifo );
tran (cceip_validate_kop_fifo_override[5], \cceip_validate_kop_fifo_override.r.part0 [5]);
tran (cceip_validate_kop_fifo_override[5], \cceip_validate_kop_fifo_override.f.tlv_sb_data_fifo );
tran (cceip_validate_kop_fifo_override[4], \cceip_validate_kop_fifo_override.r.part0 [4]);
tran (cceip_validate_kop_fifo_override[4], \cceip_validate_kop_fifo_override.f.kdf_cmd_fifo );
tran (cceip_validate_kop_fifo_override[3], \cceip_validate_kop_fifo_override.r.part0 [3]);
tran (cceip_validate_kop_fifo_override[3], \cceip_validate_kop_fifo_override.f.kdfstream_cmd_fifo );
tran (cceip_validate_kop_fifo_override[2], \cceip_validate_kop_fifo_override.r.part0 [2]);
tran (cceip_validate_kop_fifo_override[2], \cceip_validate_kop_fifo_override.f.keyfilter_cmd_fifo );
tran (cceip_validate_kop_fifo_override[1], \cceip_validate_kop_fifo_override.r.part0 [1]);
tran (cceip_validate_kop_fifo_override[1], \cceip_validate_kop_fifo_override.f.gcm_tag_data_fifo );
tran (cceip_validate_kop_fifo_override[0], \cceip_validate_kop_fifo_override.r.part0 [0]);
tran (cceip_validate_kop_fifo_override[0], \cceip_validate_kop_fifo_override.f.gcm_cmd_fifo );
tran (cddip_decrypt_kop_fifo_override[6], \cddip_decrypt_kop_fifo_override.r.part0 [6]);
tran (cddip_decrypt_kop_fifo_override[6], \cddip_decrypt_kop_fifo_override.f.gcm_status_data_fifo );
tran (cddip_decrypt_kop_fifo_override[5], \cddip_decrypt_kop_fifo_override.r.part0 [5]);
tran (cddip_decrypt_kop_fifo_override[5], \cddip_decrypt_kop_fifo_override.f.tlv_sb_data_fifo );
tran (cddip_decrypt_kop_fifo_override[4], \cddip_decrypt_kop_fifo_override.r.part0 [4]);
tran (cddip_decrypt_kop_fifo_override[4], \cddip_decrypt_kop_fifo_override.f.kdf_cmd_fifo );
tran (cddip_decrypt_kop_fifo_override[3], \cddip_decrypt_kop_fifo_override.r.part0 [3]);
tran (cddip_decrypt_kop_fifo_override[3], \cddip_decrypt_kop_fifo_override.f.kdfstream_cmd_fifo );
tran (cddip_decrypt_kop_fifo_override[2], \cddip_decrypt_kop_fifo_override.r.part0 [2]);
tran (cddip_decrypt_kop_fifo_override[2], \cddip_decrypt_kop_fifo_override.f.keyfilter_cmd_fifo );
tran (cddip_decrypt_kop_fifo_override[1], \cddip_decrypt_kop_fifo_override.r.part0 [1]);
tran (cddip_decrypt_kop_fifo_override[1], \cddip_decrypt_kop_fifo_override.f.gcm_tag_data_fifo );
tran (cddip_decrypt_kop_fifo_override[0], \cddip_decrypt_kop_fifo_override.r.part0 [0]);
tran (cddip_decrypt_kop_fifo_override[0], \cddip_decrypt_kop_fifo_override.f.gcm_cmd_fifo );
tran (sa_global_ctrl[31], \sa_global_ctrl.r.part0 [31]);
tran (sa_global_ctrl[31], \sa_global_ctrl.f.spare [29]);
tran (sa_global_ctrl[30], \sa_global_ctrl.r.part0 [30]);
tran (sa_global_ctrl[30], \sa_global_ctrl.f.spare [28]);
tran (sa_global_ctrl[29], \sa_global_ctrl.r.part0 [29]);
tran (sa_global_ctrl[29], \sa_global_ctrl.f.spare [27]);
tran (sa_global_ctrl[28], \sa_global_ctrl.r.part0 [28]);
tran (sa_global_ctrl[28], \sa_global_ctrl.f.spare [26]);
tran (sa_global_ctrl[27], \sa_global_ctrl.r.part0 [27]);
tran (sa_global_ctrl[27], \sa_global_ctrl.f.spare [25]);
tran (sa_global_ctrl[26], \sa_global_ctrl.r.part0 [26]);
tran (sa_global_ctrl[26], \sa_global_ctrl.f.spare [24]);
tran (sa_global_ctrl[25], \sa_global_ctrl.r.part0 [25]);
tran (sa_global_ctrl[25], \sa_global_ctrl.f.spare [23]);
tran (sa_global_ctrl[24], \sa_global_ctrl.r.part0 [24]);
tran (sa_global_ctrl[24], \sa_global_ctrl.f.spare [22]);
tran (sa_global_ctrl[23], \sa_global_ctrl.r.part0 [23]);
tran (sa_global_ctrl[23], \sa_global_ctrl.f.spare [21]);
tran (sa_global_ctrl[22], \sa_global_ctrl.r.part0 [22]);
tran (sa_global_ctrl[22], \sa_global_ctrl.f.spare [20]);
tran (sa_global_ctrl[21], \sa_global_ctrl.r.part0 [21]);
tran (sa_global_ctrl[21], \sa_global_ctrl.f.spare [19]);
tran (sa_global_ctrl[20], \sa_global_ctrl.r.part0 [20]);
tran (sa_global_ctrl[20], \sa_global_ctrl.f.spare [18]);
tran (sa_global_ctrl[19], \sa_global_ctrl.r.part0 [19]);
tran (sa_global_ctrl[19], \sa_global_ctrl.f.spare [17]);
tran (sa_global_ctrl[18], \sa_global_ctrl.r.part0 [18]);
tran (sa_global_ctrl[18], \sa_global_ctrl.f.spare [16]);
tran (sa_global_ctrl[17], \sa_global_ctrl.r.part0 [17]);
tran (sa_global_ctrl[17], \sa_global_ctrl.f.spare [15]);
tran (sa_global_ctrl[16], \sa_global_ctrl.r.part0 [16]);
tran (sa_global_ctrl[16], \sa_global_ctrl.f.spare [14]);
tran (sa_global_ctrl[15], \sa_global_ctrl.r.part0 [15]);
tran (sa_global_ctrl[15], \sa_global_ctrl.f.spare [13]);
tran (sa_global_ctrl[14], \sa_global_ctrl.r.part0 [14]);
tran (sa_global_ctrl[14], \sa_global_ctrl.f.spare [12]);
tran (sa_global_ctrl[13], \sa_global_ctrl.r.part0 [13]);
tran (sa_global_ctrl[13], \sa_global_ctrl.f.spare [11]);
tran (sa_global_ctrl[12], \sa_global_ctrl.r.part0 [12]);
tran (sa_global_ctrl[12], \sa_global_ctrl.f.spare [10]);
tran (sa_global_ctrl[11], \sa_global_ctrl.r.part0 [11]);
tran (sa_global_ctrl[11], \sa_global_ctrl.f.spare [9]);
tran (sa_global_ctrl[10], \sa_global_ctrl.r.part0 [10]);
tran (sa_global_ctrl[10], \sa_global_ctrl.f.spare [8]);
tran (sa_global_ctrl[9], \sa_global_ctrl.r.part0 [9]);
tran (sa_global_ctrl[9], \sa_global_ctrl.f.spare [7]);
tran (sa_global_ctrl[8], \sa_global_ctrl.r.part0 [8]);
tran (sa_global_ctrl[8], \sa_global_ctrl.f.spare [6]);
tran (sa_global_ctrl[7], \sa_global_ctrl.r.part0 [7]);
tran (sa_global_ctrl[7], \sa_global_ctrl.f.spare [5]);
tran (sa_global_ctrl[6], \sa_global_ctrl.r.part0 [6]);
tran (sa_global_ctrl[6], \sa_global_ctrl.f.spare [4]);
tran (sa_global_ctrl[5], \sa_global_ctrl.r.part0 [5]);
tran (sa_global_ctrl[5], \sa_global_ctrl.f.spare [3]);
tran (sa_global_ctrl[4], \sa_global_ctrl.r.part0 [4]);
tran (sa_global_ctrl[4], \sa_global_ctrl.f.spare [2]);
tran (sa_global_ctrl[3], \sa_global_ctrl.r.part0 [3]);
tran (sa_global_ctrl[3], \sa_global_ctrl.f.spare [1]);
tran (sa_global_ctrl[2], \sa_global_ctrl.r.part0 [2]);
tran (sa_global_ctrl[2], \sa_global_ctrl.f.spare [0]);
tran (sa_global_ctrl[1], \sa_global_ctrl.r.part0 [1]);
tran (sa_global_ctrl[1], \sa_global_ctrl.f.sa_snap );
tran (sa_global_ctrl[0], \sa_global_ctrl.r.part0 [0]);
tran (sa_global_ctrl[0], \sa_global_ctrl.f.sa_clear_live );
tran (\sa_ctrl[0][0] , \sa_ctrl[0].r.part0[0] );
tran (\sa_ctrl[0][0] , \sa_ctrl[0].f.sa_event_sel[0] );
tran (\sa_ctrl[0][1] , \sa_ctrl[0].r.part0[1] );
tran (\sa_ctrl[0][1] , \sa_ctrl[0].f.sa_event_sel[1] );
tran (\sa_ctrl[0][2] , \sa_ctrl[0].r.part0[2] );
tran (\sa_ctrl[0][2] , \sa_ctrl[0].f.sa_event_sel[2] );
tran (\sa_ctrl[0][3] , \sa_ctrl[0].r.part0[3] );
tran (\sa_ctrl[0][3] , \sa_ctrl[0].f.sa_event_sel[3] );
tran (\sa_ctrl[0][4] , \sa_ctrl[0].r.part0[4] );
tran (\sa_ctrl[0][4] , \sa_ctrl[0].f.sa_event_sel[4] );
tran (\sa_ctrl[0][5] , \sa_ctrl[0].r.part0[5] );
tran (\sa_ctrl[0][5] , \sa_ctrl[0].f.spare[0] );
tran (\sa_ctrl[0][6] , \sa_ctrl[0].r.part0[6] );
tran (\sa_ctrl[0][6] , \sa_ctrl[0].f.spare[1] );
tran (\sa_ctrl[0][7] , \sa_ctrl[0].r.part0[7] );
tran (\sa_ctrl[0][7] , \sa_ctrl[0].f.spare[2] );
tran (\sa_ctrl[0][8] , \sa_ctrl[0].r.part0[8] );
tran (\sa_ctrl[0][8] , \sa_ctrl[0].f.spare[3] );
tran (\sa_ctrl[0][9] , \sa_ctrl[0].r.part0[9] );
tran (\sa_ctrl[0][9] , \sa_ctrl[0].f.spare[4] );
tran (\sa_ctrl[0][10] , \sa_ctrl[0].r.part0[10] );
tran (\sa_ctrl[0][10] , \sa_ctrl[0].f.spare[5] );
tran (\sa_ctrl[0][11] , \sa_ctrl[0].r.part0[11] );
tran (\sa_ctrl[0][11] , \sa_ctrl[0].f.spare[6] );
tran (\sa_ctrl[0][12] , \sa_ctrl[0].r.part0[12] );
tran (\sa_ctrl[0][12] , \sa_ctrl[0].f.spare[7] );
tran (\sa_ctrl[0][13] , \sa_ctrl[0].r.part0[13] );
tran (\sa_ctrl[0][13] , \sa_ctrl[0].f.spare[8] );
tran (\sa_ctrl[0][14] , \sa_ctrl[0].r.part0[14] );
tran (\sa_ctrl[0][14] , \sa_ctrl[0].f.spare[9] );
tran (\sa_ctrl[0][15] , \sa_ctrl[0].r.part0[15] );
tran (\sa_ctrl[0][15] , \sa_ctrl[0].f.spare[10] );
tran (\sa_ctrl[0][16] , \sa_ctrl[0].r.part0[16] );
tran (\sa_ctrl[0][16] , \sa_ctrl[0].f.spare[11] );
tran (\sa_ctrl[0][17] , \sa_ctrl[0].r.part0[17] );
tran (\sa_ctrl[0][17] , \sa_ctrl[0].f.spare[12] );
tran (\sa_ctrl[0][18] , \sa_ctrl[0].r.part0[18] );
tran (\sa_ctrl[0][18] , \sa_ctrl[0].f.spare[13] );
tran (\sa_ctrl[0][19] , \sa_ctrl[0].r.part0[19] );
tran (\sa_ctrl[0][19] , \sa_ctrl[0].f.spare[14] );
tran (\sa_ctrl[0][20] , \sa_ctrl[0].r.part0[20] );
tran (\sa_ctrl[0][20] , \sa_ctrl[0].f.spare[15] );
tran (\sa_ctrl[0][21] , \sa_ctrl[0].r.part0[21] );
tran (\sa_ctrl[0][21] , \sa_ctrl[0].f.spare[16] );
tran (\sa_ctrl[0][22] , \sa_ctrl[0].r.part0[22] );
tran (\sa_ctrl[0][22] , \sa_ctrl[0].f.spare[17] );
tran (\sa_ctrl[0][23] , \sa_ctrl[0].r.part0[23] );
tran (\sa_ctrl[0][23] , \sa_ctrl[0].f.spare[18] );
tran (\sa_ctrl[0][24] , \sa_ctrl[0].r.part0[24] );
tran (\sa_ctrl[0][24] , \sa_ctrl[0].f.spare[19] );
tran (\sa_ctrl[0][25] , \sa_ctrl[0].r.part0[25] );
tran (\sa_ctrl[0][25] , \sa_ctrl[0].f.spare[20] );
tran (\sa_ctrl[0][26] , \sa_ctrl[0].r.part0[26] );
tran (\sa_ctrl[0][26] , \sa_ctrl[0].f.spare[21] );
tran (\sa_ctrl[0][27] , \sa_ctrl[0].r.part0[27] );
tran (\sa_ctrl[0][27] , \sa_ctrl[0].f.spare[22] );
tran (\sa_ctrl[0][28] , \sa_ctrl[0].r.part0[28] );
tran (\sa_ctrl[0][28] , \sa_ctrl[0].f.spare[23] );
tran (\sa_ctrl[0][29] , \sa_ctrl[0].r.part0[29] );
tran (\sa_ctrl[0][29] , \sa_ctrl[0].f.spare[24] );
tran (\sa_ctrl[0][30] , \sa_ctrl[0].r.part0[30] );
tran (\sa_ctrl[0][30] , \sa_ctrl[0].f.spare[25] );
tran (\sa_ctrl[0][31] , \sa_ctrl[0].r.part0[31] );
tran (\sa_ctrl[0][31] , \sa_ctrl[0].f.spare[26] );
tran (\sa_ctrl[1][0] , \sa_ctrl[1].r.part0[0] );
tran (\sa_ctrl[1][0] , \sa_ctrl[1].f.sa_event_sel[0] );
tran (\sa_ctrl[1][1] , \sa_ctrl[1].r.part0[1] );
tran (\sa_ctrl[1][1] , \sa_ctrl[1].f.sa_event_sel[1] );
tran (\sa_ctrl[1][2] , \sa_ctrl[1].r.part0[2] );
tran (\sa_ctrl[1][2] , \sa_ctrl[1].f.sa_event_sel[2] );
tran (\sa_ctrl[1][3] , \sa_ctrl[1].r.part0[3] );
tran (\sa_ctrl[1][3] , \sa_ctrl[1].f.sa_event_sel[3] );
tran (\sa_ctrl[1][4] , \sa_ctrl[1].r.part0[4] );
tran (\sa_ctrl[1][4] , \sa_ctrl[1].f.sa_event_sel[4] );
tran (\sa_ctrl[1][5] , \sa_ctrl[1].r.part0[5] );
tran (\sa_ctrl[1][5] , \sa_ctrl[1].f.spare[0] );
tran (\sa_ctrl[1][6] , \sa_ctrl[1].r.part0[6] );
tran (\sa_ctrl[1][6] , \sa_ctrl[1].f.spare[1] );
tran (\sa_ctrl[1][7] , \sa_ctrl[1].r.part0[7] );
tran (\sa_ctrl[1][7] , \sa_ctrl[1].f.spare[2] );
tran (\sa_ctrl[1][8] , \sa_ctrl[1].r.part0[8] );
tran (\sa_ctrl[1][8] , \sa_ctrl[1].f.spare[3] );
tran (\sa_ctrl[1][9] , \sa_ctrl[1].r.part0[9] );
tran (\sa_ctrl[1][9] , \sa_ctrl[1].f.spare[4] );
tran (\sa_ctrl[1][10] , \sa_ctrl[1].r.part0[10] );
tran (\sa_ctrl[1][10] , \sa_ctrl[1].f.spare[5] );
tran (\sa_ctrl[1][11] , \sa_ctrl[1].r.part0[11] );
tran (\sa_ctrl[1][11] , \sa_ctrl[1].f.spare[6] );
tran (\sa_ctrl[1][12] , \sa_ctrl[1].r.part0[12] );
tran (\sa_ctrl[1][12] , \sa_ctrl[1].f.spare[7] );
tran (\sa_ctrl[1][13] , \sa_ctrl[1].r.part0[13] );
tran (\sa_ctrl[1][13] , \sa_ctrl[1].f.spare[8] );
tran (\sa_ctrl[1][14] , \sa_ctrl[1].r.part0[14] );
tran (\sa_ctrl[1][14] , \sa_ctrl[1].f.spare[9] );
tran (\sa_ctrl[1][15] , \sa_ctrl[1].r.part0[15] );
tran (\sa_ctrl[1][15] , \sa_ctrl[1].f.spare[10] );
tran (\sa_ctrl[1][16] , \sa_ctrl[1].r.part0[16] );
tran (\sa_ctrl[1][16] , \sa_ctrl[1].f.spare[11] );
tran (\sa_ctrl[1][17] , \sa_ctrl[1].r.part0[17] );
tran (\sa_ctrl[1][17] , \sa_ctrl[1].f.spare[12] );
tran (\sa_ctrl[1][18] , \sa_ctrl[1].r.part0[18] );
tran (\sa_ctrl[1][18] , \sa_ctrl[1].f.spare[13] );
tran (\sa_ctrl[1][19] , \sa_ctrl[1].r.part0[19] );
tran (\sa_ctrl[1][19] , \sa_ctrl[1].f.spare[14] );
tran (\sa_ctrl[1][20] , \sa_ctrl[1].r.part0[20] );
tran (\sa_ctrl[1][20] , \sa_ctrl[1].f.spare[15] );
tran (\sa_ctrl[1][21] , \sa_ctrl[1].r.part0[21] );
tran (\sa_ctrl[1][21] , \sa_ctrl[1].f.spare[16] );
tran (\sa_ctrl[1][22] , \sa_ctrl[1].r.part0[22] );
tran (\sa_ctrl[1][22] , \sa_ctrl[1].f.spare[17] );
tran (\sa_ctrl[1][23] , \sa_ctrl[1].r.part0[23] );
tran (\sa_ctrl[1][23] , \sa_ctrl[1].f.spare[18] );
tran (\sa_ctrl[1][24] , \sa_ctrl[1].r.part0[24] );
tran (\sa_ctrl[1][24] , \sa_ctrl[1].f.spare[19] );
tran (\sa_ctrl[1][25] , \sa_ctrl[1].r.part0[25] );
tran (\sa_ctrl[1][25] , \sa_ctrl[1].f.spare[20] );
tran (\sa_ctrl[1][26] , \sa_ctrl[1].r.part0[26] );
tran (\sa_ctrl[1][26] , \sa_ctrl[1].f.spare[21] );
tran (\sa_ctrl[1][27] , \sa_ctrl[1].r.part0[27] );
tran (\sa_ctrl[1][27] , \sa_ctrl[1].f.spare[22] );
tran (\sa_ctrl[1][28] , \sa_ctrl[1].r.part0[28] );
tran (\sa_ctrl[1][28] , \sa_ctrl[1].f.spare[23] );
tran (\sa_ctrl[1][29] , \sa_ctrl[1].r.part0[29] );
tran (\sa_ctrl[1][29] , \sa_ctrl[1].f.spare[24] );
tran (\sa_ctrl[1][30] , \sa_ctrl[1].r.part0[30] );
tran (\sa_ctrl[1][30] , \sa_ctrl[1].f.spare[25] );
tran (\sa_ctrl[1][31] , \sa_ctrl[1].r.part0[31] );
tran (\sa_ctrl[1][31] , \sa_ctrl[1].f.spare[26] );
tran (\sa_ctrl[2][0] , \sa_ctrl[2].r.part0[0] );
tran (\sa_ctrl[2][0] , \sa_ctrl[2].f.sa_event_sel[0] );
tran (\sa_ctrl[2][1] , \sa_ctrl[2].r.part0[1] );
tran (\sa_ctrl[2][1] , \sa_ctrl[2].f.sa_event_sel[1] );
tran (\sa_ctrl[2][2] , \sa_ctrl[2].r.part0[2] );
tran (\sa_ctrl[2][2] , \sa_ctrl[2].f.sa_event_sel[2] );
tran (\sa_ctrl[2][3] , \sa_ctrl[2].r.part0[3] );
tran (\sa_ctrl[2][3] , \sa_ctrl[2].f.sa_event_sel[3] );
tran (\sa_ctrl[2][4] , \sa_ctrl[2].r.part0[4] );
tran (\sa_ctrl[2][4] , \sa_ctrl[2].f.sa_event_sel[4] );
tran (\sa_ctrl[2][5] , \sa_ctrl[2].r.part0[5] );
tran (\sa_ctrl[2][5] , \sa_ctrl[2].f.spare[0] );
tran (\sa_ctrl[2][6] , \sa_ctrl[2].r.part0[6] );
tran (\sa_ctrl[2][6] , \sa_ctrl[2].f.spare[1] );
tran (\sa_ctrl[2][7] , \sa_ctrl[2].r.part0[7] );
tran (\sa_ctrl[2][7] , \sa_ctrl[2].f.spare[2] );
tran (\sa_ctrl[2][8] , \sa_ctrl[2].r.part0[8] );
tran (\sa_ctrl[2][8] , \sa_ctrl[2].f.spare[3] );
tran (\sa_ctrl[2][9] , \sa_ctrl[2].r.part0[9] );
tran (\sa_ctrl[2][9] , \sa_ctrl[2].f.spare[4] );
tran (\sa_ctrl[2][10] , \sa_ctrl[2].r.part0[10] );
tran (\sa_ctrl[2][10] , \sa_ctrl[2].f.spare[5] );
tran (\sa_ctrl[2][11] , \sa_ctrl[2].r.part0[11] );
tran (\sa_ctrl[2][11] , \sa_ctrl[2].f.spare[6] );
tran (\sa_ctrl[2][12] , \sa_ctrl[2].r.part0[12] );
tran (\sa_ctrl[2][12] , \sa_ctrl[2].f.spare[7] );
tran (\sa_ctrl[2][13] , \sa_ctrl[2].r.part0[13] );
tran (\sa_ctrl[2][13] , \sa_ctrl[2].f.spare[8] );
tran (\sa_ctrl[2][14] , \sa_ctrl[2].r.part0[14] );
tran (\sa_ctrl[2][14] , \sa_ctrl[2].f.spare[9] );
tran (\sa_ctrl[2][15] , \sa_ctrl[2].r.part0[15] );
tran (\sa_ctrl[2][15] , \sa_ctrl[2].f.spare[10] );
tran (\sa_ctrl[2][16] , \sa_ctrl[2].r.part0[16] );
tran (\sa_ctrl[2][16] , \sa_ctrl[2].f.spare[11] );
tran (\sa_ctrl[2][17] , \sa_ctrl[2].r.part0[17] );
tran (\sa_ctrl[2][17] , \sa_ctrl[2].f.spare[12] );
tran (\sa_ctrl[2][18] , \sa_ctrl[2].r.part0[18] );
tran (\sa_ctrl[2][18] , \sa_ctrl[2].f.spare[13] );
tran (\sa_ctrl[2][19] , \sa_ctrl[2].r.part0[19] );
tran (\sa_ctrl[2][19] , \sa_ctrl[2].f.spare[14] );
tran (\sa_ctrl[2][20] , \sa_ctrl[2].r.part0[20] );
tran (\sa_ctrl[2][20] , \sa_ctrl[2].f.spare[15] );
tran (\sa_ctrl[2][21] , \sa_ctrl[2].r.part0[21] );
tran (\sa_ctrl[2][21] , \sa_ctrl[2].f.spare[16] );
tran (\sa_ctrl[2][22] , \sa_ctrl[2].r.part0[22] );
tran (\sa_ctrl[2][22] , \sa_ctrl[2].f.spare[17] );
tran (\sa_ctrl[2][23] , \sa_ctrl[2].r.part0[23] );
tran (\sa_ctrl[2][23] , \sa_ctrl[2].f.spare[18] );
tran (\sa_ctrl[2][24] , \sa_ctrl[2].r.part0[24] );
tran (\sa_ctrl[2][24] , \sa_ctrl[2].f.spare[19] );
tran (\sa_ctrl[2][25] , \sa_ctrl[2].r.part0[25] );
tran (\sa_ctrl[2][25] , \sa_ctrl[2].f.spare[20] );
tran (\sa_ctrl[2][26] , \sa_ctrl[2].r.part0[26] );
tran (\sa_ctrl[2][26] , \sa_ctrl[2].f.spare[21] );
tran (\sa_ctrl[2][27] , \sa_ctrl[2].r.part0[27] );
tran (\sa_ctrl[2][27] , \sa_ctrl[2].f.spare[22] );
tran (\sa_ctrl[2][28] , \sa_ctrl[2].r.part0[28] );
tran (\sa_ctrl[2][28] , \sa_ctrl[2].f.spare[23] );
tran (\sa_ctrl[2][29] , \sa_ctrl[2].r.part0[29] );
tran (\sa_ctrl[2][29] , \sa_ctrl[2].f.spare[24] );
tran (\sa_ctrl[2][30] , \sa_ctrl[2].r.part0[30] );
tran (\sa_ctrl[2][30] , \sa_ctrl[2].f.spare[25] );
tran (\sa_ctrl[2][31] , \sa_ctrl[2].r.part0[31] );
tran (\sa_ctrl[2][31] , \sa_ctrl[2].f.spare[26] );
tran (\sa_ctrl[3][0] , \sa_ctrl[3].r.part0[0] );
tran (\sa_ctrl[3][0] , \sa_ctrl[3].f.sa_event_sel[0] );
tran (\sa_ctrl[3][1] , \sa_ctrl[3].r.part0[1] );
tran (\sa_ctrl[3][1] , \sa_ctrl[3].f.sa_event_sel[1] );
tran (\sa_ctrl[3][2] , \sa_ctrl[3].r.part0[2] );
tran (\sa_ctrl[3][2] , \sa_ctrl[3].f.sa_event_sel[2] );
tran (\sa_ctrl[3][3] , \sa_ctrl[3].r.part0[3] );
tran (\sa_ctrl[3][3] , \sa_ctrl[3].f.sa_event_sel[3] );
tran (\sa_ctrl[3][4] , \sa_ctrl[3].r.part0[4] );
tran (\sa_ctrl[3][4] , \sa_ctrl[3].f.sa_event_sel[4] );
tran (\sa_ctrl[3][5] , \sa_ctrl[3].r.part0[5] );
tran (\sa_ctrl[3][5] , \sa_ctrl[3].f.spare[0] );
tran (\sa_ctrl[3][6] , \sa_ctrl[3].r.part0[6] );
tran (\sa_ctrl[3][6] , \sa_ctrl[3].f.spare[1] );
tran (\sa_ctrl[3][7] , \sa_ctrl[3].r.part0[7] );
tran (\sa_ctrl[3][7] , \sa_ctrl[3].f.spare[2] );
tran (\sa_ctrl[3][8] , \sa_ctrl[3].r.part0[8] );
tran (\sa_ctrl[3][8] , \sa_ctrl[3].f.spare[3] );
tran (\sa_ctrl[3][9] , \sa_ctrl[3].r.part0[9] );
tran (\sa_ctrl[3][9] , \sa_ctrl[3].f.spare[4] );
tran (\sa_ctrl[3][10] , \sa_ctrl[3].r.part0[10] );
tran (\sa_ctrl[3][10] , \sa_ctrl[3].f.spare[5] );
tran (\sa_ctrl[3][11] , \sa_ctrl[3].r.part0[11] );
tran (\sa_ctrl[3][11] , \sa_ctrl[3].f.spare[6] );
tran (\sa_ctrl[3][12] , \sa_ctrl[3].r.part0[12] );
tran (\sa_ctrl[3][12] , \sa_ctrl[3].f.spare[7] );
tran (\sa_ctrl[3][13] , \sa_ctrl[3].r.part0[13] );
tran (\sa_ctrl[3][13] , \sa_ctrl[3].f.spare[8] );
tran (\sa_ctrl[3][14] , \sa_ctrl[3].r.part0[14] );
tran (\sa_ctrl[3][14] , \sa_ctrl[3].f.spare[9] );
tran (\sa_ctrl[3][15] , \sa_ctrl[3].r.part0[15] );
tran (\sa_ctrl[3][15] , \sa_ctrl[3].f.spare[10] );
tran (\sa_ctrl[3][16] , \sa_ctrl[3].r.part0[16] );
tran (\sa_ctrl[3][16] , \sa_ctrl[3].f.spare[11] );
tran (\sa_ctrl[3][17] , \sa_ctrl[3].r.part0[17] );
tran (\sa_ctrl[3][17] , \sa_ctrl[3].f.spare[12] );
tran (\sa_ctrl[3][18] , \sa_ctrl[3].r.part0[18] );
tran (\sa_ctrl[3][18] , \sa_ctrl[3].f.spare[13] );
tran (\sa_ctrl[3][19] , \sa_ctrl[3].r.part0[19] );
tran (\sa_ctrl[3][19] , \sa_ctrl[3].f.spare[14] );
tran (\sa_ctrl[3][20] , \sa_ctrl[3].r.part0[20] );
tran (\sa_ctrl[3][20] , \sa_ctrl[3].f.spare[15] );
tran (\sa_ctrl[3][21] , \sa_ctrl[3].r.part0[21] );
tran (\sa_ctrl[3][21] , \sa_ctrl[3].f.spare[16] );
tran (\sa_ctrl[3][22] , \sa_ctrl[3].r.part0[22] );
tran (\sa_ctrl[3][22] , \sa_ctrl[3].f.spare[17] );
tran (\sa_ctrl[3][23] , \sa_ctrl[3].r.part0[23] );
tran (\sa_ctrl[3][23] , \sa_ctrl[3].f.spare[18] );
tran (\sa_ctrl[3][24] , \sa_ctrl[3].r.part0[24] );
tran (\sa_ctrl[3][24] , \sa_ctrl[3].f.spare[19] );
tran (\sa_ctrl[3][25] , \sa_ctrl[3].r.part0[25] );
tran (\sa_ctrl[3][25] , \sa_ctrl[3].f.spare[20] );
tran (\sa_ctrl[3][26] , \sa_ctrl[3].r.part0[26] );
tran (\sa_ctrl[3][26] , \sa_ctrl[3].f.spare[21] );
tran (\sa_ctrl[3][27] , \sa_ctrl[3].r.part0[27] );
tran (\sa_ctrl[3][27] , \sa_ctrl[3].f.spare[22] );
tran (\sa_ctrl[3][28] , \sa_ctrl[3].r.part0[28] );
tran (\sa_ctrl[3][28] , \sa_ctrl[3].f.spare[23] );
tran (\sa_ctrl[3][29] , \sa_ctrl[3].r.part0[29] );
tran (\sa_ctrl[3][29] , \sa_ctrl[3].f.spare[24] );
tran (\sa_ctrl[3][30] , \sa_ctrl[3].r.part0[30] );
tran (\sa_ctrl[3][30] , \sa_ctrl[3].f.spare[25] );
tran (\sa_ctrl[3][31] , \sa_ctrl[3].r.part0[31] );
tran (\sa_ctrl[3][31] , \sa_ctrl[3].f.spare[26] );
tran (\sa_ctrl[4][0] , \sa_ctrl[4].r.part0[0] );
tran (\sa_ctrl[4][0] , \sa_ctrl[4].f.sa_event_sel[0] );
tran (\sa_ctrl[4][1] , \sa_ctrl[4].r.part0[1] );
tran (\sa_ctrl[4][1] , \sa_ctrl[4].f.sa_event_sel[1] );
tran (\sa_ctrl[4][2] , \sa_ctrl[4].r.part0[2] );
tran (\sa_ctrl[4][2] , \sa_ctrl[4].f.sa_event_sel[2] );
tran (\sa_ctrl[4][3] , \sa_ctrl[4].r.part0[3] );
tran (\sa_ctrl[4][3] , \sa_ctrl[4].f.sa_event_sel[3] );
tran (\sa_ctrl[4][4] , \sa_ctrl[4].r.part0[4] );
tran (\sa_ctrl[4][4] , \sa_ctrl[4].f.sa_event_sel[4] );
tran (\sa_ctrl[4][5] , \sa_ctrl[4].r.part0[5] );
tran (\sa_ctrl[4][5] , \sa_ctrl[4].f.spare[0] );
tran (\sa_ctrl[4][6] , \sa_ctrl[4].r.part0[6] );
tran (\sa_ctrl[4][6] , \sa_ctrl[4].f.spare[1] );
tran (\sa_ctrl[4][7] , \sa_ctrl[4].r.part0[7] );
tran (\sa_ctrl[4][7] , \sa_ctrl[4].f.spare[2] );
tran (\sa_ctrl[4][8] , \sa_ctrl[4].r.part0[8] );
tran (\sa_ctrl[4][8] , \sa_ctrl[4].f.spare[3] );
tran (\sa_ctrl[4][9] , \sa_ctrl[4].r.part0[9] );
tran (\sa_ctrl[4][9] , \sa_ctrl[4].f.spare[4] );
tran (\sa_ctrl[4][10] , \sa_ctrl[4].r.part0[10] );
tran (\sa_ctrl[4][10] , \sa_ctrl[4].f.spare[5] );
tran (\sa_ctrl[4][11] , \sa_ctrl[4].r.part0[11] );
tran (\sa_ctrl[4][11] , \sa_ctrl[4].f.spare[6] );
tran (\sa_ctrl[4][12] , \sa_ctrl[4].r.part0[12] );
tran (\sa_ctrl[4][12] , \sa_ctrl[4].f.spare[7] );
tran (\sa_ctrl[4][13] , \sa_ctrl[4].r.part0[13] );
tran (\sa_ctrl[4][13] , \sa_ctrl[4].f.spare[8] );
tran (\sa_ctrl[4][14] , \sa_ctrl[4].r.part0[14] );
tran (\sa_ctrl[4][14] , \sa_ctrl[4].f.spare[9] );
tran (\sa_ctrl[4][15] , \sa_ctrl[4].r.part0[15] );
tran (\sa_ctrl[4][15] , \sa_ctrl[4].f.spare[10] );
tran (\sa_ctrl[4][16] , \sa_ctrl[4].r.part0[16] );
tran (\sa_ctrl[4][16] , \sa_ctrl[4].f.spare[11] );
tran (\sa_ctrl[4][17] , \sa_ctrl[4].r.part0[17] );
tran (\sa_ctrl[4][17] , \sa_ctrl[4].f.spare[12] );
tran (\sa_ctrl[4][18] , \sa_ctrl[4].r.part0[18] );
tran (\sa_ctrl[4][18] , \sa_ctrl[4].f.spare[13] );
tran (\sa_ctrl[4][19] , \sa_ctrl[4].r.part0[19] );
tran (\sa_ctrl[4][19] , \sa_ctrl[4].f.spare[14] );
tran (\sa_ctrl[4][20] , \sa_ctrl[4].r.part0[20] );
tran (\sa_ctrl[4][20] , \sa_ctrl[4].f.spare[15] );
tran (\sa_ctrl[4][21] , \sa_ctrl[4].r.part0[21] );
tran (\sa_ctrl[4][21] , \sa_ctrl[4].f.spare[16] );
tran (\sa_ctrl[4][22] , \sa_ctrl[4].r.part0[22] );
tran (\sa_ctrl[4][22] , \sa_ctrl[4].f.spare[17] );
tran (\sa_ctrl[4][23] , \sa_ctrl[4].r.part0[23] );
tran (\sa_ctrl[4][23] , \sa_ctrl[4].f.spare[18] );
tran (\sa_ctrl[4][24] , \sa_ctrl[4].r.part0[24] );
tran (\sa_ctrl[4][24] , \sa_ctrl[4].f.spare[19] );
tran (\sa_ctrl[4][25] , \sa_ctrl[4].r.part0[25] );
tran (\sa_ctrl[4][25] , \sa_ctrl[4].f.spare[20] );
tran (\sa_ctrl[4][26] , \sa_ctrl[4].r.part0[26] );
tran (\sa_ctrl[4][26] , \sa_ctrl[4].f.spare[21] );
tran (\sa_ctrl[4][27] , \sa_ctrl[4].r.part0[27] );
tran (\sa_ctrl[4][27] , \sa_ctrl[4].f.spare[22] );
tran (\sa_ctrl[4][28] , \sa_ctrl[4].r.part0[28] );
tran (\sa_ctrl[4][28] , \sa_ctrl[4].f.spare[23] );
tran (\sa_ctrl[4][29] , \sa_ctrl[4].r.part0[29] );
tran (\sa_ctrl[4][29] , \sa_ctrl[4].f.spare[24] );
tran (\sa_ctrl[4][30] , \sa_ctrl[4].r.part0[30] );
tran (\sa_ctrl[4][30] , \sa_ctrl[4].f.spare[25] );
tran (\sa_ctrl[4][31] , \sa_ctrl[4].r.part0[31] );
tran (\sa_ctrl[4][31] , \sa_ctrl[4].f.spare[26] );
tran (\sa_ctrl[5][0] , \sa_ctrl[5].r.part0[0] );
tran (\sa_ctrl[5][0] , \sa_ctrl[5].f.sa_event_sel[0] );
tran (\sa_ctrl[5][1] , \sa_ctrl[5].r.part0[1] );
tran (\sa_ctrl[5][1] , \sa_ctrl[5].f.sa_event_sel[1] );
tran (\sa_ctrl[5][2] , \sa_ctrl[5].r.part0[2] );
tran (\sa_ctrl[5][2] , \sa_ctrl[5].f.sa_event_sel[2] );
tran (\sa_ctrl[5][3] , \sa_ctrl[5].r.part0[3] );
tran (\sa_ctrl[5][3] , \sa_ctrl[5].f.sa_event_sel[3] );
tran (\sa_ctrl[5][4] , \sa_ctrl[5].r.part0[4] );
tran (\sa_ctrl[5][4] , \sa_ctrl[5].f.sa_event_sel[4] );
tran (\sa_ctrl[5][5] , \sa_ctrl[5].r.part0[5] );
tran (\sa_ctrl[5][5] , \sa_ctrl[5].f.spare[0] );
tran (\sa_ctrl[5][6] , \sa_ctrl[5].r.part0[6] );
tran (\sa_ctrl[5][6] , \sa_ctrl[5].f.spare[1] );
tran (\sa_ctrl[5][7] , \sa_ctrl[5].r.part0[7] );
tran (\sa_ctrl[5][7] , \sa_ctrl[5].f.spare[2] );
tran (\sa_ctrl[5][8] , \sa_ctrl[5].r.part0[8] );
tran (\sa_ctrl[5][8] , \sa_ctrl[5].f.spare[3] );
tran (\sa_ctrl[5][9] , \sa_ctrl[5].r.part0[9] );
tran (\sa_ctrl[5][9] , \sa_ctrl[5].f.spare[4] );
tran (\sa_ctrl[5][10] , \sa_ctrl[5].r.part0[10] );
tran (\sa_ctrl[5][10] , \sa_ctrl[5].f.spare[5] );
tran (\sa_ctrl[5][11] , \sa_ctrl[5].r.part0[11] );
tran (\sa_ctrl[5][11] , \sa_ctrl[5].f.spare[6] );
tran (\sa_ctrl[5][12] , \sa_ctrl[5].r.part0[12] );
tran (\sa_ctrl[5][12] , \sa_ctrl[5].f.spare[7] );
tran (\sa_ctrl[5][13] , \sa_ctrl[5].r.part0[13] );
tran (\sa_ctrl[5][13] , \sa_ctrl[5].f.spare[8] );
tran (\sa_ctrl[5][14] , \sa_ctrl[5].r.part0[14] );
tran (\sa_ctrl[5][14] , \sa_ctrl[5].f.spare[9] );
tran (\sa_ctrl[5][15] , \sa_ctrl[5].r.part0[15] );
tran (\sa_ctrl[5][15] , \sa_ctrl[5].f.spare[10] );
tran (\sa_ctrl[5][16] , \sa_ctrl[5].r.part0[16] );
tran (\sa_ctrl[5][16] , \sa_ctrl[5].f.spare[11] );
tran (\sa_ctrl[5][17] , \sa_ctrl[5].r.part0[17] );
tran (\sa_ctrl[5][17] , \sa_ctrl[5].f.spare[12] );
tran (\sa_ctrl[5][18] , \sa_ctrl[5].r.part0[18] );
tran (\sa_ctrl[5][18] , \sa_ctrl[5].f.spare[13] );
tran (\sa_ctrl[5][19] , \sa_ctrl[5].r.part0[19] );
tran (\sa_ctrl[5][19] , \sa_ctrl[5].f.spare[14] );
tran (\sa_ctrl[5][20] , \sa_ctrl[5].r.part0[20] );
tran (\sa_ctrl[5][20] , \sa_ctrl[5].f.spare[15] );
tran (\sa_ctrl[5][21] , \sa_ctrl[5].r.part0[21] );
tran (\sa_ctrl[5][21] , \sa_ctrl[5].f.spare[16] );
tran (\sa_ctrl[5][22] , \sa_ctrl[5].r.part0[22] );
tran (\sa_ctrl[5][22] , \sa_ctrl[5].f.spare[17] );
tran (\sa_ctrl[5][23] , \sa_ctrl[5].r.part0[23] );
tran (\sa_ctrl[5][23] , \sa_ctrl[5].f.spare[18] );
tran (\sa_ctrl[5][24] , \sa_ctrl[5].r.part0[24] );
tran (\sa_ctrl[5][24] , \sa_ctrl[5].f.spare[19] );
tran (\sa_ctrl[5][25] , \sa_ctrl[5].r.part0[25] );
tran (\sa_ctrl[5][25] , \sa_ctrl[5].f.spare[20] );
tran (\sa_ctrl[5][26] , \sa_ctrl[5].r.part0[26] );
tran (\sa_ctrl[5][26] , \sa_ctrl[5].f.spare[21] );
tran (\sa_ctrl[5][27] , \sa_ctrl[5].r.part0[27] );
tran (\sa_ctrl[5][27] , \sa_ctrl[5].f.spare[22] );
tran (\sa_ctrl[5][28] , \sa_ctrl[5].r.part0[28] );
tran (\sa_ctrl[5][28] , \sa_ctrl[5].f.spare[23] );
tran (\sa_ctrl[5][29] , \sa_ctrl[5].r.part0[29] );
tran (\sa_ctrl[5][29] , \sa_ctrl[5].f.spare[24] );
tran (\sa_ctrl[5][30] , \sa_ctrl[5].r.part0[30] );
tran (\sa_ctrl[5][30] , \sa_ctrl[5].f.spare[25] );
tran (\sa_ctrl[5][31] , \sa_ctrl[5].r.part0[31] );
tran (\sa_ctrl[5][31] , \sa_ctrl[5].f.spare[26] );
tran (\sa_ctrl[6][0] , \sa_ctrl[6].r.part0[0] );
tran (\sa_ctrl[6][0] , \sa_ctrl[6].f.sa_event_sel[0] );
tran (\sa_ctrl[6][1] , \sa_ctrl[6].r.part0[1] );
tran (\sa_ctrl[6][1] , \sa_ctrl[6].f.sa_event_sel[1] );
tran (\sa_ctrl[6][2] , \sa_ctrl[6].r.part0[2] );
tran (\sa_ctrl[6][2] , \sa_ctrl[6].f.sa_event_sel[2] );
tran (\sa_ctrl[6][3] , \sa_ctrl[6].r.part0[3] );
tran (\sa_ctrl[6][3] , \sa_ctrl[6].f.sa_event_sel[3] );
tran (\sa_ctrl[6][4] , \sa_ctrl[6].r.part0[4] );
tran (\sa_ctrl[6][4] , \sa_ctrl[6].f.sa_event_sel[4] );
tran (\sa_ctrl[6][5] , \sa_ctrl[6].r.part0[5] );
tran (\sa_ctrl[6][5] , \sa_ctrl[6].f.spare[0] );
tran (\sa_ctrl[6][6] , \sa_ctrl[6].r.part0[6] );
tran (\sa_ctrl[6][6] , \sa_ctrl[6].f.spare[1] );
tran (\sa_ctrl[6][7] , \sa_ctrl[6].r.part0[7] );
tran (\sa_ctrl[6][7] , \sa_ctrl[6].f.spare[2] );
tran (\sa_ctrl[6][8] , \sa_ctrl[6].r.part0[8] );
tran (\sa_ctrl[6][8] , \sa_ctrl[6].f.spare[3] );
tran (\sa_ctrl[6][9] , \sa_ctrl[6].r.part0[9] );
tran (\sa_ctrl[6][9] , \sa_ctrl[6].f.spare[4] );
tran (\sa_ctrl[6][10] , \sa_ctrl[6].r.part0[10] );
tran (\sa_ctrl[6][10] , \sa_ctrl[6].f.spare[5] );
tran (\sa_ctrl[6][11] , \sa_ctrl[6].r.part0[11] );
tran (\sa_ctrl[6][11] , \sa_ctrl[6].f.spare[6] );
tran (\sa_ctrl[6][12] , \sa_ctrl[6].r.part0[12] );
tran (\sa_ctrl[6][12] , \sa_ctrl[6].f.spare[7] );
tran (\sa_ctrl[6][13] , \sa_ctrl[6].r.part0[13] );
tran (\sa_ctrl[6][13] , \sa_ctrl[6].f.spare[8] );
tran (\sa_ctrl[6][14] , \sa_ctrl[6].r.part0[14] );
tran (\sa_ctrl[6][14] , \sa_ctrl[6].f.spare[9] );
tran (\sa_ctrl[6][15] , \sa_ctrl[6].r.part0[15] );
tran (\sa_ctrl[6][15] , \sa_ctrl[6].f.spare[10] );
tran (\sa_ctrl[6][16] , \sa_ctrl[6].r.part0[16] );
tran (\sa_ctrl[6][16] , \sa_ctrl[6].f.spare[11] );
tran (\sa_ctrl[6][17] , \sa_ctrl[6].r.part0[17] );
tran (\sa_ctrl[6][17] , \sa_ctrl[6].f.spare[12] );
tran (\sa_ctrl[6][18] , \sa_ctrl[6].r.part0[18] );
tran (\sa_ctrl[6][18] , \sa_ctrl[6].f.spare[13] );
tran (\sa_ctrl[6][19] , \sa_ctrl[6].r.part0[19] );
tran (\sa_ctrl[6][19] , \sa_ctrl[6].f.spare[14] );
tran (\sa_ctrl[6][20] , \sa_ctrl[6].r.part0[20] );
tran (\sa_ctrl[6][20] , \sa_ctrl[6].f.spare[15] );
tran (\sa_ctrl[6][21] , \sa_ctrl[6].r.part0[21] );
tran (\sa_ctrl[6][21] , \sa_ctrl[6].f.spare[16] );
tran (\sa_ctrl[6][22] , \sa_ctrl[6].r.part0[22] );
tran (\sa_ctrl[6][22] , \sa_ctrl[6].f.spare[17] );
tran (\sa_ctrl[6][23] , \sa_ctrl[6].r.part0[23] );
tran (\sa_ctrl[6][23] , \sa_ctrl[6].f.spare[18] );
tran (\sa_ctrl[6][24] , \sa_ctrl[6].r.part0[24] );
tran (\sa_ctrl[6][24] , \sa_ctrl[6].f.spare[19] );
tran (\sa_ctrl[6][25] , \sa_ctrl[6].r.part0[25] );
tran (\sa_ctrl[6][25] , \sa_ctrl[6].f.spare[20] );
tran (\sa_ctrl[6][26] , \sa_ctrl[6].r.part0[26] );
tran (\sa_ctrl[6][26] , \sa_ctrl[6].f.spare[21] );
tran (\sa_ctrl[6][27] , \sa_ctrl[6].r.part0[27] );
tran (\sa_ctrl[6][27] , \sa_ctrl[6].f.spare[22] );
tran (\sa_ctrl[6][28] , \sa_ctrl[6].r.part0[28] );
tran (\sa_ctrl[6][28] , \sa_ctrl[6].f.spare[23] );
tran (\sa_ctrl[6][29] , \sa_ctrl[6].r.part0[29] );
tran (\sa_ctrl[6][29] , \sa_ctrl[6].f.spare[24] );
tran (\sa_ctrl[6][30] , \sa_ctrl[6].r.part0[30] );
tran (\sa_ctrl[6][30] , \sa_ctrl[6].f.spare[25] );
tran (\sa_ctrl[6][31] , \sa_ctrl[6].r.part0[31] );
tran (\sa_ctrl[6][31] , \sa_ctrl[6].f.spare[26] );
tran (\sa_ctrl[7][0] , \sa_ctrl[7].r.part0[0] );
tran (\sa_ctrl[7][0] , \sa_ctrl[7].f.sa_event_sel[0] );
tran (\sa_ctrl[7][1] , \sa_ctrl[7].r.part0[1] );
tran (\sa_ctrl[7][1] , \sa_ctrl[7].f.sa_event_sel[1] );
tran (\sa_ctrl[7][2] , \sa_ctrl[7].r.part0[2] );
tran (\sa_ctrl[7][2] , \sa_ctrl[7].f.sa_event_sel[2] );
tran (\sa_ctrl[7][3] , \sa_ctrl[7].r.part0[3] );
tran (\sa_ctrl[7][3] , \sa_ctrl[7].f.sa_event_sel[3] );
tran (\sa_ctrl[7][4] , \sa_ctrl[7].r.part0[4] );
tran (\sa_ctrl[7][4] , \sa_ctrl[7].f.sa_event_sel[4] );
tran (\sa_ctrl[7][5] , \sa_ctrl[7].r.part0[5] );
tran (\sa_ctrl[7][5] , \sa_ctrl[7].f.spare[0] );
tran (\sa_ctrl[7][6] , \sa_ctrl[7].r.part0[6] );
tran (\sa_ctrl[7][6] , \sa_ctrl[7].f.spare[1] );
tran (\sa_ctrl[7][7] , \sa_ctrl[7].r.part0[7] );
tran (\sa_ctrl[7][7] , \sa_ctrl[7].f.spare[2] );
tran (\sa_ctrl[7][8] , \sa_ctrl[7].r.part0[8] );
tran (\sa_ctrl[7][8] , \sa_ctrl[7].f.spare[3] );
tran (\sa_ctrl[7][9] , \sa_ctrl[7].r.part0[9] );
tran (\sa_ctrl[7][9] , \sa_ctrl[7].f.spare[4] );
tran (\sa_ctrl[7][10] , \sa_ctrl[7].r.part0[10] );
tran (\sa_ctrl[7][10] , \sa_ctrl[7].f.spare[5] );
tran (\sa_ctrl[7][11] , \sa_ctrl[7].r.part0[11] );
tran (\sa_ctrl[7][11] , \sa_ctrl[7].f.spare[6] );
tran (\sa_ctrl[7][12] , \sa_ctrl[7].r.part0[12] );
tran (\sa_ctrl[7][12] , \sa_ctrl[7].f.spare[7] );
tran (\sa_ctrl[7][13] , \sa_ctrl[7].r.part0[13] );
tran (\sa_ctrl[7][13] , \sa_ctrl[7].f.spare[8] );
tran (\sa_ctrl[7][14] , \sa_ctrl[7].r.part0[14] );
tran (\sa_ctrl[7][14] , \sa_ctrl[7].f.spare[9] );
tran (\sa_ctrl[7][15] , \sa_ctrl[7].r.part0[15] );
tran (\sa_ctrl[7][15] , \sa_ctrl[7].f.spare[10] );
tran (\sa_ctrl[7][16] , \sa_ctrl[7].r.part0[16] );
tran (\sa_ctrl[7][16] , \sa_ctrl[7].f.spare[11] );
tran (\sa_ctrl[7][17] , \sa_ctrl[7].r.part0[17] );
tran (\sa_ctrl[7][17] , \sa_ctrl[7].f.spare[12] );
tran (\sa_ctrl[7][18] , \sa_ctrl[7].r.part0[18] );
tran (\sa_ctrl[7][18] , \sa_ctrl[7].f.spare[13] );
tran (\sa_ctrl[7][19] , \sa_ctrl[7].r.part0[19] );
tran (\sa_ctrl[7][19] , \sa_ctrl[7].f.spare[14] );
tran (\sa_ctrl[7][20] , \sa_ctrl[7].r.part0[20] );
tran (\sa_ctrl[7][20] , \sa_ctrl[7].f.spare[15] );
tran (\sa_ctrl[7][21] , \sa_ctrl[7].r.part0[21] );
tran (\sa_ctrl[7][21] , \sa_ctrl[7].f.spare[16] );
tran (\sa_ctrl[7][22] , \sa_ctrl[7].r.part0[22] );
tran (\sa_ctrl[7][22] , \sa_ctrl[7].f.spare[17] );
tran (\sa_ctrl[7][23] , \sa_ctrl[7].r.part0[23] );
tran (\sa_ctrl[7][23] , \sa_ctrl[7].f.spare[18] );
tran (\sa_ctrl[7][24] , \sa_ctrl[7].r.part0[24] );
tran (\sa_ctrl[7][24] , \sa_ctrl[7].f.spare[19] );
tran (\sa_ctrl[7][25] , \sa_ctrl[7].r.part0[25] );
tran (\sa_ctrl[7][25] , \sa_ctrl[7].f.spare[20] );
tran (\sa_ctrl[7][26] , \sa_ctrl[7].r.part0[26] );
tran (\sa_ctrl[7][26] , \sa_ctrl[7].f.spare[21] );
tran (\sa_ctrl[7][27] , \sa_ctrl[7].r.part0[27] );
tran (\sa_ctrl[7][27] , \sa_ctrl[7].f.spare[22] );
tran (\sa_ctrl[7][28] , \sa_ctrl[7].r.part0[28] );
tran (\sa_ctrl[7][28] , \sa_ctrl[7].f.spare[23] );
tran (\sa_ctrl[7][29] , \sa_ctrl[7].r.part0[29] );
tran (\sa_ctrl[7][29] , \sa_ctrl[7].f.spare[24] );
tran (\sa_ctrl[7][30] , \sa_ctrl[7].r.part0[30] );
tran (\sa_ctrl[7][30] , \sa_ctrl[7].f.spare[25] );
tran (\sa_ctrl[7][31] , \sa_ctrl[7].r.part0[31] );
tran (\sa_ctrl[7][31] , \sa_ctrl[7].f.spare[26] );
tran (\sa_ctrl[8][0] , \sa_ctrl[8].r.part0[0] );
tran (\sa_ctrl[8][0] , \sa_ctrl[8].f.sa_event_sel[0] );
tran (\sa_ctrl[8][1] , \sa_ctrl[8].r.part0[1] );
tran (\sa_ctrl[8][1] , \sa_ctrl[8].f.sa_event_sel[1] );
tran (\sa_ctrl[8][2] , \sa_ctrl[8].r.part0[2] );
tran (\sa_ctrl[8][2] , \sa_ctrl[8].f.sa_event_sel[2] );
tran (\sa_ctrl[8][3] , \sa_ctrl[8].r.part0[3] );
tran (\sa_ctrl[8][3] , \sa_ctrl[8].f.sa_event_sel[3] );
tran (\sa_ctrl[8][4] , \sa_ctrl[8].r.part0[4] );
tran (\sa_ctrl[8][4] , \sa_ctrl[8].f.sa_event_sel[4] );
tran (\sa_ctrl[8][5] , \sa_ctrl[8].r.part0[5] );
tran (\sa_ctrl[8][5] , \sa_ctrl[8].f.spare[0] );
tran (\sa_ctrl[8][6] , \sa_ctrl[8].r.part0[6] );
tran (\sa_ctrl[8][6] , \sa_ctrl[8].f.spare[1] );
tran (\sa_ctrl[8][7] , \sa_ctrl[8].r.part0[7] );
tran (\sa_ctrl[8][7] , \sa_ctrl[8].f.spare[2] );
tran (\sa_ctrl[8][8] , \sa_ctrl[8].r.part0[8] );
tran (\sa_ctrl[8][8] , \sa_ctrl[8].f.spare[3] );
tran (\sa_ctrl[8][9] , \sa_ctrl[8].r.part0[9] );
tran (\sa_ctrl[8][9] , \sa_ctrl[8].f.spare[4] );
tran (\sa_ctrl[8][10] , \sa_ctrl[8].r.part0[10] );
tran (\sa_ctrl[8][10] , \sa_ctrl[8].f.spare[5] );
tran (\sa_ctrl[8][11] , \sa_ctrl[8].r.part0[11] );
tran (\sa_ctrl[8][11] , \sa_ctrl[8].f.spare[6] );
tran (\sa_ctrl[8][12] , \sa_ctrl[8].r.part0[12] );
tran (\sa_ctrl[8][12] , \sa_ctrl[8].f.spare[7] );
tran (\sa_ctrl[8][13] , \sa_ctrl[8].r.part0[13] );
tran (\sa_ctrl[8][13] , \sa_ctrl[8].f.spare[8] );
tran (\sa_ctrl[8][14] , \sa_ctrl[8].r.part0[14] );
tran (\sa_ctrl[8][14] , \sa_ctrl[8].f.spare[9] );
tran (\sa_ctrl[8][15] , \sa_ctrl[8].r.part0[15] );
tran (\sa_ctrl[8][15] , \sa_ctrl[8].f.spare[10] );
tran (\sa_ctrl[8][16] , \sa_ctrl[8].r.part0[16] );
tran (\sa_ctrl[8][16] , \sa_ctrl[8].f.spare[11] );
tran (\sa_ctrl[8][17] , \sa_ctrl[8].r.part0[17] );
tran (\sa_ctrl[8][17] , \sa_ctrl[8].f.spare[12] );
tran (\sa_ctrl[8][18] , \sa_ctrl[8].r.part0[18] );
tran (\sa_ctrl[8][18] , \sa_ctrl[8].f.spare[13] );
tran (\sa_ctrl[8][19] , \sa_ctrl[8].r.part0[19] );
tran (\sa_ctrl[8][19] , \sa_ctrl[8].f.spare[14] );
tran (\sa_ctrl[8][20] , \sa_ctrl[8].r.part0[20] );
tran (\sa_ctrl[8][20] , \sa_ctrl[8].f.spare[15] );
tran (\sa_ctrl[8][21] , \sa_ctrl[8].r.part0[21] );
tran (\sa_ctrl[8][21] , \sa_ctrl[8].f.spare[16] );
tran (\sa_ctrl[8][22] , \sa_ctrl[8].r.part0[22] );
tran (\sa_ctrl[8][22] , \sa_ctrl[8].f.spare[17] );
tran (\sa_ctrl[8][23] , \sa_ctrl[8].r.part0[23] );
tran (\sa_ctrl[8][23] , \sa_ctrl[8].f.spare[18] );
tran (\sa_ctrl[8][24] , \sa_ctrl[8].r.part0[24] );
tran (\sa_ctrl[8][24] , \sa_ctrl[8].f.spare[19] );
tran (\sa_ctrl[8][25] , \sa_ctrl[8].r.part0[25] );
tran (\sa_ctrl[8][25] , \sa_ctrl[8].f.spare[20] );
tran (\sa_ctrl[8][26] , \sa_ctrl[8].r.part0[26] );
tran (\sa_ctrl[8][26] , \sa_ctrl[8].f.spare[21] );
tran (\sa_ctrl[8][27] , \sa_ctrl[8].r.part0[27] );
tran (\sa_ctrl[8][27] , \sa_ctrl[8].f.spare[22] );
tran (\sa_ctrl[8][28] , \sa_ctrl[8].r.part0[28] );
tran (\sa_ctrl[8][28] , \sa_ctrl[8].f.spare[23] );
tran (\sa_ctrl[8][29] , \sa_ctrl[8].r.part0[29] );
tran (\sa_ctrl[8][29] , \sa_ctrl[8].f.spare[24] );
tran (\sa_ctrl[8][30] , \sa_ctrl[8].r.part0[30] );
tran (\sa_ctrl[8][30] , \sa_ctrl[8].f.spare[25] );
tran (\sa_ctrl[8][31] , \sa_ctrl[8].r.part0[31] );
tran (\sa_ctrl[8][31] , \sa_ctrl[8].f.spare[26] );
tran (\sa_ctrl[9][0] , \sa_ctrl[9].r.part0[0] );
tran (\sa_ctrl[9][0] , \sa_ctrl[9].f.sa_event_sel[0] );
tran (\sa_ctrl[9][1] , \sa_ctrl[9].r.part0[1] );
tran (\sa_ctrl[9][1] , \sa_ctrl[9].f.sa_event_sel[1] );
tran (\sa_ctrl[9][2] , \sa_ctrl[9].r.part0[2] );
tran (\sa_ctrl[9][2] , \sa_ctrl[9].f.sa_event_sel[2] );
tran (\sa_ctrl[9][3] , \sa_ctrl[9].r.part0[3] );
tran (\sa_ctrl[9][3] , \sa_ctrl[9].f.sa_event_sel[3] );
tran (\sa_ctrl[9][4] , \sa_ctrl[9].r.part0[4] );
tran (\sa_ctrl[9][4] , \sa_ctrl[9].f.sa_event_sel[4] );
tran (\sa_ctrl[9][5] , \sa_ctrl[9].r.part0[5] );
tran (\sa_ctrl[9][5] , \sa_ctrl[9].f.spare[0] );
tran (\sa_ctrl[9][6] , \sa_ctrl[9].r.part0[6] );
tran (\sa_ctrl[9][6] , \sa_ctrl[9].f.spare[1] );
tran (\sa_ctrl[9][7] , \sa_ctrl[9].r.part0[7] );
tran (\sa_ctrl[9][7] , \sa_ctrl[9].f.spare[2] );
tran (\sa_ctrl[9][8] , \sa_ctrl[9].r.part0[8] );
tran (\sa_ctrl[9][8] , \sa_ctrl[9].f.spare[3] );
tran (\sa_ctrl[9][9] , \sa_ctrl[9].r.part0[9] );
tran (\sa_ctrl[9][9] , \sa_ctrl[9].f.spare[4] );
tran (\sa_ctrl[9][10] , \sa_ctrl[9].r.part0[10] );
tran (\sa_ctrl[9][10] , \sa_ctrl[9].f.spare[5] );
tran (\sa_ctrl[9][11] , \sa_ctrl[9].r.part0[11] );
tran (\sa_ctrl[9][11] , \sa_ctrl[9].f.spare[6] );
tran (\sa_ctrl[9][12] , \sa_ctrl[9].r.part0[12] );
tran (\sa_ctrl[9][12] , \sa_ctrl[9].f.spare[7] );
tran (\sa_ctrl[9][13] , \sa_ctrl[9].r.part0[13] );
tran (\sa_ctrl[9][13] , \sa_ctrl[9].f.spare[8] );
tran (\sa_ctrl[9][14] , \sa_ctrl[9].r.part0[14] );
tran (\sa_ctrl[9][14] , \sa_ctrl[9].f.spare[9] );
tran (\sa_ctrl[9][15] , \sa_ctrl[9].r.part0[15] );
tran (\sa_ctrl[9][15] , \sa_ctrl[9].f.spare[10] );
tran (\sa_ctrl[9][16] , \sa_ctrl[9].r.part0[16] );
tran (\sa_ctrl[9][16] , \sa_ctrl[9].f.spare[11] );
tran (\sa_ctrl[9][17] , \sa_ctrl[9].r.part0[17] );
tran (\sa_ctrl[9][17] , \sa_ctrl[9].f.spare[12] );
tran (\sa_ctrl[9][18] , \sa_ctrl[9].r.part0[18] );
tran (\sa_ctrl[9][18] , \sa_ctrl[9].f.spare[13] );
tran (\sa_ctrl[9][19] , \sa_ctrl[9].r.part0[19] );
tran (\sa_ctrl[9][19] , \sa_ctrl[9].f.spare[14] );
tran (\sa_ctrl[9][20] , \sa_ctrl[9].r.part0[20] );
tran (\sa_ctrl[9][20] , \sa_ctrl[9].f.spare[15] );
tran (\sa_ctrl[9][21] , \sa_ctrl[9].r.part0[21] );
tran (\sa_ctrl[9][21] , \sa_ctrl[9].f.spare[16] );
tran (\sa_ctrl[9][22] , \sa_ctrl[9].r.part0[22] );
tran (\sa_ctrl[9][22] , \sa_ctrl[9].f.spare[17] );
tran (\sa_ctrl[9][23] , \sa_ctrl[9].r.part0[23] );
tran (\sa_ctrl[9][23] , \sa_ctrl[9].f.spare[18] );
tran (\sa_ctrl[9][24] , \sa_ctrl[9].r.part0[24] );
tran (\sa_ctrl[9][24] , \sa_ctrl[9].f.spare[19] );
tran (\sa_ctrl[9][25] , \sa_ctrl[9].r.part0[25] );
tran (\sa_ctrl[9][25] , \sa_ctrl[9].f.spare[20] );
tran (\sa_ctrl[9][26] , \sa_ctrl[9].r.part0[26] );
tran (\sa_ctrl[9][26] , \sa_ctrl[9].f.spare[21] );
tran (\sa_ctrl[9][27] , \sa_ctrl[9].r.part0[27] );
tran (\sa_ctrl[9][27] , \sa_ctrl[9].f.spare[22] );
tran (\sa_ctrl[9][28] , \sa_ctrl[9].r.part0[28] );
tran (\sa_ctrl[9][28] , \sa_ctrl[9].f.spare[23] );
tran (\sa_ctrl[9][29] , \sa_ctrl[9].r.part0[29] );
tran (\sa_ctrl[9][29] , \sa_ctrl[9].f.spare[24] );
tran (\sa_ctrl[9][30] , \sa_ctrl[9].r.part0[30] );
tran (\sa_ctrl[9][30] , \sa_ctrl[9].f.spare[25] );
tran (\sa_ctrl[9][31] , \sa_ctrl[9].r.part0[31] );
tran (\sa_ctrl[9][31] , \sa_ctrl[9].f.spare[26] );
tran (\sa_ctrl[10][0] , \sa_ctrl[10].r.part0[0] );
tran (\sa_ctrl[10][0] , \sa_ctrl[10].f.sa_event_sel[0] );
tran (\sa_ctrl[10][1] , \sa_ctrl[10].r.part0[1] );
tran (\sa_ctrl[10][1] , \sa_ctrl[10].f.sa_event_sel[1] );
tran (\sa_ctrl[10][2] , \sa_ctrl[10].r.part0[2] );
tran (\sa_ctrl[10][2] , \sa_ctrl[10].f.sa_event_sel[2] );
tran (\sa_ctrl[10][3] , \sa_ctrl[10].r.part0[3] );
tran (\sa_ctrl[10][3] , \sa_ctrl[10].f.sa_event_sel[3] );
tran (\sa_ctrl[10][4] , \sa_ctrl[10].r.part0[4] );
tran (\sa_ctrl[10][4] , \sa_ctrl[10].f.sa_event_sel[4] );
tran (\sa_ctrl[10][5] , \sa_ctrl[10].r.part0[5] );
tran (\sa_ctrl[10][5] , \sa_ctrl[10].f.spare[0] );
tran (\sa_ctrl[10][6] , \sa_ctrl[10].r.part0[6] );
tran (\sa_ctrl[10][6] , \sa_ctrl[10].f.spare[1] );
tran (\sa_ctrl[10][7] , \sa_ctrl[10].r.part0[7] );
tran (\sa_ctrl[10][7] , \sa_ctrl[10].f.spare[2] );
tran (\sa_ctrl[10][8] , \sa_ctrl[10].r.part0[8] );
tran (\sa_ctrl[10][8] , \sa_ctrl[10].f.spare[3] );
tran (\sa_ctrl[10][9] , \sa_ctrl[10].r.part0[9] );
tran (\sa_ctrl[10][9] , \sa_ctrl[10].f.spare[4] );
tran (\sa_ctrl[10][10] , \sa_ctrl[10].r.part0[10] );
tran (\sa_ctrl[10][10] , \sa_ctrl[10].f.spare[5] );
tran (\sa_ctrl[10][11] , \sa_ctrl[10].r.part0[11] );
tran (\sa_ctrl[10][11] , \sa_ctrl[10].f.spare[6] );
tran (\sa_ctrl[10][12] , \sa_ctrl[10].r.part0[12] );
tran (\sa_ctrl[10][12] , \sa_ctrl[10].f.spare[7] );
tran (\sa_ctrl[10][13] , \sa_ctrl[10].r.part0[13] );
tran (\sa_ctrl[10][13] , \sa_ctrl[10].f.spare[8] );
tran (\sa_ctrl[10][14] , \sa_ctrl[10].r.part0[14] );
tran (\sa_ctrl[10][14] , \sa_ctrl[10].f.spare[9] );
tran (\sa_ctrl[10][15] , \sa_ctrl[10].r.part0[15] );
tran (\sa_ctrl[10][15] , \sa_ctrl[10].f.spare[10] );
tran (\sa_ctrl[10][16] , \sa_ctrl[10].r.part0[16] );
tran (\sa_ctrl[10][16] , \sa_ctrl[10].f.spare[11] );
tran (\sa_ctrl[10][17] , \sa_ctrl[10].r.part0[17] );
tran (\sa_ctrl[10][17] , \sa_ctrl[10].f.spare[12] );
tran (\sa_ctrl[10][18] , \sa_ctrl[10].r.part0[18] );
tran (\sa_ctrl[10][18] , \sa_ctrl[10].f.spare[13] );
tran (\sa_ctrl[10][19] , \sa_ctrl[10].r.part0[19] );
tran (\sa_ctrl[10][19] , \sa_ctrl[10].f.spare[14] );
tran (\sa_ctrl[10][20] , \sa_ctrl[10].r.part0[20] );
tran (\sa_ctrl[10][20] , \sa_ctrl[10].f.spare[15] );
tran (\sa_ctrl[10][21] , \sa_ctrl[10].r.part0[21] );
tran (\sa_ctrl[10][21] , \sa_ctrl[10].f.spare[16] );
tran (\sa_ctrl[10][22] , \sa_ctrl[10].r.part0[22] );
tran (\sa_ctrl[10][22] , \sa_ctrl[10].f.spare[17] );
tran (\sa_ctrl[10][23] , \sa_ctrl[10].r.part0[23] );
tran (\sa_ctrl[10][23] , \sa_ctrl[10].f.spare[18] );
tran (\sa_ctrl[10][24] , \sa_ctrl[10].r.part0[24] );
tran (\sa_ctrl[10][24] , \sa_ctrl[10].f.spare[19] );
tran (\sa_ctrl[10][25] , \sa_ctrl[10].r.part0[25] );
tran (\sa_ctrl[10][25] , \sa_ctrl[10].f.spare[20] );
tran (\sa_ctrl[10][26] , \sa_ctrl[10].r.part0[26] );
tran (\sa_ctrl[10][26] , \sa_ctrl[10].f.spare[21] );
tran (\sa_ctrl[10][27] , \sa_ctrl[10].r.part0[27] );
tran (\sa_ctrl[10][27] , \sa_ctrl[10].f.spare[22] );
tran (\sa_ctrl[10][28] , \sa_ctrl[10].r.part0[28] );
tran (\sa_ctrl[10][28] , \sa_ctrl[10].f.spare[23] );
tran (\sa_ctrl[10][29] , \sa_ctrl[10].r.part0[29] );
tran (\sa_ctrl[10][29] , \sa_ctrl[10].f.spare[24] );
tran (\sa_ctrl[10][30] , \sa_ctrl[10].r.part0[30] );
tran (\sa_ctrl[10][30] , \sa_ctrl[10].f.spare[25] );
tran (\sa_ctrl[10][31] , \sa_ctrl[10].r.part0[31] );
tran (\sa_ctrl[10][31] , \sa_ctrl[10].f.spare[26] );
tran (\sa_ctrl[11][0] , \sa_ctrl[11].r.part0[0] );
tran (\sa_ctrl[11][0] , \sa_ctrl[11].f.sa_event_sel[0] );
tran (\sa_ctrl[11][1] , \sa_ctrl[11].r.part0[1] );
tran (\sa_ctrl[11][1] , \sa_ctrl[11].f.sa_event_sel[1] );
tran (\sa_ctrl[11][2] , \sa_ctrl[11].r.part0[2] );
tran (\sa_ctrl[11][2] , \sa_ctrl[11].f.sa_event_sel[2] );
tran (\sa_ctrl[11][3] , \sa_ctrl[11].r.part0[3] );
tran (\sa_ctrl[11][3] , \sa_ctrl[11].f.sa_event_sel[3] );
tran (\sa_ctrl[11][4] , \sa_ctrl[11].r.part0[4] );
tran (\sa_ctrl[11][4] , \sa_ctrl[11].f.sa_event_sel[4] );
tran (\sa_ctrl[11][5] , \sa_ctrl[11].r.part0[5] );
tran (\sa_ctrl[11][5] , \sa_ctrl[11].f.spare[0] );
tran (\sa_ctrl[11][6] , \sa_ctrl[11].r.part0[6] );
tran (\sa_ctrl[11][6] , \sa_ctrl[11].f.spare[1] );
tran (\sa_ctrl[11][7] , \sa_ctrl[11].r.part0[7] );
tran (\sa_ctrl[11][7] , \sa_ctrl[11].f.spare[2] );
tran (\sa_ctrl[11][8] , \sa_ctrl[11].r.part0[8] );
tran (\sa_ctrl[11][8] , \sa_ctrl[11].f.spare[3] );
tran (\sa_ctrl[11][9] , \sa_ctrl[11].r.part0[9] );
tran (\sa_ctrl[11][9] , \sa_ctrl[11].f.spare[4] );
tran (\sa_ctrl[11][10] , \sa_ctrl[11].r.part0[10] );
tran (\sa_ctrl[11][10] , \sa_ctrl[11].f.spare[5] );
tran (\sa_ctrl[11][11] , \sa_ctrl[11].r.part0[11] );
tran (\sa_ctrl[11][11] , \sa_ctrl[11].f.spare[6] );
tran (\sa_ctrl[11][12] , \sa_ctrl[11].r.part0[12] );
tran (\sa_ctrl[11][12] , \sa_ctrl[11].f.spare[7] );
tran (\sa_ctrl[11][13] , \sa_ctrl[11].r.part0[13] );
tran (\sa_ctrl[11][13] , \sa_ctrl[11].f.spare[8] );
tran (\sa_ctrl[11][14] , \sa_ctrl[11].r.part0[14] );
tran (\sa_ctrl[11][14] , \sa_ctrl[11].f.spare[9] );
tran (\sa_ctrl[11][15] , \sa_ctrl[11].r.part0[15] );
tran (\sa_ctrl[11][15] , \sa_ctrl[11].f.spare[10] );
tran (\sa_ctrl[11][16] , \sa_ctrl[11].r.part0[16] );
tran (\sa_ctrl[11][16] , \sa_ctrl[11].f.spare[11] );
tran (\sa_ctrl[11][17] , \sa_ctrl[11].r.part0[17] );
tran (\sa_ctrl[11][17] , \sa_ctrl[11].f.spare[12] );
tran (\sa_ctrl[11][18] , \sa_ctrl[11].r.part0[18] );
tran (\sa_ctrl[11][18] , \sa_ctrl[11].f.spare[13] );
tran (\sa_ctrl[11][19] , \sa_ctrl[11].r.part0[19] );
tran (\sa_ctrl[11][19] , \sa_ctrl[11].f.spare[14] );
tran (\sa_ctrl[11][20] , \sa_ctrl[11].r.part0[20] );
tran (\sa_ctrl[11][20] , \sa_ctrl[11].f.spare[15] );
tran (\sa_ctrl[11][21] , \sa_ctrl[11].r.part0[21] );
tran (\sa_ctrl[11][21] , \sa_ctrl[11].f.spare[16] );
tran (\sa_ctrl[11][22] , \sa_ctrl[11].r.part0[22] );
tran (\sa_ctrl[11][22] , \sa_ctrl[11].f.spare[17] );
tran (\sa_ctrl[11][23] , \sa_ctrl[11].r.part0[23] );
tran (\sa_ctrl[11][23] , \sa_ctrl[11].f.spare[18] );
tran (\sa_ctrl[11][24] , \sa_ctrl[11].r.part0[24] );
tran (\sa_ctrl[11][24] , \sa_ctrl[11].f.spare[19] );
tran (\sa_ctrl[11][25] , \sa_ctrl[11].r.part0[25] );
tran (\sa_ctrl[11][25] , \sa_ctrl[11].f.spare[20] );
tran (\sa_ctrl[11][26] , \sa_ctrl[11].r.part0[26] );
tran (\sa_ctrl[11][26] , \sa_ctrl[11].f.spare[21] );
tran (\sa_ctrl[11][27] , \sa_ctrl[11].r.part0[27] );
tran (\sa_ctrl[11][27] , \sa_ctrl[11].f.spare[22] );
tran (\sa_ctrl[11][28] , \sa_ctrl[11].r.part0[28] );
tran (\sa_ctrl[11][28] , \sa_ctrl[11].f.spare[23] );
tran (\sa_ctrl[11][29] , \sa_ctrl[11].r.part0[29] );
tran (\sa_ctrl[11][29] , \sa_ctrl[11].f.spare[24] );
tran (\sa_ctrl[11][30] , \sa_ctrl[11].r.part0[30] );
tran (\sa_ctrl[11][30] , \sa_ctrl[11].f.spare[25] );
tran (\sa_ctrl[11][31] , \sa_ctrl[11].r.part0[31] );
tran (\sa_ctrl[11][31] , \sa_ctrl[11].f.spare[26] );
tran (\sa_ctrl[12][0] , \sa_ctrl[12].r.part0[0] );
tran (\sa_ctrl[12][0] , \sa_ctrl[12].f.sa_event_sel[0] );
tran (\sa_ctrl[12][1] , \sa_ctrl[12].r.part0[1] );
tran (\sa_ctrl[12][1] , \sa_ctrl[12].f.sa_event_sel[1] );
tran (\sa_ctrl[12][2] , \sa_ctrl[12].r.part0[2] );
tran (\sa_ctrl[12][2] , \sa_ctrl[12].f.sa_event_sel[2] );
tran (\sa_ctrl[12][3] , \sa_ctrl[12].r.part0[3] );
tran (\sa_ctrl[12][3] , \sa_ctrl[12].f.sa_event_sel[3] );
tran (\sa_ctrl[12][4] , \sa_ctrl[12].r.part0[4] );
tran (\sa_ctrl[12][4] , \sa_ctrl[12].f.sa_event_sel[4] );
tran (\sa_ctrl[12][5] , \sa_ctrl[12].r.part0[5] );
tran (\sa_ctrl[12][5] , \sa_ctrl[12].f.spare[0] );
tran (\sa_ctrl[12][6] , \sa_ctrl[12].r.part0[6] );
tran (\sa_ctrl[12][6] , \sa_ctrl[12].f.spare[1] );
tran (\sa_ctrl[12][7] , \sa_ctrl[12].r.part0[7] );
tran (\sa_ctrl[12][7] , \sa_ctrl[12].f.spare[2] );
tran (\sa_ctrl[12][8] , \sa_ctrl[12].r.part0[8] );
tran (\sa_ctrl[12][8] , \sa_ctrl[12].f.spare[3] );
tran (\sa_ctrl[12][9] , \sa_ctrl[12].r.part0[9] );
tran (\sa_ctrl[12][9] , \sa_ctrl[12].f.spare[4] );
tran (\sa_ctrl[12][10] , \sa_ctrl[12].r.part0[10] );
tran (\sa_ctrl[12][10] , \sa_ctrl[12].f.spare[5] );
tran (\sa_ctrl[12][11] , \sa_ctrl[12].r.part0[11] );
tran (\sa_ctrl[12][11] , \sa_ctrl[12].f.spare[6] );
tran (\sa_ctrl[12][12] , \sa_ctrl[12].r.part0[12] );
tran (\sa_ctrl[12][12] , \sa_ctrl[12].f.spare[7] );
tran (\sa_ctrl[12][13] , \sa_ctrl[12].r.part0[13] );
tran (\sa_ctrl[12][13] , \sa_ctrl[12].f.spare[8] );
tran (\sa_ctrl[12][14] , \sa_ctrl[12].r.part0[14] );
tran (\sa_ctrl[12][14] , \sa_ctrl[12].f.spare[9] );
tran (\sa_ctrl[12][15] , \sa_ctrl[12].r.part0[15] );
tran (\sa_ctrl[12][15] , \sa_ctrl[12].f.spare[10] );
tran (\sa_ctrl[12][16] , \sa_ctrl[12].r.part0[16] );
tran (\sa_ctrl[12][16] , \sa_ctrl[12].f.spare[11] );
tran (\sa_ctrl[12][17] , \sa_ctrl[12].r.part0[17] );
tran (\sa_ctrl[12][17] , \sa_ctrl[12].f.spare[12] );
tran (\sa_ctrl[12][18] , \sa_ctrl[12].r.part0[18] );
tran (\sa_ctrl[12][18] , \sa_ctrl[12].f.spare[13] );
tran (\sa_ctrl[12][19] , \sa_ctrl[12].r.part0[19] );
tran (\sa_ctrl[12][19] , \sa_ctrl[12].f.spare[14] );
tran (\sa_ctrl[12][20] , \sa_ctrl[12].r.part0[20] );
tran (\sa_ctrl[12][20] , \sa_ctrl[12].f.spare[15] );
tran (\sa_ctrl[12][21] , \sa_ctrl[12].r.part0[21] );
tran (\sa_ctrl[12][21] , \sa_ctrl[12].f.spare[16] );
tran (\sa_ctrl[12][22] , \sa_ctrl[12].r.part0[22] );
tran (\sa_ctrl[12][22] , \sa_ctrl[12].f.spare[17] );
tran (\sa_ctrl[12][23] , \sa_ctrl[12].r.part0[23] );
tran (\sa_ctrl[12][23] , \sa_ctrl[12].f.spare[18] );
tran (\sa_ctrl[12][24] , \sa_ctrl[12].r.part0[24] );
tran (\sa_ctrl[12][24] , \sa_ctrl[12].f.spare[19] );
tran (\sa_ctrl[12][25] , \sa_ctrl[12].r.part0[25] );
tran (\sa_ctrl[12][25] , \sa_ctrl[12].f.spare[20] );
tran (\sa_ctrl[12][26] , \sa_ctrl[12].r.part0[26] );
tran (\sa_ctrl[12][26] , \sa_ctrl[12].f.spare[21] );
tran (\sa_ctrl[12][27] , \sa_ctrl[12].r.part0[27] );
tran (\sa_ctrl[12][27] , \sa_ctrl[12].f.spare[22] );
tran (\sa_ctrl[12][28] , \sa_ctrl[12].r.part0[28] );
tran (\sa_ctrl[12][28] , \sa_ctrl[12].f.spare[23] );
tran (\sa_ctrl[12][29] , \sa_ctrl[12].r.part0[29] );
tran (\sa_ctrl[12][29] , \sa_ctrl[12].f.spare[24] );
tran (\sa_ctrl[12][30] , \sa_ctrl[12].r.part0[30] );
tran (\sa_ctrl[12][30] , \sa_ctrl[12].f.spare[25] );
tran (\sa_ctrl[12][31] , \sa_ctrl[12].r.part0[31] );
tran (\sa_ctrl[12][31] , \sa_ctrl[12].f.spare[26] );
tran (\sa_ctrl[13][0] , \sa_ctrl[13].r.part0[0] );
tran (\sa_ctrl[13][0] , \sa_ctrl[13].f.sa_event_sel[0] );
tran (\sa_ctrl[13][1] , \sa_ctrl[13].r.part0[1] );
tran (\sa_ctrl[13][1] , \sa_ctrl[13].f.sa_event_sel[1] );
tran (\sa_ctrl[13][2] , \sa_ctrl[13].r.part0[2] );
tran (\sa_ctrl[13][2] , \sa_ctrl[13].f.sa_event_sel[2] );
tran (\sa_ctrl[13][3] , \sa_ctrl[13].r.part0[3] );
tran (\sa_ctrl[13][3] , \sa_ctrl[13].f.sa_event_sel[3] );
tran (\sa_ctrl[13][4] , \sa_ctrl[13].r.part0[4] );
tran (\sa_ctrl[13][4] , \sa_ctrl[13].f.sa_event_sel[4] );
tran (\sa_ctrl[13][5] , \sa_ctrl[13].r.part0[5] );
tran (\sa_ctrl[13][5] , \sa_ctrl[13].f.spare[0] );
tran (\sa_ctrl[13][6] , \sa_ctrl[13].r.part0[6] );
tran (\sa_ctrl[13][6] , \sa_ctrl[13].f.spare[1] );
tran (\sa_ctrl[13][7] , \sa_ctrl[13].r.part0[7] );
tran (\sa_ctrl[13][7] , \sa_ctrl[13].f.spare[2] );
tran (\sa_ctrl[13][8] , \sa_ctrl[13].r.part0[8] );
tran (\sa_ctrl[13][8] , \sa_ctrl[13].f.spare[3] );
tran (\sa_ctrl[13][9] , \sa_ctrl[13].r.part0[9] );
tran (\sa_ctrl[13][9] , \sa_ctrl[13].f.spare[4] );
tran (\sa_ctrl[13][10] , \sa_ctrl[13].r.part0[10] );
tran (\sa_ctrl[13][10] , \sa_ctrl[13].f.spare[5] );
tran (\sa_ctrl[13][11] , \sa_ctrl[13].r.part0[11] );
tran (\sa_ctrl[13][11] , \sa_ctrl[13].f.spare[6] );
tran (\sa_ctrl[13][12] , \sa_ctrl[13].r.part0[12] );
tran (\sa_ctrl[13][12] , \sa_ctrl[13].f.spare[7] );
tran (\sa_ctrl[13][13] , \sa_ctrl[13].r.part0[13] );
tran (\sa_ctrl[13][13] , \sa_ctrl[13].f.spare[8] );
tran (\sa_ctrl[13][14] , \sa_ctrl[13].r.part0[14] );
tran (\sa_ctrl[13][14] , \sa_ctrl[13].f.spare[9] );
tran (\sa_ctrl[13][15] , \sa_ctrl[13].r.part0[15] );
tran (\sa_ctrl[13][15] , \sa_ctrl[13].f.spare[10] );
tran (\sa_ctrl[13][16] , \sa_ctrl[13].r.part0[16] );
tran (\sa_ctrl[13][16] , \sa_ctrl[13].f.spare[11] );
tran (\sa_ctrl[13][17] , \sa_ctrl[13].r.part0[17] );
tran (\sa_ctrl[13][17] , \sa_ctrl[13].f.spare[12] );
tran (\sa_ctrl[13][18] , \sa_ctrl[13].r.part0[18] );
tran (\sa_ctrl[13][18] , \sa_ctrl[13].f.spare[13] );
tran (\sa_ctrl[13][19] , \sa_ctrl[13].r.part0[19] );
tran (\sa_ctrl[13][19] , \sa_ctrl[13].f.spare[14] );
tran (\sa_ctrl[13][20] , \sa_ctrl[13].r.part0[20] );
tran (\sa_ctrl[13][20] , \sa_ctrl[13].f.spare[15] );
tran (\sa_ctrl[13][21] , \sa_ctrl[13].r.part0[21] );
tran (\sa_ctrl[13][21] , \sa_ctrl[13].f.spare[16] );
tran (\sa_ctrl[13][22] , \sa_ctrl[13].r.part0[22] );
tran (\sa_ctrl[13][22] , \sa_ctrl[13].f.spare[17] );
tran (\sa_ctrl[13][23] , \sa_ctrl[13].r.part0[23] );
tran (\sa_ctrl[13][23] , \sa_ctrl[13].f.spare[18] );
tran (\sa_ctrl[13][24] , \sa_ctrl[13].r.part0[24] );
tran (\sa_ctrl[13][24] , \sa_ctrl[13].f.spare[19] );
tran (\sa_ctrl[13][25] , \sa_ctrl[13].r.part0[25] );
tran (\sa_ctrl[13][25] , \sa_ctrl[13].f.spare[20] );
tran (\sa_ctrl[13][26] , \sa_ctrl[13].r.part0[26] );
tran (\sa_ctrl[13][26] , \sa_ctrl[13].f.spare[21] );
tran (\sa_ctrl[13][27] , \sa_ctrl[13].r.part0[27] );
tran (\sa_ctrl[13][27] , \sa_ctrl[13].f.spare[22] );
tran (\sa_ctrl[13][28] , \sa_ctrl[13].r.part0[28] );
tran (\sa_ctrl[13][28] , \sa_ctrl[13].f.spare[23] );
tran (\sa_ctrl[13][29] , \sa_ctrl[13].r.part0[29] );
tran (\sa_ctrl[13][29] , \sa_ctrl[13].f.spare[24] );
tran (\sa_ctrl[13][30] , \sa_ctrl[13].r.part0[30] );
tran (\sa_ctrl[13][30] , \sa_ctrl[13].f.spare[25] );
tran (\sa_ctrl[13][31] , \sa_ctrl[13].r.part0[31] );
tran (\sa_ctrl[13][31] , \sa_ctrl[13].f.spare[26] );
tran (\sa_ctrl[14][0] , \sa_ctrl[14].r.part0[0] );
tran (\sa_ctrl[14][0] , \sa_ctrl[14].f.sa_event_sel[0] );
tran (\sa_ctrl[14][1] , \sa_ctrl[14].r.part0[1] );
tran (\sa_ctrl[14][1] , \sa_ctrl[14].f.sa_event_sel[1] );
tran (\sa_ctrl[14][2] , \sa_ctrl[14].r.part0[2] );
tran (\sa_ctrl[14][2] , \sa_ctrl[14].f.sa_event_sel[2] );
tran (\sa_ctrl[14][3] , \sa_ctrl[14].r.part0[3] );
tran (\sa_ctrl[14][3] , \sa_ctrl[14].f.sa_event_sel[3] );
tran (\sa_ctrl[14][4] , \sa_ctrl[14].r.part0[4] );
tran (\sa_ctrl[14][4] , \sa_ctrl[14].f.sa_event_sel[4] );
tran (\sa_ctrl[14][5] , \sa_ctrl[14].r.part0[5] );
tran (\sa_ctrl[14][5] , \sa_ctrl[14].f.spare[0] );
tran (\sa_ctrl[14][6] , \sa_ctrl[14].r.part0[6] );
tran (\sa_ctrl[14][6] , \sa_ctrl[14].f.spare[1] );
tran (\sa_ctrl[14][7] , \sa_ctrl[14].r.part0[7] );
tran (\sa_ctrl[14][7] , \sa_ctrl[14].f.spare[2] );
tran (\sa_ctrl[14][8] , \sa_ctrl[14].r.part0[8] );
tran (\sa_ctrl[14][8] , \sa_ctrl[14].f.spare[3] );
tran (\sa_ctrl[14][9] , \sa_ctrl[14].r.part0[9] );
tran (\sa_ctrl[14][9] , \sa_ctrl[14].f.spare[4] );
tran (\sa_ctrl[14][10] , \sa_ctrl[14].r.part0[10] );
tran (\sa_ctrl[14][10] , \sa_ctrl[14].f.spare[5] );
tran (\sa_ctrl[14][11] , \sa_ctrl[14].r.part0[11] );
tran (\sa_ctrl[14][11] , \sa_ctrl[14].f.spare[6] );
tran (\sa_ctrl[14][12] , \sa_ctrl[14].r.part0[12] );
tran (\sa_ctrl[14][12] , \sa_ctrl[14].f.spare[7] );
tran (\sa_ctrl[14][13] , \sa_ctrl[14].r.part0[13] );
tran (\sa_ctrl[14][13] , \sa_ctrl[14].f.spare[8] );
tran (\sa_ctrl[14][14] , \sa_ctrl[14].r.part0[14] );
tran (\sa_ctrl[14][14] , \sa_ctrl[14].f.spare[9] );
tran (\sa_ctrl[14][15] , \sa_ctrl[14].r.part0[15] );
tran (\sa_ctrl[14][15] , \sa_ctrl[14].f.spare[10] );
tran (\sa_ctrl[14][16] , \sa_ctrl[14].r.part0[16] );
tran (\sa_ctrl[14][16] , \sa_ctrl[14].f.spare[11] );
tran (\sa_ctrl[14][17] , \sa_ctrl[14].r.part0[17] );
tran (\sa_ctrl[14][17] , \sa_ctrl[14].f.spare[12] );
tran (\sa_ctrl[14][18] , \sa_ctrl[14].r.part0[18] );
tran (\sa_ctrl[14][18] , \sa_ctrl[14].f.spare[13] );
tran (\sa_ctrl[14][19] , \sa_ctrl[14].r.part0[19] );
tran (\sa_ctrl[14][19] , \sa_ctrl[14].f.spare[14] );
tran (\sa_ctrl[14][20] , \sa_ctrl[14].r.part0[20] );
tran (\sa_ctrl[14][20] , \sa_ctrl[14].f.spare[15] );
tran (\sa_ctrl[14][21] , \sa_ctrl[14].r.part0[21] );
tran (\sa_ctrl[14][21] , \sa_ctrl[14].f.spare[16] );
tran (\sa_ctrl[14][22] , \sa_ctrl[14].r.part0[22] );
tran (\sa_ctrl[14][22] , \sa_ctrl[14].f.spare[17] );
tran (\sa_ctrl[14][23] , \sa_ctrl[14].r.part0[23] );
tran (\sa_ctrl[14][23] , \sa_ctrl[14].f.spare[18] );
tran (\sa_ctrl[14][24] , \sa_ctrl[14].r.part0[24] );
tran (\sa_ctrl[14][24] , \sa_ctrl[14].f.spare[19] );
tran (\sa_ctrl[14][25] , \sa_ctrl[14].r.part0[25] );
tran (\sa_ctrl[14][25] , \sa_ctrl[14].f.spare[20] );
tran (\sa_ctrl[14][26] , \sa_ctrl[14].r.part0[26] );
tran (\sa_ctrl[14][26] , \sa_ctrl[14].f.spare[21] );
tran (\sa_ctrl[14][27] , \sa_ctrl[14].r.part0[27] );
tran (\sa_ctrl[14][27] , \sa_ctrl[14].f.spare[22] );
tran (\sa_ctrl[14][28] , \sa_ctrl[14].r.part0[28] );
tran (\sa_ctrl[14][28] , \sa_ctrl[14].f.spare[23] );
tran (\sa_ctrl[14][29] , \sa_ctrl[14].r.part0[29] );
tran (\sa_ctrl[14][29] , \sa_ctrl[14].f.spare[24] );
tran (\sa_ctrl[14][30] , \sa_ctrl[14].r.part0[30] );
tran (\sa_ctrl[14][30] , \sa_ctrl[14].f.spare[25] );
tran (\sa_ctrl[14][31] , \sa_ctrl[14].r.part0[31] );
tran (\sa_ctrl[14][31] , \sa_ctrl[14].f.spare[26] );
tran (\sa_ctrl[15][0] , \sa_ctrl[15].r.part0[0] );
tran (\sa_ctrl[15][0] , \sa_ctrl[15].f.sa_event_sel[0] );
tran (\sa_ctrl[15][1] , \sa_ctrl[15].r.part0[1] );
tran (\sa_ctrl[15][1] , \sa_ctrl[15].f.sa_event_sel[1] );
tran (\sa_ctrl[15][2] , \sa_ctrl[15].r.part0[2] );
tran (\sa_ctrl[15][2] , \sa_ctrl[15].f.sa_event_sel[2] );
tran (\sa_ctrl[15][3] , \sa_ctrl[15].r.part0[3] );
tran (\sa_ctrl[15][3] , \sa_ctrl[15].f.sa_event_sel[3] );
tran (\sa_ctrl[15][4] , \sa_ctrl[15].r.part0[4] );
tran (\sa_ctrl[15][4] , \sa_ctrl[15].f.sa_event_sel[4] );
tran (\sa_ctrl[15][5] , \sa_ctrl[15].r.part0[5] );
tran (\sa_ctrl[15][5] , \sa_ctrl[15].f.spare[0] );
tran (\sa_ctrl[15][6] , \sa_ctrl[15].r.part0[6] );
tran (\sa_ctrl[15][6] , \sa_ctrl[15].f.spare[1] );
tran (\sa_ctrl[15][7] , \sa_ctrl[15].r.part0[7] );
tran (\sa_ctrl[15][7] , \sa_ctrl[15].f.spare[2] );
tran (\sa_ctrl[15][8] , \sa_ctrl[15].r.part0[8] );
tran (\sa_ctrl[15][8] , \sa_ctrl[15].f.spare[3] );
tran (\sa_ctrl[15][9] , \sa_ctrl[15].r.part0[9] );
tran (\sa_ctrl[15][9] , \sa_ctrl[15].f.spare[4] );
tran (\sa_ctrl[15][10] , \sa_ctrl[15].r.part0[10] );
tran (\sa_ctrl[15][10] , \sa_ctrl[15].f.spare[5] );
tran (\sa_ctrl[15][11] , \sa_ctrl[15].r.part0[11] );
tran (\sa_ctrl[15][11] , \sa_ctrl[15].f.spare[6] );
tran (\sa_ctrl[15][12] , \sa_ctrl[15].r.part0[12] );
tran (\sa_ctrl[15][12] , \sa_ctrl[15].f.spare[7] );
tran (\sa_ctrl[15][13] , \sa_ctrl[15].r.part0[13] );
tran (\sa_ctrl[15][13] , \sa_ctrl[15].f.spare[8] );
tran (\sa_ctrl[15][14] , \sa_ctrl[15].r.part0[14] );
tran (\sa_ctrl[15][14] , \sa_ctrl[15].f.spare[9] );
tran (\sa_ctrl[15][15] , \sa_ctrl[15].r.part0[15] );
tran (\sa_ctrl[15][15] , \sa_ctrl[15].f.spare[10] );
tran (\sa_ctrl[15][16] , \sa_ctrl[15].r.part0[16] );
tran (\sa_ctrl[15][16] , \sa_ctrl[15].f.spare[11] );
tran (\sa_ctrl[15][17] , \sa_ctrl[15].r.part0[17] );
tran (\sa_ctrl[15][17] , \sa_ctrl[15].f.spare[12] );
tran (\sa_ctrl[15][18] , \sa_ctrl[15].r.part0[18] );
tran (\sa_ctrl[15][18] , \sa_ctrl[15].f.spare[13] );
tran (\sa_ctrl[15][19] , \sa_ctrl[15].r.part0[19] );
tran (\sa_ctrl[15][19] , \sa_ctrl[15].f.spare[14] );
tran (\sa_ctrl[15][20] , \sa_ctrl[15].r.part0[20] );
tran (\sa_ctrl[15][20] , \sa_ctrl[15].f.spare[15] );
tran (\sa_ctrl[15][21] , \sa_ctrl[15].r.part0[21] );
tran (\sa_ctrl[15][21] , \sa_ctrl[15].f.spare[16] );
tran (\sa_ctrl[15][22] , \sa_ctrl[15].r.part0[22] );
tran (\sa_ctrl[15][22] , \sa_ctrl[15].f.spare[17] );
tran (\sa_ctrl[15][23] , \sa_ctrl[15].r.part0[23] );
tran (\sa_ctrl[15][23] , \sa_ctrl[15].f.spare[18] );
tran (\sa_ctrl[15][24] , \sa_ctrl[15].r.part0[24] );
tran (\sa_ctrl[15][24] , \sa_ctrl[15].f.spare[19] );
tran (\sa_ctrl[15][25] , \sa_ctrl[15].r.part0[25] );
tran (\sa_ctrl[15][25] , \sa_ctrl[15].f.spare[20] );
tran (\sa_ctrl[15][26] , \sa_ctrl[15].r.part0[26] );
tran (\sa_ctrl[15][26] , \sa_ctrl[15].f.spare[21] );
tran (\sa_ctrl[15][27] , \sa_ctrl[15].r.part0[27] );
tran (\sa_ctrl[15][27] , \sa_ctrl[15].f.spare[22] );
tran (\sa_ctrl[15][28] , \sa_ctrl[15].r.part0[28] );
tran (\sa_ctrl[15][28] , \sa_ctrl[15].f.spare[23] );
tran (\sa_ctrl[15][29] , \sa_ctrl[15].r.part0[29] );
tran (\sa_ctrl[15][29] , \sa_ctrl[15].f.spare[24] );
tran (\sa_ctrl[15][30] , \sa_ctrl[15].r.part0[30] );
tran (\sa_ctrl[15][30] , \sa_ctrl[15].f.spare[25] );
tran (\sa_ctrl[15][31] , \sa_ctrl[15].r.part0[31] );
tran (\sa_ctrl[15][31] , \sa_ctrl[15].f.spare[26] );
tran (\sa_ctrl[16][0] , \sa_ctrl[16].r.part0[0] );
tran (\sa_ctrl[16][0] , \sa_ctrl[16].f.sa_event_sel[0] );
tran (\sa_ctrl[16][1] , \sa_ctrl[16].r.part0[1] );
tran (\sa_ctrl[16][1] , \sa_ctrl[16].f.sa_event_sel[1] );
tran (\sa_ctrl[16][2] , \sa_ctrl[16].r.part0[2] );
tran (\sa_ctrl[16][2] , \sa_ctrl[16].f.sa_event_sel[2] );
tran (\sa_ctrl[16][3] , \sa_ctrl[16].r.part0[3] );
tran (\sa_ctrl[16][3] , \sa_ctrl[16].f.sa_event_sel[3] );
tran (\sa_ctrl[16][4] , \sa_ctrl[16].r.part0[4] );
tran (\sa_ctrl[16][4] , \sa_ctrl[16].f.sa_event_sel[4] );
tran (\sa_ctrl[16][5] , \sa_ctrl[16].r.part0[5] );
tran (\sa_ctrl[16][5] , \sa_ctrl[16].f.spare[0] );
tran (\sa_ctrl[16][6] , \sa_ctrl[16].r.part0[6] );
tran (\sa_ctrl[16][6] , \sa_ctrl[16].f.spare[1] );
tran (\sa_ctrl[16][7] , \sa_ctrl[16].r.part0[7] );
tran (\sa_ctrl[16][7] , \sa_ctrl[16].f.spare[2] );
tran (\sa_ctrl[16][8] , \sa_ctrl[16].r.part0[8] );
tran (\sa_ctrl[16][8] , \sa_ctrl[16].f.spare[3] );
tran (\sa_ctrl[16][9] , \sa_ctrl[16].r.part0[9] );
tran (\sa_ctrl[16][9] , \sa_ctrl[16].f.spare[4] );
tran (\sa_ctrl[16][10] , \sa_ctrl[16].r.part0[10] );
tran (\sa_ctrl[16][10] , \sa_ctrl[16].f.spare[5] );
tran (\sa_ctrl[16][11] , \sa_ctrl[16].r.part0[11] );
tran (\sa_ctrl[16][11] , \sa_ctrl[16].f.spare[6] );
tran (\sa_ctrl[16][12] , \sa_ctrl[16].r.part0[12] );
tran (\sa_ctrl[16][12] , \sa_ctrl[16].f.spare[7] );
tran (\sa_ctrl[16][13] , \sa_ctrl[16].r.part0[13] );
tran (\sa_ctrl[16][13] , \sa_ctrl[16].f.spare[8] );
tran (\sa_ctrl[16][14] , \sa_ctrl[16].r.part0[14] );
tran (\sa_ctrl[16][14] , \sa_ctrl[16].f.spare[9] );
tran (\sa_ctrl[16][15] , \sa_ctrl[16].r.part0[15] );
tran (\sa_ctrl[16][15] , \sa_ctrl[16].f.spare[10] );
tran (\sa_ctrl[16][16] , \sa_ctrl[16].r.part0[16] );
tran (\sa_ctrl[16][16] , \sa_ctrl[16].f.spare[11] );
tran (\sa_ctrl[16][17] , \sa_ctrl[16].r.part0[17] );
tran (\sa_ctrl[16][17] , \sa_ctrl[16].f.spare[12] );
tran (\sa_ctrl[16][18] , \sa_ctrl[16].r.part0[18] );
tran (\sa_ctrl[16][18] , \sa_ctrl[16].f.spare[13] );
tran (\sa_ctrl[16][19] , \sa_ctrl[16].r.part0[19] );
tran (\sa_ctrl[16][19] , \sa_ctrl[16].f.spare[14] );
tran (\sa_ctrl[16][20] , \sa_ctrl[16].r.part0[20] );
tran (\sa_ctrl[16][20] , \sa_ctrl[16].f.spare[15] );
tran (\sa_ctrl[16][21] , \sa_ctrl[16].r.part0[21] );
tran (\sa_ctrl[16][21] , \sa_ctrl[16].f.spare[16] );
tran (\sa_ctrl[16][22] , \sa_ctrl[16].r.part0[22] );
tran (\sa_ctrl[16][22] , \sa_ctrl[16].f.spare[17] );
tran (\sa_ctrl[16][23] , \sa_ctrl[16].r.part0[23] );
tran (\sa_ctrl[16][23] , \sa_ctrl[16].f.spare[18] );
tran (\sa_ctrl[16][24] , \sa_ctrl[16].r.part0[24] );
tran (\sa_ctrl[16][24] , \sa_ctrl[16].f.spare[19] );
tran (\sa_ctrl[16][25] , \sa_ctrl[16].r.part0[25] );
tran (\sa_ctrl[16][25] , \sa_ctrl[16].f.spare[20] );
tran (\sa_ctrl[16][26] , \sa_ctrl[16].r.part0[26] );
tran (\sa_ctrl[16][26] , \sa_ctrl[16].f.spare[21] );
tran (\sa_ctrl[16][27] , \sa_ctrl[16].r.part0[27] );
tran (\sa_ctrl[16][27] , \sa_ctrl[16].f.spare[22] );
tran (\sa_ctrl[16][28] , \sa_ctrl[16].r.part0[28] );
tran (\sa_ctrl[16][28] , \sa_ctrl[16].f.spare[23] );
tran (\sa_ctrl[16][29] , \sa_ctrl[16].r.part0[29] );
tran (\sa_ctrl[16][29] , \sa_ctrl[16].f.spare[24] );
tran (\sa_ctrl[16][30] , \sa_ctrl[16].r.part0[30] );
tran (\sa_ctrl[16][30] , \sa_ctrl[16].f.spare[25] );
tran (\sa_ctrl[16][31] , \sa_ctrl[16].r.part0[31] );
tran (\sa_ctrl[16][31] , \sa_ctrl[16].f.spare[26] );
tran (\sa_ctrl[17][0] , \sa_ctrl[17].r.part0[0] );
tran (\sa_ctrl[17][0] , \sa_ctrl[17].f.sa_event_sel[0] );
tran (\sa_ctrl[17][1] , \sa_ctrl[17].r.part0[1] );
tran (\sa_ctrl[17][1] , \sa_ctrl[17].f.sa_event_sel[1] );
tran (\sa_ctrl[17][2] , \sa_ctrl[17].r.part0[2] );
tran (\sa_ctrl[17][2] , \sa_ctrl[17].f.sa_event_sel[2] );
tran (\sa_ctrl[17][3] , \sa_ctrl[17].r.part0[3] );
tran (\sa_ctrl[17][3] , \sa_ctrl[17].f.sa_event_sel[3] );
tran (\sa_ctrl[17][4] , \sa_ctrl[17].r.part0[4] );
tran (\sa_ctrl[17][4] , \sa_ctrl[17].f.sa_event_sel[4] );
tran (\sa_ctrl[17][5] , \sa_ctrl[17].r.part0[5] );
tran (\sa_ctrl[17][5] , \sa_ctrl[17].f.spare[0] );
tran (\sa_ctrl[17][6] , \sa_ctrl[17].r.part0[6] );
tran (\sa_ctrl[17][6] , \sa_ctrl[17].f.spare[1] );
tran (\sa_ctrl[17][7] , \sa_ctrl[17].r.part0[7] );
tran (\sa_ctrl[17][7] , \sa_ctrl[17].f.spare[2] );
tran (\sa_ctrl[17][8] , \sa_ctrl[17].r.part0[8] );
tran (\sa_ctrl[17][8] , \sa_ctrl[17].f.spare[3] );
tran (\sa_ctrl[17][9] , \sa_ctrl[17].r.part0[9] );
tran (\sa_ctrl[17][9] , \sa_ctrl[17].f.spare[4] );
tran (\sa_ctrl[17][10] , \sa_ctrl[17].r.part0[10] );
tran (\sa_ctrl[17][10] , \sa_ctrl[17].f.spare[5] );
tran (\sa_ctrl[17][11] , \sa_ctrl[17].r.part0[11] );
tran (\sa_ctrl[17][11] , \sa_ctrl[17].f.spare[6] );
tran (\sa_ctrl[17][12] , \sa_ctrl[17].r.part0[12] );
tran (\sa_ctrl[17][12] , \sa_ctrl[17].f.spare[7] );
tran (\sa_ctrl[17][13] , \sa_ctrl[17].r.part0[13] );
tran (\sa_ctrl[17][13] , \sa_ctrl[17].f.spare[8] );
tran (\sa_ctrl[17][14] , \sa_ctrl[17].r.part0[14] );
tran (\sa_ctrl[17][14] , \sa_ctrl[17].f.spare[9] );
tran (\sa_ctrl[17][15] , \sa_ctrl[17].r.part0[15] );
tran (\sa_ctrl[17][15] , \sa_ctrl[17].f.spare[10] );
tran (\sa_ctrl[17][16] , \sa_ctrl[17].r.part0[16] );
tran (\sa_ctrl[17][16] , \sa_ctrl[17].f.spare[11] );
tran (\sa_ctrl[17][17] , \sa_ctrl[17].r.part0[17] );
tran (\sa_ctrl[17][17] , \sa_ctrl[17].f.spare[12] );
tran (\sa_ctrl[17][18] , \sa_ctrl[17].r.part0[18] );
tran (\sa_ctrl[17][18] , \sa_ctrl[17].f.spare[13] );
tran (\sa_ctrl[17][19] , \sa_ctrl[17].r.part0[19] );
tran (\sa_ctrl[17][19] , \sa_ctrl[17].f.spare[14] );
tran (\sa_ctrl[17][20] , \sa_ctrl[17].r.part0[20] );
tran (\sa_ctrl[17][20] , \sa_ctrl[17].f.spare[15] );
tran (\sa_ctrl[17][21] , \sa_ctrl[17].r.part0[21] );
tran (\sa_ctrl[17][21] , \sa_ctrl[17].f.spare[16] );
tran (\sa_ctrl[17][22] , \sa_ctrl[17].r.part0[22] );
tran (\sa_ctrl[17][22] , \sa_ctrl[17].f.spare[17] );
tran (\sa_ctrl[17][23] , \sa_ctrl[17].r.part0[23] );
tran (\sa_ctrl[17][23] , \sa_ctrl[17].f.spare[18] );
tran (\sa_ctrl[17][24] , \sa_ctrl[17].r.part0[24] );
tran (\sa_ctrl[17][24] , \sa_ctrl[17].f.spare[19] );
tran (\sa_ctrl[17][25] , \sa_ctrl[17].r.part0[25] );
tran (\sa_ctrl[17][25] , \sa_ctrl[17].f.spare[20] );
tran (\sa_ctrl[17][26] , \sa_ctrl[17].r.part0[26] );
tran (\sa_ctrl[17][26] , \sa_ctrl[17].f.spare[21] );
tran (\sa_ctrl[17][27] , \sa_ctrl[17].r.part0[27] );
tran (\sa_ctrl[17][27] , \sa_ctrl[17].f.spare[22] );
tran (\sa_ctrl[17][28] , \sa_ctrl[17].r.part0[28] );
tran (\sa_ctrl[17][28] , \sa_ctrl[17].f.spare[23] );
tran (\sa_ctrl[17][29] , \sa_ctrl[17].r.part0[29] );
tran (\sa_ctrl[17][29] , \sa_ctrl[17].f.spare[24] );
tran (\sa_ctrl[17][30] , \sa_ctrl[17].r.part0[30] );
tran (\sa_ctrl[17][30] , \sa_ctrl[17].f.spare[25] );
tran (\sa_ctrl[17][31] , \sa_ctrl[17].r.part0[31] );
tran (\sa_ctrl[17][31] , \sa_ctrl[17].f.spare[26] );
tran (\sa_ctrl[18][0] , \sa_ctrl[18].r.part0[0] );
tran (\sa_ctrl[18][0] , \sa_ctrl[18].f.sa_event_sel[0] );
tran (\sa_ctrl[18][1] , \sa_ctrl[18].r.part0[1] );
tran (\sa_ctrl[18][1] , \sa_ctrl[18].f.sa_event_sel[1] );
tran (\sa_ctrl[18][2] , \sa_ctrl[18].r.part0[2] );
tran (\sa_ctrl[18][2] , \sa_ctrl[18].f.sa_event_sel[2] );
tran (\sa_ctrl[18][3] , \sa_ctrl[18].r.part0[3] );
tran (\sa_ctrl[18][3] , \sa_ctrl[18].f.sa_event_sel[3] );
tran (\sa_ctrl[18][4] , \sa_ctrl[18].r.part0[4] );
tran (\sa_ctrl[18][4] , \sa_ctrl[18].f.sa_event_sel[4] );
tran (\sa_ctrl[18][5] , \sa_ctrl[18].r.part0[5] );
tran (\sa_ctrl[18][5] , \sa_ctrl[18].f.spare[0] );
tran (\sa_ctrl[18][6] , \sa_ctrl[18].r.part0[6] );
tran (\sa_ctrl[18][6] , \sa_ctrl[18].f.spare[1] );
tran (\sa_ctrl[18][7] , \sa_ctrl[18].r.part0[7] );
tran (\sa_ctrl[18][7] , \sa_ctrl[18].f.spare[2] );
tran (\sa_ctrl[18][8] , \sa_ctrl[18].r.part0[8] );
tran (\sa_ctrl[18][8] , \sa_ctrl[18].f.spare[3] );
tran (\sa_ctrl[18][9] , \sa_ctrl[18].r.part0[9] );
tran (\sa_ctrl[18][9] , \sa_ctrl[18].f.spare[4] );
tran (\sa_ctrl[18][10] , \sa_ctrl[18].r.part0[10] );
tran (\sa_ctrl[18][10] , \sa_ctrl[18].f.spare[5] );
tran (\sa_ctrl[18][11] , \sa_ctrl[18].r.part0[11] );
tran (\sa_ctrl[18][11] , \sa_ctrl[18].f.spare[6] );
tran (\sa_ctrl[18][12] , \sa_ctrl[18].r.part0[12] );
tran (\sa_ctrl[18][12] , \sa_ctrl[18].f.spare[7] );
tran (\sa_ctrl[18][13] , \sa_ctrl[18].r.part0[13] );
tran (\sa_ctrl[18][13] , \sa_ctrl[18].f.spare[8] );
tran (\sa_ctrl[18][14] , \sa_ctrl[18].r.part0[14] );
tran (\sa_ctrl[18][14] , \sa_ctrl[18].f.spare[9] );
tran (\sa_ctrl[18][15] , \sa_ctrl[18].r.part0[15] );
tran (\sa_ctrl[18][15] , \sa_ctrl[18].f.spare[10] );
tran (\sa_ctrl[18][16] , \sa_ctrl[18].r.part0[16] );
tran (\sa_ctrl[18][16] , \sa_ctrl[18].f.spare[11] );
tran (\sa_ctrl[18][17] , \sa_ctrl[18].r.part0[17] );
tran (\sa_ctrl[18][17] , \sa_ctrl[18].f.spare[12] );
tran (\sa_ctrl[18][18] , \sa_ctrl[18].r.part0[18] );
tran (\sa_ctrl[18][18] , \sa_ctrl[18].f.spare[13] );
tran (\sa_ctrl[18][19] , \sa_ctrl[18].r.part0[19] );
tran (\sa_ctrl[18][19] , \sa_ctrl[18].f.spare[14] );
tran (\sa_ctrl[18][20] , \sa_ctrl[18].r.part0[20] );
tran (\sa_ctrl[18][20] , \sa_ctrl[18].f.spare[15] );
tran (\sa_ctrl[18][21] , \sa_ctrl[18].r.part0[21] );
tran (\sa_ctrl[18][21] , \sa_ctrl[18].f.spare[16] );
tran (\sa_ctrl[18][22] , \sa_ctrl[18].r.part0[22] );
tran (\sa_ctrl[18][22] , \sa_ctrl[18].f.spare[17] );
tran (\sa_ctrl[18][23] , \sa_ctrl[18].r.part0[23] );
tran (\sa_ctrl[18][23] , \sa_ctrl[18].f.spare[18] );
tran (\sa_ctrl[18][24] , \sa_ctrl[18].r.part0[24] );
tran (\sa_ctrl[18][24] , \sa_ctrl[18].f.spare[19] );
tran (\sa_ctrl[18][25] , \sa_ctrl[18].r.part0[25] );
tran (\sa_ctrl[18][25] , \sa_ctrl[18].f.spare[20] );
tran (\sa_ctrl[18][26] , \sa_ctrl[18].r.part0[26] );
tran (\sa_ctrl[18][26] , \sa_ctrl[18].f.spare[21] );
tran (\sa_ctrl[18][27] , \sa_ctrl[18].r.part0[27] );
tran (\sa_ctrl[18][27] , \sa_ctrl[18].f.spare[22] );
tran (\sa_ctrl[18][28] , \sa_ctrl[18].r.part0[28] );
tran (\sa_ctrl[18][28] , \sa_ctrl[18].f.spare[23] );
tran (\sa_ctrl[18][29] , \sa_ctrl[18].r.part0[29] );
tran (\sa_ctrl[18][29] , \sa_ctrl[18].f.spare[24] );
tran (\sa_ctrl[18][30] , \sa_ctrl[18].r.part0[30] );
tran (\sa_ctrl[18][30] , \sa_ctrl[18].f.spare[25] );
tran (\sa_ctrl[18][31] , \sa_ctrl[18].r.part0[31] );
tran (\sa_ctrl[18][31] , \sa_ctrl[18].f.spare[26] );
tran (\sa_ctrl[19][0] , \sa_ctrl[19].r.part0[0] );
tran (\sa_ctrl[19][0] , \sa_ctrl[19].f.sa_event_sel[0] );
tran (\sa_ctrl[19][1] , \sa_ctrl[19].r.part0[1] );
tran (\sa_ctrl[19][1] , \sa_ctrl[19].f.sa_event_sel[1] );
tran (\sa_ctrl[19][2] , \sa_ctrl[19].r.part0[2] );
tran (\sa_ctrl[19][2] , \sa_ctrl[19].f.sa_event_sel[2] );
tran (\sa_ctrl[19][3] , \sa_ctrl[19].r.part0[3] );
tran (\sa_ctrl[19][3] , \sa_ctrl[19].f.sa_event_sel[3] );
tran (\sa_ctrl[19][4] , \sa_ctrl[19].r.part0[4] );
tran (\sa_ctrl[19][4] , \sa_ctrl[19].f.sa_event_sel[4] );
tran (\sa_ctrl[19][5] , \sa_ctrl[19].r.part0[5] );
tran (\sa_ctrl[19][5] , \sa_ctrl[19].f.spare[0] );
tran (\sa_ctrl[19][6] , \sa_ctrl[19].r.part0[6] );
tran (\sa_ctrl[19][6] , \sa_ctrl[19].f.spare[1] );
tran (\sa_ctrl[19][7] , \sa_ctrl[19].r.part0[7] );
tran (\sa_ctrl[19][7] , \sa_ctrl[19].f.spare[2] );
tran (\sa_ctrl[19][8] , \sa_ctrl[19].r.part0[8] );
tran (\sa_ctrl[19][8] , \sa_ctrl[19].f.spare[3] );
tran (\sa_ctrl[19][9] , \sa_ctrl[19].r.part0[9] );
tran (\sa_ctrl[19][9] , \sa_ctrl[19].f.spare[4] );
tran (\sa_ctrl[19][10] , \sa_ctrl[19].r.part0[10] );
tran (\sa_ctrl[19][10] , \sa_ctrl[19].f.spare[5] );
tran (\sa_ctrl[19][11] , \sa_ctrl[19].r.part0[11] );
tran (\sa_ctrl[19][11] , \sa_ctrl[19].f.spare[6] );
tran (\sa_ctrl[19][12] , \sa_ctrl[19].r.part0[12] );
tran (\sa_ctrl[19][12] , \sa_ctrl[19].f.spare[7] );
tran (\sa_ctrl[19][13] , \sa_ctrl[19].r.part0[13] );
tran (\sa_ctrl[19][13] , \sa_ctrl[19].f.spare[8] );
tran (\sa_ctrl[19][14] , \sa_ctrl[19].r.part0[14] );
tran (\sa_ctrl[19][14] , \sa_ctrl[19].f.spare[9] );
tran (\sa_ctrl[19][15] , \sa_ctrl[19].r.part0[15] );
tran (\sa_ctrl[19][15] , \sa_ctrl[19].f.spare[10] );
tran (\sa_ctrl[19][16] , \sa_ctrl[19].r.part0[16] );
tran (\sa_ctrl[19][16] , \sa_ctrl[19].f.spare[11] );
tran (\sa_ctrl[19][17] , \sa_ctrl[19].r.part0[17] );
tran (\sa_ctrl[19][17] , \sa_ctrl[19].f.spare[12] );
tran (\sa_ctrl[19][18] , \sa_ctrl[19].r.part0[18] );
tran (\sa_ctrl[19][18] , \sa_ctrl[19].f.spare[13] );
tran (\sa_ctrl[19][19] , \sa_ctrl[19].r.part0[19] );
tran (\sa_ctrl[19][19] , \sa_ctrl[19].f.spare[14] );
tran (\sa_ctrl[19][20] , \sa_ctrl[19].r.part0[20] );
tran (\sa_ctrl[19][20] , \sa_ctrl[19].f.spare[15] );
tran (\sa_ctrl[19][21] , \sa_ctrl[19].r.part0[21] );
tran (\sa_ctrl[19][21] , \sa_ctrl[19].f.spare[16] );
tran (\sa_ctrl[19][22] , \sa_ctrl[19].r.part0[22] );
tran (\sa_ctrl[19][22] , \sa_ctrl[19].f.spare[17] );
tran (\sa_ctrl[19][23] , \sa_ctrl[19].r.part0[23] );
tran (\sa_ctrl[19][23] , \sa_ctrl[19].f.spare[18] );
tran (\sa_ctrl[19][24] , \sa_ctrl[19].r.part0[24] );
tran (\sa_ctrl[19][24] , \sa_ctrl[19].f.spare[19] );
tran (\sa_ctrl[19][25] , \sa_ctrl[19].r.part0[25] );
tran (\sa_ctrl[19][25] , \sa_ctrl[19].f.spare[20] );
tran (\sa_ctrl[19][26] , \sa_ctrl[19].r.part0[26] );
tran (\sa_ctrl[19][26] , \sa_ctrl[19].f.spare[21] );
tran (\sa_ctrl[19][27] , \sa_ctrl[19].r.part0[27] );
tran (\sa_ctrl[19][27] , \sa_ctrl[19].f.spare[22] );
tran (\sa_ctrl[19][28] , \sa_ctrl[19].r.part0[28] );
tran (\sa_ctrl[19][28] , \sa_ctrl[19].f.spare[23] );
tran (\sa_ctrl[19][29] , \sa_ctrl[19].r.part0[29] );
tran (\sa_ctrl[19][29] , \sa_ctrl[19].f.spare[24] );
tran (\sa_ctrl[19][30] , \sa_ctrl[19].r.part0[30] );
tran (\sa_ctrl[19][30] , \sa_ctrl[19].f.spare[25] );
tran (\sa_ctrl[19][31] , \sa_ctrl[19].r.part0[31] );
tran (\sa_ctrl[19][31] , \sa_ctrl[19].f.spare[26] );
tran (\sa_ctrl[20][0] , \sa_ctrl[20].r.part0[0] );
tran (\sa_ctrl[20][0] , \sa_ctrl[20].f.sa_event_sel[0] );
tran (\sa_ctrl[20][1] , \sa_ctrl[20].r.part0[1] );
tran (\sa_ctrl[20][1] , \sa_ctrl[20].f.sa_event_sel[1] );
tran (\sa_ctrl[20][2] , \sa_ctrl[20].r.part0[2] );
tran (\sa_ctrl[20][2] , \sa_ctrl[20].f.sa_event_sel[2] );
tran (\sa_ctrl[20][3] , \sa_ctrl[20].r.part0[3] );
tran (\sa_ctrl[20][3] , \sa_ctrl[20].f.sa_event_sel[3] );
tran (\sa_ctrl[20][4] , \sa_ctrl[20].r.part0[4] );
tran (\sa_ctrl[20][4] , \sa_ctrl[20].f.sa_event_sel[4] );
tran (\sa_ctrl[20][5] , \sa_ctrl[20].r.part0[5] );
tran (\sa_ctrl[20][5] , \sa_ctrl[20].f.spare[0] );
tran (\sa_ctrl[20][6] , \sa_ctrl[20].r.part0[6] );
tran (\sa_ctrl[20][6] , \sa_ctrl[20].f.spare[1] );
tran (\sa_ctrl[20][7] , \sa_ctrl[20].r.part0[7] );
tran (\sa_ctrl[20][7] , \sa_ctrl[20].f.spare[2] );
tran (\sa_ctrl[20][8] , \sa_ctrl[20].r.part0[8] );
tran (\sa_ctrl[20][8] , \sa_ctrl[20].f.spare[3] );
tran (\sa_ctrl[20][9] , \sa_ctrl[20].r.part0[9] );
tran (\sa_ctrl[20][9] , \sa_ctrl[20].f.spare[4] );
tran (\sa_ctrl[20][10] , \sa_ctrl[20].r.part0[10] );
tran (\sa_ctrl[20][10] , \sa_ctrl[20].f.spare[5] );
tran (\sa_ctrl[20][11] , \sa_ctrl[20].r.part0[11] );
tran (\sa_ctrl[20][11] , \sa_ctrl[20].f.spare[6] );
tran (\sa_ctrl[20][12] , \sa_ctrl[20].r.part0[12] );
tran (\sa_ctrl[20][12] , \sa_ctrl[20].f.spare[7] );
tran (\sa_ctrl[20][13] , \sa_ctrl[20].r.part0[13] );
tran (\sa_ctrl[20][13] , \sa_ctrl[20].f.spare[8] );
tran (\sa_ctrl[20][14] , \sa_ctrl[20].r.part0[14] );
tran (\sa_ctrl[20][14] , \sa_ctrl[20].f.spare[9] );
tran (\sa_ctrl[20][15] , \sa_ctrl[20].r.part0[15] );
tran (\sa_ctrl[20][15] , \sa_ctrl[20].f.spare[10] );
tran (\sa_ctrl[20][16] , \sa_ctrl[20].r.part0[16] );
tran (\sa_ctrl[20][16] , \sa_ctrl[20].f.spare[11] );
tran (\sa_ctrl[20][17] , \sa_ctrl[20].r.part0[17] );
tran (\sa_ctrl[20][17] , \sa_ctrl[20].f.spare[12] );
tran (\sa_ctrl[20][18] , \sa_ctrl[20].r.part0[18] );
tran (\sa_ctrl[20][18] , \sa_ctrl[20].f.spare[13] );
tran (\sa_ctrl[20][19] , \sa_ctrl[20].r.part0[19] );
tran (\sa_ctrl[20][19] , \sa_ctrl[20].f.spare[14] );
tran (\sa_ctrl[20][20] , \sa_ctrl[20].r.part0[20] );
tran (\sa_ctrl[20][20] , \sa_ctrl[20].f.spare[15] );
tran (\sa_ctrl[20][21] , \sa_ctrl[20].r.part0[21] );
tran (\sa_ctrl[20][21] , \sa_ctrl[20].f.spare[16] );
tran (\sa_ctrl[20][22] , \sa_ctrl[20].r.part0[22] );
tran (\sa_ctrl[20][22] , \sa_ctrl[20].f.spare[17] );
tran (\sa_ctrl[20][23] , \sa_ctrl[20].r.part0[23] );
tran (\sa_ctrl[20][23] , \sa_ctrl[20].f.spare[18] );
tran (\sa_ctrl[20][24] , \sa_ctrl[20].r.part0[24] );
tran (\sa_ctrl[20][24] , \sa_ctrl[20].f.spare[19] );
tran (\sa_ctrl[20][25] , \sa_ctrl[20].r.part0[25] );
tran (\sa_ctrl[20][25] , \sa_ctrl[20].f.spare[20] );
tran (\sa_ctrl[20][26] , \sa_ctrl[20].r.part0[26] );
tran (\sa_ctrl[20][26] , \sa_ctrl[20].f.spare[21] );
tran (\sa_ctrl[20][27] , \sa_ctrl[20].r.part0[27] );
tran (\sa_ctrl[20][27] , \sa_ctrl[20].f.spare[22] );
tran (\sa_ctrl[20][28] , \sa_ctrl[20].r.part0[28] );
tran (\sa_ctrl[20][28] , \sa_ctrl[20].f.spare[23] );
tran (\sa_ctrl[20][29] , \sa_ctrl[20].r.part0[29] );
tran (\sa_ctrl[20][29] , \sa_ctrl[20].f.spare[24] );
tran (\sa_ctrl[20][30] , \sa_ctrl[20].r.part0[30] );
tran (\sa_ctrl[20][30] , \sa_ctrl[20].f.spare[25] );
tran (\sa_ctrl[20][31] , \sa_ctrl[20].r.part0[31] );
tran (\sa_ctrl[20][31] , \sa_ctrl[20].f.spare[26] );
tran (\sa_ctrl[21][0] , \sa_ctrl[21].r.part0[0] );
tran (\sa_ctrl[21][0] , \sa_ctrl[21].f.sa_event_sel[0] );
tran (\sa_ctrl[21][1] , \sa_ctrl[21].r.part0[1] );
tran (\sa_ctrl[21][1] , \sa_ctrl[21].f.sa_event_sel[1] );
tran (\sa_ctrl[21][2] , \sa_ctrl[21].r.part0[2] );
tran (\sa_ctrl[21][2] , \sa_ctrl[21].f.sa_event_sel[2] );
tran (\sa_ctrl[21][3] , \sa_ctrl[21].r.part0[3] );
tran (\sa_ctrl[21][3] , \sa_ctrl[21].f.sa_event_sel[3] );
tran (\sa_ctrl[21][4] , \sa_ctrl[21].r.part0[4] );
tran (\sa_ctrl[21][4] , \sa_ctrl[21].f.sa_event_sel[4] );
tran (\sa_ctrl[21][5] , \sa_ctrl[21].r.part0[5] );
tran (\sa_ctrl[21][5] , \sa_ctrl[21].f.spare[0] );
tran (\sa_ctrl[21][6] , \sa_ctrl[21].r.part0[6] );
tran (\sa_ctrl[21][6] , \sa_ctrl[21].f.spare[1] );
tran (\sa_ctrl[21][7] , \sa_ctrl[21].r.part0[7] );
tran (\sa_ctrl[21][7] , \sa_ctrl[21].f.spare[2] );
tran (\sa_ctrl[21][8] , \sa_ctrl[21].r.part0[8] );
tran (\sa_ctrl[21][8] , \sa_ctrl[21].f.spare[3] );
tran (\sa_ctrl[21][9] , \sa_ctrl[21].r.part0[9] );
tran (\sa_ctrl[21][9] , \sa_ctrl[21].f.spare[4] );
tran (\sa_ctrl[21][10] , \sa_ctrl[21].r.part0[10] );
tran (\sa_ctrl[21][10] , \sa_ctrl[21].f.spare[5] );
tran (\sa_ctrl[21][11] , \sa_ctrl[21].r.part0[11] );
tran (\sa_ctrl[21][11] , \sa_ctrl[21].f.spare[6] );
tran (\sa_ctrl[21][12] , \sa_ctrl[21].r.part0[12] );
tran (\sa_ctrl[21][12] , \sa_ctrl[21].f.spare[7] );
tran (\sa_ctrl[21][13] , \sa_ctrl[21].r.part0[13] );
tran (\sa_ctrl[21][13] , \sa_ctrl[21].f.spare[8] );
tran (\sa_ctrl[21][14] , \sa_ctrl[21].r.part0[14] );
tran (\sa_ctrl[21][14] , \sa_ctrl[21].f.spare[9] );
tran (\sa_ctrl[21][15] , \sa_ctrl[21].r.part0[15] );
tran (\sa_ctrl[21][15] , \sa_ctrl[21].f.spare[10] );
tran (\sa_ctrl[21][16] , \sa_ctrl[21].r.part0[16] );
tran (\sa_ctrl[21][16] , \sa_ctrl[21].f.spare[11] );
tran (\sa_ctrl[21][17] , \sa_ctrl[21].r.part0[17] );
tran (\sa_ctrl[21][17] , \sa_ctrl[21].f.spare[12] );
tran (\sa_ctrl[21][18] , \sa_ctrl[21].r.part0[18] );
tran (\sa_ctrl[21][18] , \sa_ctrl[21].f.spare[13] );
tran (\sa_ctrl[21][19] , \sa_ctrl[21].r.part0[19] );
tran (\sa_ctrl[21][19] , \sa_ctrl[21].f.spare[14] );
tran (\sa_ctrl[21][20] , \sa_ctrl[21].r.part0[20] );
tran (\sa_ctrl[21][20] , \sa_ctrl[21].f.spare[15] );
tran (\sa_ctrl[21][21] , \sa_ctrl[21].r.part0[21] );
tran (\sa_ctrl[21][21] , \sa_ctrl[21].f.spare[16] );
tran (\sa_ctrl[21][22] , \sa_ctrl[21].r.part0[22] );
tran (\sa_ctrl[21][22] , \sa_ctrl[21].f.spare[17] );
tran (\sa_ctrl[21][23] , \sa_ctrl[21].r.part0[23] );
tran (\sa_ctrl[21][23] , \sa_ctrl[21].f.spare[18] );
tran (\sa_ctrl[21][24] , \sa_ctrl[21].r.part0[24] );
tran (\sa_ctrl[21][24] , \sa_ctrl[21].f.spare[19] );
tran (\sa_ctrl[21][25] , \sa_ctrl[21].r.part0[25] );
tran (\sa_ctrl[21][25] , \sa_ctrl[21].f.spare[20] );
tran (\sa_ctrl[21][26] , \sa_ctrl[21].r.part0[26] );
tran (\sa_ctrl[21][26] , \sa_ctrl[21].f.spare[21] );
tran (\sa_ctrl[21][27] , \sa_ctrl[21].r.part0[27] );
tran (\sa_ctrl[21][27] , \sa_ctrl[21].f.spare[22] );
tran (\sa_ctrl[21][28] , \sa_ctrl[21].r.part0[28] );
tran (\sa_ctrl[21][28] , \sa_ctrl[21].f.spare[23] );
tran (\sa_ctrl[21][29] , \sa_ctrl[21].r.part0[29] );
tran (\sa_ctrl[21][29] , \sa_ctrl[21].f.spare[24] );
tran (\sa_ctrl[21][30] , \sa_ctrl[21].r.part0[30] );
tran (\sa_ctrl[21][30] , \sa_ctrl[21].f.spare[25] );
tran (\sa_ctrl[21][31] , \sa_ctrl[21].r.part0[31] );
tran (\sa_ctrl[21][31] , \sa_ctrl[21].f.spare[26] );
tran (\sa_ctrl[22][0] , \sa_ctrl[22].r.part0[0] );
tran (\sa_ctrl[22][0] , \sa_ctrl[22].f.sa_event_sel[0] );
tran (\sa_ctrl[22][1] , \sa_ctrl[22].r.part0[1] );
tran (\sa_ctrl[22][1] , \sa_ctrl[22].f.sa_event_sel[1] );
tran (\sa_ctrl[22][2] , \sa_ctrl[22].r.part0[2] );
tran (\sa_ctrl[22][2] , \sa_ctrl[22].f.sa_event_sel[2] );
tran (\sa_ctrl[22][3] , \sa_ctrl[22].r.part0[3] );
tran (\sa_ctrl[22][3] , \sa_ctrl[22].f.sa_event_sel[3] );
tran (\sa_ctrl[22][4] , \sa_ctrl[22].r.part0[4] );
tran (\sa_ctrl[22][4] , \sa_ctrl[22].f.sa_event_sel[4] );
tran (\sa_ctrl[22][5] , \sa_ctrl[22].r.part0[5] );
tran (\sa_ctrl[22][5] , \sa_ctrl[22].f.spare[0] );
tran (\sa_ctrl[22][6] , \sa_ctrl[22].r.part0[6] );
tran (\sa_ctrl[22][6] , \sa_ctrl[22].f.spare[1] );
tran (\sa_ctrl[22][7] , \sa_ctrl[22].r.part0[7] );
tran (\sa_ctrl[22][7] , \sa_ctrl[22].f.spare[2] );
tran (\sa_ctrl[22][8] , \sa_ctrl[22].r.part0[8] );
tran (\sa_ctrl[22][8] , \sa_ctrl[22].f.spare[3] );
tran (\sa_ctrl[22][9] , \sa_ctrl[22].r.part0[9] );
tran (\sa_ctrl[22][9] , \sa_ctrl[22].f.spare[4] );
tran (\sa_ctrl[22][10] , \sa_ctrl[22].r.part0[10] );
tran (\sa_ctrl[22][10] , \sa_ctrl[22].f.spare[5] );
tran (\sa_ctrl[22][11] , \sa_ctrl[22].r.part0[11] );
tran (\sa_ctrl[22][11] , \sa_ctrl[22].f.spare[6] );
tran (\sa_ctrl[22][12] , \sa_ctrl[22].r.part0[12] );
tran (\sa_ctrl[22][12] , \sa_ctrl[22].f.spare[7] );
tran (\sa_ctrl[22][13] , \sa_ctrl[22].r.part0[13] );
tran (\sa_ctrl[22][13] , \sa_ctrl[22].f.spare[8] );
tran (\sa_ctrl[22][14] , \sa_ctrl[22].r.part0[14] );
tran (\sa_ctrl[22][14] , \sa_ctrl[22].f.spare[9] );
tran (\sa_ctrl[22][15] , \sa_ctrl[22].r.part0[15] );
tran (\sa_ctrl[22][15] , \sa_ctrl[22].f.spare[10] );
tran (\sa_ctrl[22][16] , \sa_ctrl[22].r.part0[16] );
tran (\sa_ctrl[22][16] , \sa_ctrl[22].f.spare[11] );
tran (\sa_ctrl[22][17] , \sa_ctrl[22].r.part0[17] );
tran (\sa_ctrl[22][17] , \sa_ctrl[22].f.spare[12] );
tran (\sa_ctrl[22][18] , \sa_ctrl[22].r.part0[18] );
tran (\sa_ctrl[22][18] , \sa_ctrl[22].f.spare[13] );
tran (\sa_ctrl[22][19] , \sa_ctrl[22].r.part0[19] );
tran (\sa_ctrl[22][19] , \sa_ctrl[22].f.spare[14] );
tran (\sa_ctrl[22][20] , \sa_ctrl[22].r.part0[20] );
tran (\sa_ctrl[22][20] , \sa_ctrl[22].f.spare[15] );
tran (\sa_ctrl[22][21] , \sa_ctrl[22].r.part0[21] );
tran (\sa_ctrl[22][21] , \sa_ctrl[22].f.spare[16] );
tran (\sa_ctrl[22][22] , \sa_ctrl[22].r.part0[22] );
tran (\sa_ctrl[22][22] , \sa_ctrl[22].f.spare[17] );
tran (\sa_ctrl[22][23] , \sa_ctrl[22].r.part0[23] );
tran (\sa_ctrl[22][23] , \sa_ctrl[22].f.spare[18] );
tran (\sa_ctrl[22][24] , \sa_ctrl[22].r.part0[24] );
tran (\sa_ctrl[22][24] , \sa_ctrl[22].f.spare[19] );
tran (\sa_ctrl[22][25] , \sa_ctrl[22].r.part0[25] );
tran (\sa_ctrl[22][25] , \sa_ctrl[22].f.spare[20] );
tran (\sa_ctrl[22][26] , \sa_ctrl[22].r.part0[26] );
tran (\sa_ctrl[22][26] , \sa_ctrl[22].f.spare[21] );
tran (\sa_ctrl[22][27] , \sa_ctrl[22].r.part0[27] );
tran (\sa_ctrl[22][27] , \sa_ctrl[22].f.spare[22] );
tran (\sa_ctrl[22][28] , \sa_ctrl[22].r.part0[28] );
tran (\sa_ctrl[22][28] , \sa_ctrl[22].f.spare[23] );
tran (\sa_ctrl[22][29] , \sa_ctrl[22].r.part0[29] );
tran (\sa_ctrl[22][29] , \sa_ctrl[22].f.spare[24] );
tran (\sa_ctrl[22][30] , \sa_ctrl[22].r.part0[30] );
tran (\sa_ctrl[22][30] , \sa_ctrl[22].f.spare[25] );
tran (\sa_ctrl[22][31] , \sa_ctrl[22].r.part0[31] );
tran (\sa_ctrl[22][31] , \sa_ctrl[22].f.spare[26] );
tran (\sa_ctrl[23][0] , \sa_ctrl[23].r.part0[0] );
tran (\sa_ctrl[23][0] , \sa_ctrl[23].f.sa_event_sel[0] );
tran (\sa_ctrl[23][1] , \sa_ctrl[23].r.part0[1] );
tran (\sa_ctrl[23][1] , \sa_ctrl[23].f.sa_event_sel[1] );
tran (\sa_ctrl[23][2] , \sa_ctrl[23].r.part0[2] );
tran (\sa_ctrl[23][2] , \sa_ctrl[23].f.sa_event_sel[2] );
tran (\sa_ctrl[23][3] , \sa_ctrl[23].r.part0[3] );
tran (\sa_ctrl[23][3] , \sa_ctrl[23].f.sa_event_sel[3] );
tran (\sa_ctrl[23][4] , \sa_ctrl[23].r.part0[4] );
tran (\sa_ctrl[23][4] , \sa_ctrl[23].f.sa_event_sel[4] );
tran (\sa_ctrl[23][5] , \sa_ctrl[23].r.part0[5] );
tran (\sa_ctrl[23][5] , \sa_ctrl[23].f.spare[0] );
tran (\sa_ctrl[23][6] , \sa_ctrl[23].r.part0[6] );
tran (\sa_ctrl[23][6] , \sa_ctrl[23].f.spare[1] );
tran (\sa_ctrl[23][7] , \sa_ctrl[23].r.part0[7] );
tran (\sa_ctrl[23][7] , \sa_ctrl[23].f.spare[2] );
tran (\sa_ctrl[23][8] , \sa_ctrl[23].r.part0[8] );
tran (\sa_ctrl[23][8] , \sa_ctrl[23].f.spare[3] );
tran (\sa_ctrl[23][9] , \sa_ctrl[23].r.part0[9] );
tran (\sa_ctrl[23][9] , \sa_ctrl[23].f.spare[4] );
tran (\sa_ctrl[23][10] , \sa_ctrl[23].r.part0[10] );
tran (\sa_ctrl[23][10] , \sa_ctrl[23].f.spare[5] );
tran (\sa_ctrl[23][11] , \sa_ctrl[23].r.part0[11] );
tran (\sa_ctrl[23][11] , \sa_ctrl[23].f.spare[6] );
tran (\sa_ctrl[23][12] , \sa_ctrl[23].r.part0[12] );
tran (\sa_ctrl[23][12] , \sa_ctrl[23].f.spare[7] );
tran (\sa_ctrl[23][13] , \sa_ctrl[23].r.part0[13] );
tran (\sa_ctrl[23][13] , \sa_ctrl[23].f.spare[8] );
tran (\sa_ctrl[23][14] , \sa_ctrl[23].r.part0[14] );
tran (\sa_ctrl[23][14] , \sa_ctrl[23].f.spare[9] );
tran (\sa_ctrl[23][15] , \sa_ctrl[23].r.part0[15] );
tran (\sa_ctrl[23][15] , \sa_ctrl[23].f.spare[10] );
tran (\sa_ctrl[23][16] , \sa_ctrl[23].r.part0[16] );
tran (\sa_ctrl[23][16] , \sa_ctrl[23].f.spare[11] );
tran (\sa_ctrl[23][17] , \sa_ctrl[23].r.part0[17] );
tran (\sa_ctrl[23][17] , \sa_ctrl[23].f.spare[12] );
tran (\sa_ctrl[23][18] , \sa_ctrl[23].r.part0[18] );
tran (\sa_ctrl[23][18] , \sa_ctrl[23].f.spare[13] );
tran (\sa_ctrl[23][19] , \sa_ctrl[23].r.part0[19] );
tran (\sa_ctrl[23][19] , \sa_ctrl[23].f.spare[14] );
tran (\sa_ctrl[23][20] , \sa_ctrl[23].r.part0[20] );
tran (\sa_ctrl[23][20] , \sa_ctrl[23].f.spare[15] );
tran (\sa_ctrl[23][21] , \sa_ctrl[23].r.part0[21] );
tran (\sa_ctrl[23][21] , \sa_ctrl[23].f.spare[16] );
tran (\sa_ctrl[23][22] , \sa_ctrl[23].r.part0[22] );
tran (\sa_ctrl[23][22] , \sa_ctrl[23].f.spare[17] );
tran (\sa_ctrl[23][23] , \sa_ctrl[23].r.part0[23] );
tran (\sa_ctrl[23][23] , \sa_ctrl[23].f.spare[18] );
tran (\sa_ctrl[23][24] , \sa_ctrl[23].r.part0[24] );
tran (\sa_ctrl[23][24] , \sa_ctrl[23].f.spare[19] );
tran (\sa_ctrl[23][25] , \sa_ctrl[23].r.part0[25] );
tran (\sa_ctrl[23][25] , \sa_ctrl[23].f.spare[20] );
tran (\sa_ctrl[23][26] , \sa_ctrl[23].r.part0[26] );
tran (\sa_ctrl[23][26] , \sa_ctrl[23].f.spare[21] );
tran (\sa_ctrl[23][27] , \sa_ctrl[23].r.part0[27] );
tran (\sa_ctrl[23][27] , \sa_ctrl[23].f.spare[22] );
tran (\sa_ctrl[23][28] , \sa_ctrl[23].r.part0[28] );
tran (\sa_ctrl[23][28] , \sa_ctrl[23].f.spare[23] );
tran (\sa_ctrl[23][29] , \sa_ctrl[23].r.part0[29] );
tran (\sa_ctrl[23][29] , \sa_ctrl[23].f.spare[24] );
tran (\sa_ctrl[23][30] , \sa_ctrl[23].r.part0[30] );
tran (\sa_ctrl[23][30] , \sa_ctrl[23].f.spare[25] );
tran (\sa_ctrl[23][31] , \sa_ctrl[23].r.part0[31] );
tran (\sa_ctrl[23][31] , \sa_ctrl[23].f.spare[26] );
tran (\sa_ctrl[24][0] , \sa_ctrl[24].r.part0[0] );
tran (\sa_ctrl[24][0] , \sa_ctrl[24].f.sa_event_sel[0] );
tran (\sa_ctrl[24][1] , \sa_ctrl[24].r.part0[1] );
tran (\sa_ctrl[24][1] , \sa_ctrl[24].f.sa_event_sel[1] );
tran (\sa_ctrl[24][2] , \sa_ctrl[24].r.part0[2] );
tran (\sa_ctrl[24][2] , \sa_ctrl[24].f.sa_event_sel[2] );
tran (\sa_ctrl[24][3] , \sa_ctrl[24].r.part0[3] );
tran (\sa_ctrl[24][3] , \sa_ctrl[24].f.sa_event_sel[3] );
tran (\sa_ctrl[24][4] , \sa_ctrl[24].r.part0[4] );
tran (\sa_ctrl[24][4] , \sa_ctrl[24].f.sa_event_sel[4] );
tran (\sa_ctrl[24][5] , \sa_ctrl[24].r.part0[5] );
tran (\sa_ctrl[24][5] , \sa_ctrl[24].f.spare[0] );
tran (\sa_ctrl[24][6] , \sa_ctrl[24].r.part0[6] );
tran (\sa_ctrl[24][6] , \sa_ctrl[24].f.spare[1] );
tran (\sa_ctrl[24][7] , \sa_ctrl[24].r.part0[7] );
tran (\sa_ctrl[24][7] , \sa_ctrl[24].f.spare[2] );
tran (\sa_ctrl[24][8] , \sa_ctrl[24].r.part0[8] );
tran (\sa_ctrl[24][8] , \sa_ctrl[24].f.spare[3] );
tran (\sa_ctrl[24][9] , \sa_ctrl[24].r.part0[9] );
tran (\sa_ctrl[24][9] , \sa_ctrl[24].f.spare[4] );
tran (\sa_ctrl[24][10] , \sa_ctrl[24].r.part0[10] );
tran (\sa_ctrl[24][10] , \sa_ctrl[24].f.spare[5] );
tran (\sa_ctrl[24][11] , \sa_ctrl[24].r.part0[11] );
tran (\sa_ctrl[24][11] , \sa_ctrl[24].f.spare[6] );
tran (\sa_ctrl[24][12] , \sa_ctrl[24].r.part0[12] );
tran (\sa_ctrl[24][12] , \sa_ctrl[24].f.spare[7] );
tran (\sa_ctrl[24][13] , \sa_ctrl[24].r.part0[13] );
tran (\sa_ctrl[24][13] , \sa_ctrl[24].f.spare[8] );
tran (\sa_ctrl[24][14] , \sa_ctrl[24].r.part0[14] );
tran (\sa_ctrl[24][14] , \sa_ctrl[24].f.spare[9] );
tran (\sa_ctrl[24][15] , \sa_ctrl[24].r.part0[15] );
tran (\sa_ctrl[24][15] , \sa_ctrl[24].f.spare[10] );
tran (\sa_ctrl[24][16] , \sa_ctrl[24].r.part0[16] );
tran (\sa_ctrl[24][16] , \sa_ctrl[24].f.spare[11] );
tran (\sa_ctrl[24][17] , \sa_ctrl[24].r.part0[17] );
tran (\sa_ctrl[24][17] , \sa_ctrl[24].f.spare[12] );
tran (\sa_ctrl[24][18] , \sa_ctrl[24].r.part0[18] );
tran (\sa_ctrl[24][18] , \sa_ctrl[24].f.spare[13] );
tran (\sa_ctrl[24][19] , \sa_ctrl[24].r.part0[19] );
tran (\sa_ctrl[24][19] , \sa_ctrl[24].f.spare[14] );
tran (\sa_ctrl[24][20] , \sa_ctrl[24].r.part0[20] );
tran (\sa_ctrl[24][20] , \sa_ctrl[24].f.spare[15] );
tran (\sa_ctrl[24][21] , \sa_ctrl[24].r.part0[21] );
tran (\sa_ctrl[24][21] , \sa_ctrl[24].f.spare[16] );
tran (\sa_ctrl[24][22] , \sa_ctrl[24].r.part0[22] );
tran (\sa_ctrl[24][22] , \sa_ctrl[24].f.spare[17] );
tran (\sa_ctrl[24][23] , \sa_ctrl[24].r.part0[23] );
tran (\sa_ctrl[24][23] , \sa_ctrl[24].f.spare[18] );
tran (\sa_ctrl[24][24] , \sa_ctrl[24].r.part0[24] );
tran (\sa_ctrl[24][24] , \sa_ctrl[24].f.spare[19] );
tran (\sa_ctrl[24][25] , \sa_ctrl[24].r.part0[25] );
tran (\sa_ctrl[24][25] , \sa_ctrl[24].f.spare[20] );
tran (\sa_ctrl[24][26] , \sa_ctrl[24].r.part0[26] );
tran (\sa_ctrl[24][26] , \sa_ctrl[24].f.spare[21] );
tran (\sa_ctrl[24][27] , \sa_ctrl[24].r.part0[27] );
tran (\sa_ctrl[24][27] , \sa_ctrl[24].f.spare[22] );
tran (\sa_ctrl[24][28] , \sa_ctrl[24].r.part0[28] );
tran (\sa_ctrl[24][28] , \sa_ctrl[24].f.spare[23] );
tran (\sa_ctrl[24][29] , \sa_ctrl[24].r.part0[29] );
tran (\sa_ctrl[24][29] , \sa_ctrl[24].f.spare[24] );
tran (\sa_ctrl[24][30] , \sa_ctrl[24].r.part0[30] );
tran (\sa_ctrl[24][30] , \sa_ctrl[24].f.spare[25] );
tran (\sa_ctrl[24][31] , \sa_ctrl[24].r.part0[31] );
tran (\sa_ctrl[24][31] , \sa_ctrl[24].f.spare[26] );
tran (\sa_ctrl[25][0] , \sa_ctrl[25].r.part0[0] );
tran (\sa_ctrl[25][0] , \sa_ctrl[25].f.sa_event_sel[0] );
tran (\sa_ctrl[25][1] , \sa_ctrl[25].r.part0[1] );
tran (\sa_ctrl[25][1] , \sa_ctrl[25].f.sa_event_sel[1] );
tran (\sa_ctrl[25][2] , \sa_ctrl[25].r.part0[2] );
tran (\sa_ctrl[25][2] , \sa_ctrl[25].f.sa_event_sel[2] );
tran (\sa_ctrl[25][3] , \sa_ctrl[25].r.part0[3] );
tran (\sa_ctrl[25][3] , \sa_ctrl[25].f.sa_event_sel[3] );
tran (\sa_ctrl[25][4] , \sa_ctrl[25].r.part0[4] );
tran (\sa_ctrl[25][4] , \sa_ctrl[25].f.sa_event_sel[4] );
tran (\sa_ctrl[25][5] , \sa_ctrl[25].r.part0[5] );
tran (\sa_ctrl[25][5] , \sa_ctrl[25].f.spare[0] );
tran (\sa_ctrl[25][6] , \sa_ctrl[25].r.part0[6] );
tran (\sa_ctrl[25][6] , \sa_ctrl[25].f.spare[1] );
tran (\sa_ctrl[25][7] , \sa_ctrl[25].r.part0[7] );
tran (\sa_ctrl[25][7] , \sa_ctrl[25].f.spare[2] );
tran (\sa_ctrl[25][8] , \sa_ctrl[25].r.part0[8] );
tran (\sa_ctrl[25][8] , \sa_ctrl[25].f.spare[3] );
tran (\sa_ctrl[25][9] , \sa_ctrl[25].r.part0[9] );
tran (\sa_ctrl[25][9] , \sa_ctrl[25].f.spare[4] );
tran (\sa_ctrl[25][10] , \sa_ctrl[25].r.part0[10] );
tran (\sa_ctrl[25][10] , \sa_ctrl[25].f.spare[5] );
tran (\sa_ctrl[25][11] , \sa_ctrl[25].r.part0[11] );
tran (\sa_ctrl[25][11] , \sa_ctrl[25].f.spare[6] );
tran (\sa_ctrl[25][12] , \sa_ctrl[25].r.part0[12] );
tran (\sa_ctrl[25][12] , \sa_ctrl[25].f.spare[7] );
tran (\sa_ctrl[25][13] , \sa_ctrl[25].r.part0[13] );
tran (\sa_ctrl[25][13] , \sa_ctrl[25].f.spare[8] );
tran (\sa_ctrl[25][14] , \sa_ctrl[25].r.part0[14] );
tran (\sa_ctrl[25][14] , \sa_ctrl[25].f.spare[9] );
tran (\sa_ctrl[25][15] , \sa_ctrl[25].r.part0[15] );
tran (\sa_ctrl[25][15] , \sa_ctrl[25].f.spare[10] );
tran (\sa_ctrl[25][16] , \sa_ctrl[25].r.part0[16] );
tran (\sa_ctrl[25][16] , \sa_ctrl[25].f.spare[11] );
tran (\sa_ctrl[25][17] , \sa_ctrl[25].r.part0[17] );
tran (\sa_ctrl[25][17] , \sa_ctrl[25].f.spare[12] );
tran (\sa_ctrl[25][18] , \sa_ctrl[25].r.part0[18] );
tran (\sa_ctrl[25][18] , \sa_ctrl[25].f.spare[13] );
tran (\sa_ctrl[25][19] , \sa_ctrl[25].r.part0[19] );
tran (\sa_ctrl[25][19] , \sa_ctrl[25].f.spare[14] );
tran (\sa_ctrl[25][20] , \sa_ctrl[25].r.part0[20] );
tran (\sa_ctrl[25][20] , \sa_ctrl[25].f.spare[15] );
tran (\sa_ctrl[25][21] , \sa_ctrl[25].r.part0[21] );
tran (\sa_ctrl[25][21] , \sa_ctrl[25].f.spare[16] );
tran (\sa_ctrl[25][22] , \sa_ctrl[25].r.part0[22] );
tran (\sa_ctrl[25][22] , \sa_ctrl[25].f.spare[17] );
tran (\sa_ctrl[25][23] , \sa_ctrl[25].r.part0[23] );
tran (\sa_ctrl[25][23] , \sa_ctrl[25].f.spare[18] );
tran (\sa_ctrl[25][24] , \sa_ctrl[25].r.part0[24] );
tran (\sa_ctrl[25][24] , \sa_ctrl[25].f.spare[19] );
tran (\sa_ctrl[25][25] , \sa_ctrl[25].r.part0[25] );
tran (\sa_ctrl[25][25] , \sa_ctrl[25].f.spare[20] );
tran (\sa_ctrl[25][26] , \sa_ctrl[25].r.part0[26] );
tran (\sa_ctrl[25][26] , \sa_ctrl[25].f.spare[21] );
tran (\sa_ctrl[25][27] , \sa_ctrl[25].r.part0[27] );
tran (\sa_ctrl[25][27] , \sa_ctrl[25].f.spare[22] );
tran (\sa_ctrl[25][28] , \sa_ctrl[25].r.part0[28] );
tran (\sa_ctrl[25][28] , \sa_ctrl[25].f.spare[23] );
tran (\sa_ctrl[25][29] , \sa_ctrl[25].r.part0[29] );
tran (\sa_ctrl[25][29] , \sa_ctrl[25].f.spare[24] );
tran (\sa_ctrl[25][30] , \sa_ctrl[25].r.part0[30] );
tran (\sa_ctrl[25][30] , \sa_ctrl[25].f.spare[25] );
tran (\sa_ctrl[25][31] , \sa_ctrl[25].r.part0[31] );
tran (\sa_ctrl[25][31] , \sa_ctrl[25].f.spare[26] );
tran (\sa_ctrl[26][0] , \sa_ctrl[26].r.part0[0] );
tran (\sa_ctrl[26][0] , \sa_ctrl[26].f.sa_event_sel[0] );
tran (\sa_ctrl[26][1] , \sa_ctrl[26].r.part0[1] );
tran (\sa_ctrl[26][1] , \sa_ctrl[26].f.sa_event_sel[1] );
tran (\sa_ctrl[26][2] , \sa_ctrl[26].r.part0[2] );
tran (\sa_ctrl[26][2] , \sa_ctrl[26].f.sa_event_sel[2] );
tran (\sa_ctrl[26][3] , \sa_ctrl[26].r.part0[3] );
tran (\sa_ctrl[26][3] , \sa_ctrl[26].f.sa_event_sel[3] );
tran (\sa_ctrl[26][4] , \sa_ctrl[26].r.part0[4] );
tran (\sa_ctrl[26][4] , \sa_ctrl[26].f.sa_event_sel[4] );
tran (\sa_ctrl[26][5] , \sa_ctrl[26].r.part0[5] );
tran (\sa_ctrl[26][5] , \sa_ctrl[26].f.spare[0] );
tran (\sa_ctrl[26][6] , \sa_ctrl[26].r.part0[6] );
tran (\sa_ctrl[26][6] , \sa_ctrl[26].f.spare[1] );
tran (\sa_ctrl[26][7] , \sa_ctrl[26].r.part0[7] );
tran (\sa_ctrl[26][7] , \sa_ctrl[26].f.spare[2] );
tran (\sa_ctrl[26][8] , \sa_ctrl[26].r.part0[8] );
tran (\sa_ctrl[26][8] , \sa_ctrl[26].f.spare[3] );
tran (\sa_ctrl[26][9] , \sa_ctrl[26].r.part0[9] );
tran (\sa_ctrl[26][9] , \sa_ctrl[26].f.spare[4] );
tran (\sa_ctrl[26][10] , \sa_ctrl[26].r.part0[10] );
tran (\sa_ctrl[26][10] , \sa_ctrl[26].f.spare[5] );
tran (\sa_ctrl[26][11] , \sa_ctrl[26].r.part0[11] );
tran (\sa_ctrl[26][11] , \sa_ctrl[26].f.spare[6] );
tran (\sa_ctrl[26][12] , \sa_ctrl[26].r.part0[12] );
tran (\sa_ctrl[26][12] , \sa_ctrl[26].f.spare[7] );
tran (\sa_ctrl[26][13] , \sa_ctrl[26].r.part0[13] );
tran (\sa_ctrl[26][13] , \sa_ctrl[26].f.spare[8] );
tran (\sa_ctrl[26][14] , \sa_ctrl[26].r.part0[14] );
tran (\sa_ctrl[26][14] , \sa_ctrl[26].f.spare[9] );
tran (\sa_ctrl[26][15] , \sa_ctrl[26].r.part0[15] );
tran (\sa_ctrl[26][15] , \sa_ctrl[26].f.spare[10] );
tran (\sa_ctrl[26][16] , \sa_ctrl[26].r.part0[16] );
tran (\sa_ctrl[26][16] , \sa_ctrl[26].f.spare[11] );
tran (\sa_ctrl[26][17] , \sa_ctrl[26].r.part0[17] );
tran (\sa_ctrl[26][17] , \sa_ctrl[26].f.spare[12] );
tran (\sa_ctrl[26][18] , \sa_ctrl[26].r.part0[18] );
tran (\sa_ctrl[26][18] , \sa_ctrl[26].f.spare[13] );
tran (\sa_ctrl[26][19] , \sa_ctrl[26].r.part0[19] );
tran (\sa_ctrl[26][19] , \sa_ctrl[26].f.spare[14] );
tran (\sa_ctrl[26][20] , \sa_ctrl[26].r.part0[20] );
tran (\sa_ctrl[26][20] , \sa_ctrl[26].f.spare[15] );
tran (\sa_ctrl[26][21] , \sa_ctrl[26].r.part0[21] );
tran (\sa_ctrl[26][21] , \sa_ctrl[26].f.spare[16] );
tran (\sa_ctrl[26][22] , \sa_ctrl[26].r.part0[22] );
tran (\sa_ctrl[26][22] , \sa_ctrl[26].f.spare[17] );
tran (\sa_ctrl[26][23] , \sa_ctrl[26].r.part0[23] );
tran (\sa_ctrl[26][23] , \sa_ctrl[26].f.spare[18] );
tran (\sa_ctrl[26][24] , \sa_ctrl[26].r.part0[24] );
tran (\sa_ctrl[26][24] , \sa_ctrl[26].f.spare[19] );
tran (\sa_ctrl[26][25] , \sa_ctrl[26].r.part0[25] );
tran (\sa_ctrl[26][25] , \sa_ctrl[26].f.spare[20] );
tran (\sa_ctrl[26][26] , \sa_ctrl[26].r.part0[26] );
tran (\sa_ctrl[26][26] , \sa_ctrl[26].f.spare[21] );
tran (\sa_ctrl[26][27] , \sa_ctrl[26].r.part0[27] );
tran (\sa_ctrl[26][27] , \sa_ctrl[26].f.spare[22] );
tran (\sa_ctrl[26][28] , \sa_ctrl[26].r.part0[28] );
tran (\sa_ctrl[26][28] , \sa_ctrl[26].f.spare[23] );
tran (\sa_ctrl[26][29] , \sa_ctrl[26].r.part0[29] );
tran (\sa_ctrl[26][29] , \sa_ctrl[26].f.spare[24] );
tran (\sa_ctrl[26][30] , \sa_ctrl[26].r.part0[30] );
tran (\sa_ctrl[26][30] , \sa_ctrl[26].f.spare[25] );
tran (\sa_ctrl[26][31] , \sa_ctrl[26].r.part0[31] );
tran (\sa_ctrl[26][31] , \sa_ctrl[26].f.spare[26] );
tran (\sa_ctrl[27][0] , \sa_ctrl[27].r.part0[0] );
tran (\sa_ctrl[27][0] , \sa_ctrl[27].f.sa_event_sel[0] );
tran (\sa_ctrl[27][1] , \sa_ctrl[27].r.part0[1] );
tran (\sa_ctrl[27][1] , \sa_ctrl[27].f.sa_event_sel[1] );
tran (\sa_ctrl[27][2] , \sa_ctrl[27].r.part0[2] );
tran (\sa_ctrl[27][2] , \sa_ctrl[27].f.sa_event_sel[2] );
tran (\sa_ctrl[27][3] , \sa_ctrl[27].r.part0[3] );
tran (\sa_ctrl[27][3] , \sa_ctrl[27].f.sa_event_sel[3] );
tran (\sa_ctrl[27][4] , \sa_ctrl[27].r.part0[4] );
tran (\sa_ctrl[27][4] , \sa_ctrl[27].f.sa_event_sel[4] );
tran (\sa_ctrl[27][5] , \sa_ctrl[27].r.part0[5] );
tran (\sa_ctrl[27][5] , \sa_ctrl[27].f.spare[0] );
tran (\sa_ctrl[27][6] , \sa_ctrl[27].r.part0[6] );
tran (\sa_ctrl[27][6] , \sa_ctrl[27].f.spare[1] );
tran (\sa_ctrl[27][7] , \sa_ctrl[27].r.part0[7] );
tran (\sa_ctrl[27][7] , \sa_ctrl[27].f.spare[2] );
tran (\sa_ctrl[27][8] , \sa_ctrl[27].r.part0[8] );
tran (\sa_ctrl[27][8] , \sa_ctrl[27].f.spare[3] );
tran (\sa_ctrl[27][9] , \sa_ctrl[27].r.part0[9] );
tran (\sa_ctrl[27][9] , \sa_ctrl[27].f.spare[4] );
tran (\sa_ctrl[27][10] , \sa_ctrl[27].r.part0[10] );
tran (\sa_ctrl[27][10] , \sa_ctrl[27].f.spare[5] );
tran (\sa_ctrl[27][11] , \sa_ctrl[27].r.part0[11] );
tran (\sa_ctrl[27][11] , \sa_ctrl[27].f.spare[6] );
tran (\sa_ctrl[27][12] , \sa_ctrl[27].r.part0[12] );
tran (\sa_ctrl[27][12] , \sa_ctrl[27].f.spare[7] );
tran (\sa_ctrl[27][13] , \sa_ctrl[27].r.part0[13] );
tran (\sa_ctrl[27][13] , \sa_ctrl[27].f.spare[8] );
tran (\sa_ctrl[27][14] , \sa_ctrl[27].r.part0[14] );
tran (\sa_ctrl[27][14] , \sa_ctrl[27].f.spare[9] );
tran (\sa_ctrl[27][15] , \sa_ctrl[27].r.part0[15] );
tran (\sa_ctrl[27][15] , \sa_ctrl[27].f.spare[10] );
tran (\sa_ctrl[27][16] , \sa_ctrl[27].r.part0[16] );
tran (\sa_ctrl[27][16] , \sa_ctrl[27].f.spare[11] );
tran (\sa_ctrl[27][17] , \sa_ctrl[27].r.part0[17] );
tran (\sa_ctrl[27][17] , \sa_ctrl[27].f.spare[12] );
tran (\sa_ctrl[27][18] , \sa_ctrl[27].r.part0[18] );
tran (\sa_ctrl[27][18] , \sa_ctrl[27].f.spare[13] );
tran (\sa_ctrl[27][19] , \sa_ctrl[27].r.part0[19] );
tran (\sa_ctrl[27][19] , \sa_ctrl[27].f.spare[14] );
tran (\sa_ctrl[27][20] , \sa_ctrl[27].r.part0[20] );
tran (\sa_ctrl[27][20] , \sa_ctrl[27].f.spare[15] );
tran (\sa_ctrl[27][21] , \sa_ctrl[27].r.part0[21] );
tran (\sa_ctrl[27][21] , \sa_ctrl[27].f.spare[16] );
tran (\sa_ctrl[27][22] , \sa_ctrl[27].r.part0[22] );
tran (\sa_ctrl[27][22] , \sa_ctrl[27].f.spare[17] );
tran (\sa_ctrl[27][23] , \sa_ctrl[27].r.part0[23] );
tran (\sa_ctrl[27][23] , \sa_ctrl[27].f.spare[18] );
tran (\sa_ctrl[27][24] , \sa_ctrl[27].r.part0[24] );
tran (\sa_ctrl[27][24] , \sa_ctrl[27].f.spare[19] );
tran (\sa_ctrl[27][25] , \sa_ctrl[27].r.part0[25] );
tran (\sa_ctrl[27][25] , \sa_ctrl[27].f.spare[20] );
tran (\sa_ctrl[27][26] , \sa_ctrl[27].r.part0[26] );
tran (\sa_ctrl[27][26] , \sa_ctrl[27].f.spare[21] );
tran (\sa_ctrl[27][27] , \sa_ctrl[27].r.part0[27] );
tran (\sa_ctrl[27][27] , \sa_ctrl[27].f.spare[22] );
tran (\sa_ctrl[27][28] , \sa_ctrl[27].r.part0[28] );
tran (\sa_ctrl[27][28] , \sa_ctrl[27].f.spare[23] );
tran (\sa_ctrl[27][29] , \sa_ctrl[27].r.part0[29] );
tran (\sa_ctrl[27][29] , \sa_ctrl[27].f.spare[24] );
tran (\sa_ctrl[27][30] , \sa_ctrl[27].r.part0[30] );
tran (\sa_ctrl[27][30] , \sa_ctrl[27].f.spare[25] );
tran (\sa_ctrl[27][31] , \sa_ctrl[27].r.part0[31] );
tran (\sa_ctrl[27][31] , \sa_ctrl[27].f.spare[26] );
tran (\sa_ctrl[28][0] , \sa_ctrl[28].r.part0[0] );
tran (\sa_ctrl[28][0] , \sa_ctrl[28].f.sa_event_sel[0] );
tran (\sa_ctrl[28][1] , \sa_ctrl[28].r.part0[1] );
tran (\sa_ctrl[28][1] , \sa_ctrl[28].f.sa_event_sel[1] );
tran (\sa_ctrl[28][2] , \sa_ctrl[28].r.part0[2] );
tran (\sa_ctrl[28][2] , \sa_ctrl[28].f.sa_event_sel[2] );
tran (\sa_ctrl[28][3] , \sa_ctrl[28].r.part0[3] );
tran (\sa_ctrl[28][3] , \sa_ctrl[28].f.sa_event_sel[3] );
tran (\sa_ctrl[28][4] , \sa_ctrl[28].r.part0[4] );
tran (\sa_ctrl[28][4] , \sa_ctrl[28].f.sa_event_sel[4] );
tran (\sa_ctrl[28][5] , \sa_ctrl[28].r.part0[5] );
tran (\sa_ctrl[28][5] , \sa_ctrl[28].f.spare[0] );
tran (\sa_ctrl[28][6] , \sa_ctrl[28].r.part0[6] );
tran (\sa_ctrl[28][6] , \sa_ctrl[28].f.spare[1] );
tran (\sa_ctrl[28][7] , \sa_ctrl[28].r.part0[7] );
tran (\sa_ctrl[28][7] , \sa_ctrl[28].f.spare[2] );
tran (\sa_ctrl[28][8] , \sa_ctrl[28].r.part0[8] );
tran (\sa_ctrl[28][8] , \sa_ctrl[28].f.spare[3] );
tran (\sa_ctrl[28][9] , \sa_ctrl[28].r.part0[9] );
tran (\sa_ctrl[28][9] , \sa_ctrl[28].f.spare[4] );
tran (\sa_ctrl[28][10] , \sa_ctrl[28].r.part0[10] );
tran (\sa_ctrl[28][10] , \sa_ctrl[28].f.spare[5] );
tran (\sa_ctrl[28][11] , \sa_ctrl[28].r.part0[11] );
tran (\sa_ctrl[28][11] , \sa_ctrl[28].f.spare[6] );
tran (\sa_ctrl[28][12] , \sa_ctrl[28].r.part0[12] );
tran (\sa_ctrl[28][12] , \sa_ctrl[28].f.spare[7] );
tran (\sa_ctrl[28][13] , \sa_ctrl[28].r.part0[13] );
tran (\sa_ctrl[28][13] , \sa_ctrl[28].f.spare[8] );
tran (\sa_ctrl[28][14] , \sa_ctrl[28].r.part0[14] );
tran (\sa_ctrl[28][14] , \sa_ctrl[28].f.spare[9] );
tran (\sa_ctrl[28][15] , \sa_ctrl[28].r.part0[15] );
tran (\sa_ctrl[28][15] , \sa_ctrl[28].f.spare[10] );
tran (\sa_ctrl[28][16] , \sa_ctrl[28].r.part0[16] );
tran (\sa_ctrl[28][16] , \sa_ctrl[28].f.spare[11] );
tran (\sa_ctrl[28][17] , \sa_ctrl[28].r.part0[17] );
tran (\sa_ctrl[28][17] , \sa_ctrl[28].f.spare[12] );
tran (\sa_ctrl[28][18] , \sa_ctrl[28].r.part0[18] );
tran (\sa_ctrl[28][18] , \sa_ctrl[28].f.spare[13] );
tran (\sa_ctrl[28][19] , \sa_ctrl[28].r.part0[19] );
tran (\sa_ctrl[28][19] , \sa_ctrl[28].f.spare[14] );
tran (\sa_ctrl[28][20] , \sa_ctrl[28].r.part0[20] );
tran (\sa_ctrl[28][20] , \sa_ctrl[28].f.spare[15] );
tran (\sa_ctrl[28][21] , \sa_ctrl[28].r.part0[21] );
tran (\sa_ctrl[28][21] , \sa_ctrl[28].f.spare[16] );
tran (\sa_ctrl[28][22] , \sa_ctrl[28].r.part0[22] );
tran (\sa_ctrl[28][22] , \sa_ctrl[28].f.spare[17] );
tran (\sa_ctrl[28][23] , \sa_ctrl[28].r.part0[23] );
tran (\sa_ctrl[28][23] , \sa_ctrl[28].f.spare[18] );
tran (\sa_ctrl[28][24] , \sa_ctrl[28].r.part0[24] );
tran (\sa_ctrl[28][24] , \sa_ctrl[28].f.spare[19] );
tran (\sa_ctrl[28][25] , \sa_ctrl[28].r.part0[25] );
tran (\sa_ctrl[28][25] , \sa_ctrl[28].f.spare[20] );
tran (\sa_ctrl[28][26] , \sa_ctrl[28].r.part0[26] );
tran (\sa_ctrl[28][26] , \sa_ctrl[28].f.spare[21] );
tran (\sa_ctrl[28][27] , \sa_ctrl[28].r.part0[27] );
tran (\sa_ctrl[28][27] , \sa_ctrl[28].f.spare[22] );
tran (\sa_ctrl[28][28] , \sa_ctrl[28].r.part0[28] );
tran (\sa_ctrl[28][28] , \sa_ctrl[28].f.spare[23] );
tran (\sa_ctrl[28][29] , \sa_ctrl[28].r.part0[29] );
tran (\sa_ctrl[28][29] , \sa_ctrl[28].f.spare[24] );
tran (\sa_ctrl[28][30] , \sa_ctrl[28].r.part0[30] );
tran (\sa_ctrl[28][30] , \sa_ctrl[28].f.spare[25] );
tran (\sa_ctrl[28][31] , \sa_ctrl[28].r.part0[31] );
tran (\sa_ctrl[28][31] , \sa_ctrl[28].f.spare[26] );
tran (\sa_ctrl[29][0] , \sa_ctrl[29].r.part0[0] );
tran (\sa_ctrl[29][0] , \sa_ctrl[29].f.sa_event_sel[0] );
tran (\sa_ctrl[29][1] , \sa_ctrl[29].r.part0[1] );
tran (\sa_ctrl[29][1] , \sa_ctrl[29].f.sa_event_sel[1] );
tran (\sa_ctrl[29][2] , \sa_ctrl[29].r.part0[2] );
tran (\sa_ctrl[29][2] , \sa_ctrl[29].f.sa_event_sel[2] );
tran (\sa_ctrl[29][3] , \sa_ctrl[29].r.part0[3] );
tran (\sa_ctrl[29][3] , \sa_ctrl[29].f.sa_event_sel[3] );
tran (\sa_ctrl[29][4] , \sa_ctrl[29].r.part0[4] );
tran (\sa_ctrl[29][4] , \sa_ctrl[29].f.sa_event_sel[4] );
tran (\sa_ctrl[29][5] , \sa_ctrl[29].r.part0[5] );
tran (\sa_ctrl[29][5] , \sa_ctrl[29].f.spare[0] );
tran (\sa_ctrl[29][6] , \sa_ctrl[29].r.part0[6] );
tran (\sa_ctrl[29][6] , \sa_ctrl[29].f.spare[1] );
tran (\sa_ctrl[29][7] , \sa_ctrl[29].r.part0[7] );
tran (\sa_ctrl[29][7] , \sa_ctrl[29].f.spare[2] );
tran (\sa_ctrl[29][8] , \sa_ctrl[29].r.part0[8] );
tran (\sa_ctrl[29][8] , \sa_ctrl[29].f.spare[3] );
tran (\sa_ctrl[29][9] , \sa_ctrl[29].r.part0[9] );
tran (\sa_ctrl[29][9] , \sa_ctrl[29].f.spare[4] );
tran (\sa_ctrl[29][10] , \sa_ctrl[29].r.part0[10] );
tran (\sa_ctrl[29][10] , \sa_ctrl[29].f.spare[5] );
tran (\sa_ctrl[29][11] , \sa_ctrl[29].r.part0[11] );
tran (\sa_ctrl[29][11] , \sa_ctrl[29].f.spare[6] );
tran (\sa_ctrl[29][12] , \sa_ctrl[29].r.part0[12] );
tran (\sa_ctrl[29][12] , \sa_ctrl[29].f.spare[7] );
tran (\sa_ctrl[29][13] , \sa_ctrl[29].r.part0[13] );
tran (\sa_ctrl[29][13] , \sa_ctrl[29].f.spare[8] );
tran (\sa_ctrl[29][14] , \sa_ctrl[29].r.part0[14] );
tran (\sa_ctrl[29][14] , \sa_ctrl[29].f.spare[9] );
tran (\sa_ctrl[29][15] , \sa_ctrl[29].r.part0[15] );
tran (\sa_ctrl[29][15] , \sa_ctrl[29].f.spare[10] );
tran (\sa_ctrl[29][16] , \sa_ctrl[29].r.part0[16] );
tran (\sa_ctrl[29][16] , \sa_ctrl[29].f.spare[11] );
tran (\sa_ctrl[29][17] , \sa_ctrl[29].r.part0[17] );
tran (\sa_ctrl[29][17] , \sa_ctrl[29].f.spare[12] );
tran (\sa_ctrl[29][18] , \sa_ctrl[29].r.part0[18] );
tran (\sa_ctrl[29][18] , \sa_ctrl[29].f.spare[13] );
tran (\sa_ctrl[29][19] , \sa_ctrl[29].r.part0[19] );
tran (\sa_ctrl[29][19] , \sa_ctrl[29].f.spare[14] );
tran (\sa_ctrl[29][20] , \sa_ctrl[29].r.part0[20] );
tran (\sa_ctrl[29][20] , \sa_ctrl[29].f.spare[15] );
tran (\sa_ctrl[29][21] , \sa_ctrl[29].r.part0[21] );
tran (\sa_ctrl[29][21] , \sa_ctrl[29].f.spare[16] );
tran (\sa_ctrl[29][22] , \sa_ctrl[29].r.part0[22] );
tran (\sa_ctrl[29][22] , \sa_ctrl[29].f.spare[17] );
tran (\sa_ctrl[29][23] , \sa_ctrl[29].r.part0[23] );
tran (\sa_ctrl[29][23] , \sa_ctrl[29].f.spare[18] );
tran (\sa_ctrl[29][24] , \sa_ctrl[29].r.part0[24] );
tran (\sa_ctrl[29][24] , \sa_ctrl[29].f.spare[19] );
tran (\sa_ctrl[29][25] , \sa_ctrl[29].r.part0[25] );
tran (\sa_ctrl[29][25] , \sa_ctrl[29].f.spare[20] );
tran (\sa_ctrl[29][26] , \sa_ctrl[29].r.part0[26] );
tran (\sa_ctrl[29][26] , \sa_ctrl[29].f.spare[21] );
tran (\sa_ctrl[29][27] , \sa_ctrl[29].r.part0[27] );
tran (\sa_ctrl[29][27] , \sa_ctrl[29].f.spare[22] );
tran (\sa_ctrl[29][28] , \sa_ctrl[29].r.part0[28] );
tran (\sa_ctrl[29][28] , \sa_ctrl[29].f.spare[23] );
tran (\sa_ctrl[29][29] , \sa_ctrl[29].r.part0[29] );
tran (\sa_ctrl[29][29] , \sa_ctrl[29].f.spare[24] );
tran (\sa_ctrl[29][30] , \sa_ctrl[29].r.part0[30] );
tran (\sa_ctrl[29][30] , \sa_ctrl[29].f.spare[25] );
tran (\sa_ctrl[29][31] , \sa_ctrl[29].r.part0[31] );
tran (\sa_ctrl[29][31] , \sa_ctrl[29].f.spare[26] );
tran (\sa_ctrl[30][0] , \sa_ctrl[30].r.part0[0] );
tran (\sa_ctrl[30][0] , \sa_ctrl[30].f.sa_event_sel[0] );
tran (\sa_ctrl[30][1] , \sa_ctrl[30].r.part0[1] );
tran (\sa_ctrl[30][1] , \sa_ctrl[30].f.sa_event_sel[1] );
tran (\sa_ctrl[30][2] , \sa_ctrl[30].r.part0[2] );
tran (\sa_ctrl[30][2] , \sa_ctrl[30].f.sa_event_sel[2] );
tran (\sa_ctrl[30][3] , \sa_ctrl[30].r.part0[3] );
tran (\sa_ctrl[30][3] , \sa_ctrl[30].f.sa_event_sel[3] );
tran (\sa_ctrl[30][4] , \sa_ctrl[30].r.part0[4] );
tran (\sa_ctrl[30][4] , \sa_ctrl[30].f.sa_event_sel[4] );
tran (\sa_ctrl[30][5] , \sa_ctrl[30].r.part0[5] );
tran (\sa_ctrl[30][5] , \sa_ctrl[30].f.spare[0] );
tran (\sa_ctrl[30][6] , \sa_ctrl[30].r.part0[6] );
tran (\sa_ctrl[30][6] , \sa_ctrl[30].f.spare[1] );
tran (\sa_ctrl[30][7] , \sa_ctrl[30].r.part0[7] );
tran (\sa_ctrl[30][7] , \sa_ctrl[30].f.spare[2] );
tran (\sa_ctrl[30][8] , \sa_ctrl[30].r.part0[8] );
tran (\sa_ctrl[30][8] , \sa_ctrl[30].f.spare[3] );
tran (\sa_ctrl[30][9] , \sa_ctrl[30].r.part0[9] );
tran (\sa_ctrl[30][9] , \sa_ctrl[30].f.spare[4] );
tran (\sa_ctrl[30][10] , \sa_ctrl[30].r.part0[10] );
tran (\sa_ctrl[30][10] , \sa_ctrl[30].f.spare[5] );
tran (\sa_ctrl[30][11] , \sa_ctrl[30].r.part0[11] );
tran (\sa_ctrl[30][11] , \sa_ctrl[30].f.spare[6] );
tran (\sa_ctrl[30][12] , \sa_ctrl[30].r.part0[12] );
tran (\sa_ctrl[30][12] , \sa_ctrl[30].f.spare[7] );
tran (\sa_ctrl[30][13] , \sa_ctrl[30].r.part0[13] );
tran (\sa_ctrl[30][13] , \sa_ctrl[30].f.spare[8] );
tran (\sa_ctrl[30][14] , \sa_ctrl[30].r.part0[14] );
tran (\sa_ctrl[30][14] , \sa_ctrl[30].f.spare[9] );
tran (\sa_ctrl[30][15] , \sa_ctrl[30].r.part0[15] );
tran (\sa_ctrl[30][15] , \sa_ctrl[30].f.spare[10] );
tran (\sa_ctrl[30][16] , \sa_ctrl[30].r.part0[16] );
tran (\sa_ctrl[30][16] , \sa_ctrl[30].f.spare[11] );
tran (\sa_ctrl[30][17] , \sa_ctrl[30].r.part0[17] );
tran (\sa_ctrl[30][17] , \sa_ctrl[30].f.spare[12] );
tran (\sa_ctrl[30][18] , \sa_ctrl[30].r.part0[18] );
tran (\sa_ctrl[30][18] , \sa_ctrl[30].f.spare[13] );
tran (\sa_ctrl[30][19] , \sa_ctrl[30].r.part0[19] );
tran (\sa_ctrl[30][19] , \sa_ctrl[30].f.spare[14] );
tran (\sa_ctrl[30][20] , \sa_ctrl[30].r.part0[20] );
tran (\sa_ctrl[30][20] , \sa_ctrl[30].f.spare[15] );
tran (\sa_ctrl[30][21] , \sa_ctrl[30].r.part0[21] );
tran (\sa_ctrl[30][21] , \sa_ctrl[30].f.spare[16] );
tran (\sa_ctrl[30][22] , \sa_ctrl[30].r.part0[22] );
tran (\sa_ctrl[30][22] , \sa_ctrl[30].f.spare[17] );
tran (\sa_ctrl[30][23] , \sa_ctrl[30].r.part0[23] );
tran (\sa_ctrl[30][23] , \sa_ctrl[30].f.spare[18] );
tran (\sa_ctrl[30][24] , \sa_ctrl[30].r.part0[24] );
tran (\sa_ctrl[30][24] , \sa_ctrl[30].f.spare[19] );
tran (\sa_ctrl[30][25] , \sa_ctrl[30].r.part0[25] );
tran (\sa_ctrl[30][25] , \sa_ctrl[30].f.spare[20] );
tran (\sa_ctrl[30][26] , \sa_ctrl[30].r.part0[26] );
tran (\sa_ctrl[30][26] , \sa_ctrl[30].f.spare[21] );
tran (\sa_ctrl[30][27] , \sa_ctrl[30].r.part0[27] );
tran (\sa_ctrl[30][27] , \sa_ctrl[30].f.spare[22] );
tran (\sa_ctrl[30][28] , \sa_ctrl[30].r.part0[28] );
tran (\sa_ctrl[30][28] , \sa_ctrl[30].f.spare[23] );
tran (\sa_ctrl[30][29] , \sa_ctrl[30].r.part0[29] );
tran (\sa_ctrl[30][29] , \sa_ctrl[30].f.spare[24] );
tran (\sa_ctrl[30][30] , \sa_ctrl[30].r.part0[30] );
tran (\sa_ctrl[30][30] , \sa_ctrl[30].f.spare[25] );
tran (\sa_ctrl[30][31] , \sa_ctrl[30].r.part0[31] );
tran (\sa_ctrl[30][31] , \sa_ctrl[30].f.spare[26] );
tran (\sa_ctrl[31][0] , \sa_ctrl[31].r.part0[0] );
tran (\sa_ctrl[31][0] , \sa_ctrl[31].f.sa_event_sel[0] );
tran (\sa_ctrl[31][1] , \sa_ctrl[31].r.part0[1] );
tran (\sa_ctrl[31][1] , \sa_ctrl[31].f.sa_event_sel[1] );
tran (\sa_ctrl[31][2] , \sa_ctrl[31].r.part0[2] );
tran (\sa_ctrl[31][2] , \sa_ctrl[31].f.sa_event_sel[2] );
tran (\sa_ctrl[31][3] , \sa_ctrl[31].r.part0[3] );
tran (\sa_ctrl[31][3] , \sa_ctrl[31].f.sa_event_sel[3] );
tran (\sa_ctrl[31][4] , \sa_ctrl[31].r.part0[4] );
tran (\sa_ctrl[31][4] , \sa_ctrl[31].f.sa_event_sel[4] );
tran (\sa_ctrl[31][5] , \sa_ctrl[31].r.part0[5] );
tran (\sa_ctrl[31][5] , \sa_ctrl[31].f.spare[0] );
tran (\sa_ctrl[31][6] , \sa_ctrl[31].r.part0[6] );
tran (\sa_ctrl[31][6] , \sa_ctrl[31].f.spare[1] );
tran (\sa_ctrl[31][7] , \sa_ctrl[31].r.part0[7] );
tran (\sa_ctrl[31][7] , \sa_ctrl[31].f.spare[2] );
tran (\sa_ctrl[31][8] , \sa_ctrl[31].r.part0[8] );
tran (\sa_ctrl[31][8] , \sa_ctrl[31].f.spare[3] );
tran (\sa_ctrl[31][9] , \sa_ctrl[31].r.part0[9] );
tran (\sa_ctrl[31][9] , \sa_ctrl[31].f.spare[4] );
tran (\sa_ctrl[31][10] , \sa_ctrl[31].r.part0[10] );
tran (\sa_ctrl[31][10] , \sa_ctrl[31].f.spare[5] );
tran (\sa_ctrl[31][11] , \sa_ctrl[31].r.part0[11] );
tran (\sa_ctrl[31][11] , \sa_ctrl[31].f.spare[6] );
tran (\sa_ctrl[31][12] , \sa_ctrl[31].r.part0[12] );
tran (\sa_ctrl[31][12] , \sa_ctrl[31].f.spare[7] );
tran (\sa_ctrl[31][13] , \sa_ctrl[31].r.part0[13] );
tran (\sa_ctrl[31][13] , \sa_ctrl[31].f.spare[8] );
tran (\sa_ctrl[31][14] , \sa_ctrl[31].r.part0[14] );
tran (\sa_ctrl[31][14] , \sa_ctrl[31].f.spare[9] );
tran (\sa_ctrl[31][15] , \sa_ctrl[31].r.part0[15] );
tran (\sa_ctrl[31][15] , \sa_ctrl[31].f.spare[10] );
tran (\sa_ctrl[31][16] , \sa_ctrl[31].r.part0[16] );
tran (\sa_ctrl[31][16] , \sa_ctrl[31].f.spare[11] );
tran (\sa_ctrl[31][17] , \sa_ctrl[31].r.part0[17] );
tran (\sa_ctrl[31][17] , \sa_ctrl[31].f.spare[12] );
tran (\sa_ctrl[31][18] , \sa_ctrl[31].r.part0[18] );
tran (\sa_ctrl[31][18] , \sa_ctrl[31].f.spare[13] );
tran (\sa_ctrl[31][19] , \sa_ctrl[31].r.part0[19] );
tran (\sa_ctrl[31][19] , \sa_ctrl[31].f.spare[14] );
tran (\sa_ctrl[31][20] , \sa_ctrl[31].r.part0[20] );
tran (\sa_ctrl[31][20] , \sa_ctrl[31].f.spare[15] );
tran (\sa_ctrl[31][21] , \sa_ctrl[31].r.part0[21] );
tran (\sa_ctrl[31][21] , \sa_ctrl[31].f.spare[16] );
tran (\sa_ctrl[31][22] , \sa_ctrl[31].r.part0[22] );
tran (\sa_ctrl[31][22] , \sa_ctrl[31].f.spare[17] );
tran (\sa_ctrl[31][23] , \sa_ctrl[31].r.part0[23] );
tran (\sa_ctrl[31][23] , \sa_ctrl[31].f.spare[18] );
tran (\sa_ctrl[31][24] , \sa_ctrl[31].r.part0[24] );
tran (\sa_ctrl[31][24] , \sa_ctrl[31].f.spare[19] );
tran (\sa_ctrl[31][25] , \sa_ctrl[31].r.part0[25] );
tran (\sa_ctrl[31][25] , \sa_ctrl[31].f.spare[20] );
tran (\sa_ctrl[31][26] , \sa_ctrl[31].r.part0[26] );
tran (\sa_ctrl[31][26] , \sa_ctrl[31].f.spare[21] );
tran (\sa_ctrl[31][27] , \sa_ctrl[31].r.part0[27] );
tran (\sa_ctrl[31][27] , \sa_ctrl[31].f.spare[22] );
tran (\sa_ctrl[31][28] , \sa_ctrl[31].r.part0[28] );
tran (\sa_ctrl[31][28] , \sa_ctrl[31].f.spare[23] );
tran (\sa_ctrl[31][29] , \sa_ctrl[31].r.part0[29] );
tran (\sa_ctrl[31][29] , \sa_ctrl[31].f.spare[24] );
tran (\sa_ctrl[31][30] , \sa_ctrl[31].r.part0[30] );
tran (\sa_ctrl[31][30] , \sa_ctrl[31].f.spare[25] );
tran (\sa_ctrl[31][31] , \sa_ctrl[31].r.part0[31] );
tran (\sa_ctrl[31][31] , \sa_ctrl[31].f.spare[26] );
tran (rbus_ring_i[83], \rbus_ring_i.addr [15]);
tran (rbus_ring_i[82], \rbus_ring_i.addr [14]);
tran (rbus_ring_i[81], \rbus_ring_i.addr [13]);
tran (rbus_ring_i[80], \rbus_ring_i.addr [12]);
tran (rbus_ring_i[79], \rbus_ring_i.addr [11]);
tran (rbus_ring_i[78], \rbus_ring_i.addr [10]);
tran (rbus_ring_i[77], \rbus_ring_i.addr [9]);
tran (rbus_ring_i[76], \rbus_ring_i.addr [8]);
tran (rbus_ring_i[75], \rbus_ring_i.addr [7]);
tran (rbus_ring_i[74], \rbus_ring_i.addr [6]);
tran (rbus_ring_i[73], \rbus_ring_i.addr [5]);
tran (rbus_ring_i[72], \rbus_ring_i.addr [4]);
tran (rbus_ring_i[71], \rbus_ring_i.addr [3]);
tran (rbus_ring_i[70], \rbus_ring_i.addr [2]);
tran (rbus_ring_i[69], \rbus_ring_i.addr [1]);
tran (rbus_ring_i[68], \rbus_ring_i.addr [0]);
tran (rbus_ring_i[67], \rbus_ring_i.wr_strb );
tran (rbus_ring_i[66], \rbus_ring_i.wr_data [31]);
tran (rbus_ring_i[65], \rbus_ring_i.wr_data [30]);
tran (rbus_ring_i[64], \rbus_ring_i.wr_data [29]);
tran (rbus_ring_i[63], \rbus_ring_i.wr_data [28]);
tran (rbus_ring_i[62], \rbus_ring_i.wr_data [27]);
tran (rbus_ring_i[61], \rbus_ring_i.wr_data [26]);
tran (rbus_ring_i[60], \rbus_ring_i.wr_data [25]);
tran (rbus_ring_i[59], \rbus_ring_i.wr_data [24]);
tran (rbus_ring_i[58], \rbus_ring_i.wr_data [23]);
tran (rbus_ring_i[57], \rbus_ring_i.wr_data [22]);
tran (rbus_ring_i[56], \rbus_ring_i.wr_data [21]);
tran (rbus_ring_i[55], \rbus_ring_i.wr_data [20]);
tran (rbus_ring_i[54], \rbus_ring_i.wr_data [19]);
tran (rbus_ring_i[53], \rbus_ring_i.wr_data [18]);
tran (rbus_ring_i[52], \rbus_ring_i.wr_data [17]);
tran (rbus_ring_i[51], \rbus_ring_i.wr_data [16]);
tran (rbus_ring_i[50], \rbus_ring_i.wr_data [15]);
tran (rbus_ring_i[49], \rbus_ring_i.wr_data [14]);
tran (rbus_ring_i[48], \rbus_ring_i.wr_data [13]);
tran (rbus_ring_i[47], \rbus_ring_i.wr_data [12]);
tran (rbus_ring_i[46], \rbus_ring_i.wr_data [11]);
tran (rbus_ring_i[45], \rbus_ring_i.wr_data [10]);
tran (rbus_ring_i[44], \rbus_ring_i.wr_data [9]);
tran (rbus_ring_i[43], \rbus_ring_i.wr_data [8]);
tran (rbus_ring_i[42], \rbus_ring_i.wr_data [7]);
tran (rbus_ring_i[41], \rbus_ring_i.wr_data [6]);
tran (rbus_ring_i[40], \rbus_ring_i.wr_data [5]);
tran (rbus_ring_i[39], \rbus_ring_i.wr_data [4]);
tran (rbus_ring_i[38], \rbus_ring_i.wr_data [3]);
tran (rbus_ring_i[37], \rbus_ring_i.wr_data [2]);
tran (rbus_ring_i[36], \rbus_ring_i.wr_data [1]);
tran (rbus_ring_i[35], \rbus_ring_i.wr_data [0]);
tran (rbus_ring_i[34], \rbus_ring_i.rd_strb );
tran (rbus_ring_i[33], \rbus_ring_i.rd_data [31]);
tran (rbus_ring_i[32], \rbus_ring_i.rd_data [30]);
tran (rbus_ring_i[31], \rbus_ring_i.rd_data [29]);
tran (rbus_ring_i[30], \rbus_ring_i.rd_data [28]);
tran (rbus_ring_i[29], \rbus_ring_i.rd_data [27]);
tran (rbus_ring_i[28], \rbus_ring_i.rd_data [26]);
tran (rbus_ring_i[27], \rbus_ring_i.rd_data [25]);
tran (rbus_ring_i[26], \rbus_ring_i.rd_data [24]);
tran (rbus_ring_i[25], \rbus_ring_i.rd_data [23]);
tran (rbus_ring_i[24], \rbus_ring_i.rd_data [22]);
tran (rbus_ring_i[23], \rbus_ring_i.rd_data [21]);
tran (rbus_ring_i[22], \rbus_ring_i.rd_data [20]);
tran (rbus_ring_i[21], \rbus_ring_i.rd_data [19]);
tran (rbus_ring_i[20], \rbus_ring_i.rd_data [18]);
tran (rbus_ring_i[19], \rbus_ring_i.rd_data [17]);
tran (rbus_ring_i[18], \rbus_ring_i.rd_data [16]);
tran (rbus_ring_i[17], \rbus_ring_i.rd_data [15]);
tran (rbus_ring_i[16], \rbus_ring_i.rd_data [14]);
tran (rbus_ring_i[15], \rbus_ring_i.rd_data [13]);
tran (rbus_ring_i[14], \rbus_ring_i.rd_data [12]);
tran (rbus_ring_i[13], \rbus_ring_i.rd_data [11]);
tran (rbus_ring_i[12], \rbus_ring_i.rd_data [10]);
tran (rbus_ring_i[11], \rbus_ring_i.rd_data [9]);
tran (rbus_ring_i[10], \rbus_ring_i.rd_data [8]);
tran (rbus_ring_i[9], \rbus_ring_i.rd_data [7]);
tran (rbus_ring_i[8], \rbus_ring_i.rd_data [6]);
tran (rbus_ring_i[7], \rbus_ring_i.rd_data [5]);
tran (rbus_ring_i[6], \rbus_ring_i.rd_data [4]);
tran (rbus_ring_i[5], \rbus_ring_i.rd_data [3]);
tran (rbus_ring_i[4], \rbus_ring_i.rd_data [2]);
tran (rbus_ring_i[3], \rbus_ring_i.rd_data [1]);
tran (rbus_ring_i[2], \rbus_ring_i.rd_data [0]);
tran (rbus_ring_i[1], \rbus_ring_i.ack );
tran (rbus_ring_i[0], \rbus_ring_i.err_ack );
tran (kme_cceip0_ob_out_pre[82], \kme_cceip0_ob_out_pre.tvalid );
tran (kme_cceip0_ob_out_pre[81], \kme_cceip0_ob_out_pre.tlast );
tran (kme_cceip0_ob_out_pre[80], \kme_cceip0_ob_out_pre.tid [0]);
tran (kme_cceip0_ob_out_pre[79], \kme_cceip0_ob_out_pre.tstrb [7]);
tran (kme_cceip0_ob_out_pre[78], \kme_cceip0_ob_out_pre.tstrb [6]);
tran (kme_cceip0_ob_out_pre[77], \kme_cceip0_ob_out_pre.tstrb [5]);
tran (kme_cceip0_ob_out_pre[76], \kme_cceip0_ob_out_pre.tstrb [4]);
tran (kme_cceip0_ob_out_pre[75], \kme_cceip0_ob_out_pre.tstrb [3]);
tran (kme_cceip0_ob_out_pre[74], \kme_cceip0_ob_out_pre.tstrb [2]);
tran (kme_cceip0_ob_out_pre[73], \kme_cceip0_ob_out_pre.tstrb [1]);
tran (kme_cceip0_ob_out_pre[72], \kme_cceip0_ob_out_pre.tstrb [0]);
tran (kme_cceip0_ob_out_pre[71], \kme_cceip0_ob_out_pre.tuser [7]);
tran (kme_cceip0_ob_out_pre[70], \kme_cceip0_ob_out_pre.tuser [6]);
tran (kme_cceip0_ob_out_pre[69], \kme_cceip0_ob_out_pre.tuser [5]);
tran (kme_cceip0_ob_out_pre[68], \kme_cceip0_ob_out_pre.tuser [4]);
tran (kme_cceip0_ob_out_pre[67], \kme_cceip0_ob_out_pre.tuser [3]);
tran (kme_cceip0_ob_out_pre[66], \kme_cceip0_ob_out_pre.tuser [2]);
tran (kme_cceip0_ob_out_pre[65], \kme_cceip0_ob_out_pre.tuser [1]);
tran (kme_cceip0_ob_out_pre[64], \kme_cceip0_ob_out_pre.tuser [0]);
tran (kme_cceip0_ob_out_pre[63], \kme_cceip0_ob_out_pre.tdata [63]);
tran (kme_cceip0_ob_out_pre[62], \kme_cceip0_ob_out_pre.tdata [62]);
tran (kme_cceip0_ob_out_pre[61], \kme_cceip0_ob_out_pre.tdata [61]);
tran (kme_cceip0_ob_out_pre[60], \kme_cceip0_ob_out_pre.tdata [60]);
tran (kme_cceip0_ob_out_pre[59], \kme_cceip0_ob_out_pre.tdata [59]);
tran (kme_cceip0_ob_out_pre[58], \kme_cceip0_ob_out_pre.tdata [58]);
tran (kme_cceip0_ob_out_pre[57], \kme_cceip0_ob_out_pre.tdata [57]);
tran (kme_cceip0_ob_out_pre[56], \kme_cceip0_ob_out_pre.tdata [56]);
tran (kme_cceip0_ob_out_pre[55], \kme_cceip0_ob_out_pre.tdata [55]);
tran (kme_cceip0_ob_out_pre[54], \kme_cceip0_ob_out_pre.tdata [54]);
tran (kme_cceip0_ob_out_pre[53], \kme_cceip0_ob_out_pre.tdata [53]);
tran (kme_cceip0_ob_out_pre[52], \kme_cceip0_ob_out_pre.tdata [52]);
tran (kme_cceip0_ob_out_pre[51], \kme_cceip0_ob_out_pre.tdata [51]);
tran (kme_cceip0_ob_out_pre[50], \kme_cceip0_ob_out_pre.tdata [50]);
tran (kme_cceip0_ob_out_pre[49], \kme_cceip0_ob_out_pre.tdata [49]);
tran (kme_cceip0_ob_out_pre[48], \kme_cceip0_ob_out_pre.tdata [48]);
tran (kme_cceip0_ob_out_pre[47], \kme_cceip0_ob_out_pre.tdata [47]);
tran (kme_cceip0_ob_out_pre[46], \kme_cceip0_ob_out_pre.tdata [46]);
tran (kme_cceip0_ob_out_pre[45], \kme_cceip0_ob_out_pre.tdata [45]);
tran (kme_cceip0_ob_out_pre[44], \kme_cceip0_ob_out_pre.tdata [44]);
tran (kme_cceip0_ob_out_pre[43], \kme_cceip0_ob_out_pre.tdata [43]);
tran (kme_cceip0_ob_out_pre[42], \kme_cceip0_ob_out_pre.tdata [42]);
tran (kme_cceip0_ob_out_pre[41], \kme_cceip0_ob_out_pre.tdata [41]);
tran (kme_cceip0_ob_out_pre[40], \kme_cceip0_ob_out_pre.tdata [40]);
tran (kme_cceip0_ob_out_pre[39], \kme_cceip0_ob_out_pre.tdata [39]);
tran (kme_cceip0_ob_out_pre[38], \kme_cceip0_ob_out_pre.tdata [38]);
tran (kme_cceip0_ob_out_pre[37], \kme_cceip0_ob_out_pre.tdata [37]);
tran (kme_cceip0_ob_out_pre[36], \kme_cceip0_ob_out_pre.tdata [36]);
tran (kme_cceip0_ob_out_pre[35], \kme_cceip0_ob_out_pre.tdata [35]);
tran (kme_cceip0_ob_out_pre[34], \kme_cceip0_ob_out_pre.tdata [34]);
tran (kme_cceip0_ob_out_pre[33], \kme_cceip0_ob_out_pre.tdata [33]);
tran (kme_cceip0_ob_out_pre[32], \kme_cceip0_ob_out_pre.tdata [32]);
tran (kme_cceip0_ob_out_pre[31], \kme_cceip0_ob_out_pre.tdata [31]);
tran (kme_cceip0_ob_out_pre[30], \kme_cceip0_ob_out_pre.tdata [30]);
tran (kme_cceip0_ob_out_pre[29], \kme_cceip0_ob_out_pre.tdata [29]);
tran (kme_cceip0_ob_out_pre[28], \kme_cceip0_ob_out_pre.tdata [28]);
tran (kme_cceip0_ob_out_pre[27], \kme_cceip0_ob_out_pre.tdata [27]);
tran (kme_cceip0_ob_out_pre[26], \kme_cceip0_ob_out_pre.tdata [26]);
tran (kme_cceip0_ob_out_pre[25], \kme_cceip0_ob_out_pre.tdata [25]);
tran (kme_cceip0_ob_out_pre[24], \kme_cceip0_ob_out_pre.tdata [24]);
tran (kme_cceip0_ob_out_pre[23], \kme_cceip0_ob_out_pre.tdata [23]);
tran (kme_cceip0_ob_out_pre[22], \kme_cceip0_ob_out_pre.tdata [22]);
tran (kme_cceip0_ob_out_pre[21], \kme_cceip0_ob_out_pre.tdata [21]);
tran (kme_cceip0_ob_out_pre[20], \kme_cceip0_ob_out_pre.tdata [20]);
tran (kme_cceip0_ob_out_pre[19], \kme_cceip0_ob_out_pre.tdata [19]);
tran (kme_cceip0_ob_out_pre[18], \kme_cceip0_ob_out_pre.tdata [18]);
tran (kme_cceip0_ob_out_pre[17], \kme_cceip0_ob_out_pre.tdata [17]);
tran (kme_cceip0_ob_out_pre[16], \kme_cceip0_ob_out_pre.tdata [16]);
tran (kme_cceip0_ob_out_pre[15], \kme_cceip0_ob_out_pre.tdata [15]);
tran (kme_cceip0_ob_out_pre[14], \kme_cceip0_ob_out_pre.tdata [14]);
tran (kme_cceip0_ob_out_pre[13], \kme_cceip0_ob_out_pre.tdata [13]);
tran (kme_cceip0_ob_out_pre[12], \kme_cceip0_ob_out_pre.tdata [12]);
tran (kme_cceip0_ob_out_pre[11], \kme_cceip0_ob_out_pre.tdata [11]);
tran (kme_cceip0_ob_out_pre[10], \kme_cceip0_ob_out_pre.tdata [10]);
tran (kme_cceip0_ob_out_pre[9], \kme_cceip0_ob_out_pre.tdata [9]);
tran (kme_cceip0_ob_out_pre[8], \kme_cceip0_ob_out_pre.tdata [8]);
tran (kme_cceip0_ob_out_pre[7], \kme_cceip0_ob_out_pre.tdata [7]);
tran (kme_cceip0_ob_out_pre[6], \kme_cceip0_ob_out_pre.tdata [6]);
tran (kme_cceip0_ob_out_pre[5], \kme_cceip0_ob_out_pre.tdata [5]);
tran (kme_cceip0_ob_out_pre[4], \kme_cceip0_ob_out_pre.tdata [4]);
tran (kme_cceip0_ob_out_pre[3], \kme_cceip0_ob_out_pre.tdata [3]);
tran (kme_cceip0_ob_out_pre[2], \kme_cceip0_ob_out_pre.tdata [2]);
tran (kme_cceip0_ob_out_pre[1], \kme_cceip0_ob_out_pre.tdata [1]);
tran (kme_cceip0_ob_out_pre[0], \kme_cceip0_ob_out_pre.tdata [0]);
tran (kme_cceip0_ob_in[0], \kme_cceip0_ob_in.tready );
tran (kme_cceip1_ob_out_pre[82], \kme_cceip1_ob_out_pre.tvalid );
tran (kme_cceip1_ob_out_pre[81], \kme_cceip1_ob_out_pre.tlast );
tran (kme_cceip1_ob_out_pre[80], \kme_cceip1_ob_out_pre.tid [0]);
tran (kme_cceip1_ob_out_pre[79], \kme_cceip1_ob_out_pre.tstrb [7]);
tran (kme_cceip1_ob_out_pre[78], \kme_cceip1_ob_out_pre.tstrb [6]);
tran (kme_cceip1_ob_out_pre[77], \kme_cceip1_ob_out_pre.tstrb [5]);
tran (kme_cceip1_ob_out_pre[76], \kme_cceip1_ob_out_pre.tstrb [4]);
tran (kme_cceip1_ob_out_pre[75], \kme_cceip1_ob_out_pre.tstrb [3]);
tran (kme_cceip1_ob_out_pre[74], \kme_cceip1_ob_out_pre.tstrb [2]);
tran (kme_cceip1_ob_out_pre[73], \kme_cceip1_ob_out_pre.tstrb [1]);
tran (kme_cceip1_ob_out_pre[72], \kme_cceip1_ob_out_pre.tstrb [0]);
tran (kme_cceip1_ob_out_pre[71], \kme_cceip1_ob_out_pre.tuser [7]);
tran (kme_cceip1_ob_out_pre[70], \kme_cceip1_ob_out_pre.tuser [6]);
tran (kme_cceip1_ob_out_pre[69], \kme_cceip1_ob_out_pre.tuser [5]);
tran (kme_cceip1_ob_out_pre[68], \kme_cceip1_ob_out_pre.tuser [4]);
tran (kme_cceip1_ob_out_pre[67], \kme_cceip1_ob_out_pre.tuser [3]);
tran (kme_cceip1_ob_out_pre[66], \kme_cceip1_ob_out_pre.tuser [2]);
tran (kme_cceip1_ob_out_pre[65], \kme_cceip1_ob_out_pre.tuser [1]);
tran (kme_cceip1_ob_out_pre[64], \kme_cceip1_ob_out_pre.tuser [0]);
tran (kme_cceip1_ob_out_pre[63], \kme_cceip1_ob_out_pre.tdata [63]);
tran (kme_cceip1_ob_out_pre[62], \kme_cceip1_ob_out_pre.tdata [62]);
tran (kme_cceip1_ob_out_pre[61], \kme_cceip1_ob_out_pre.tdata [61]);
tran (kme_cceip1_ob_out_pre[60], \kme_cceip1_ob_out_pre.tdata [60]);
tran (kme_cceip1_ob_out_pre[59], \kme_cceip1_ob_out_pre.tdata [59]);
tran (kme_cceip1_ob_out_pre[58], \kme_cceip1_ob_out_pre.tdata [58]);
tran (kme_cceip1_ob_out_pre[57], \kme_cceip1_ob_out_pre.tdata [57]);
tran (kme_cceip1_ob_out_pre[56], \kme_cceip1_ob_out_pre.tdata [56]);
tran (kme_cceip1_ob_out_pre[55], \kme_cceip1_ob_out_pre.tdata [55]);
tran (kme_cceip1_ob_out_pre[54], \kme_cceip1_ob_out_pre.tdata [54]);
tran (kme_cceip1_ob_out_pre[53], \kme_cceip1_ob_out_pre.tdata [53]);
tran (kme_cceip1_ob_out_pre[52], \kme_cceip1_ob_out_pre.tdata [52]);
tran (kme_cceip1_ob_out_pre[51], \kme_cceip1_ob_out_pre.tdata [51]);
tran (kme_cceip1_ob_out_pre[50], \kme_cceip1_ob_out_pre.tdata [50]);
tran (kme_cceip1_ob_out_pre[49], \kme_cceip1_ob_out_pre.tdata [49]);
tran (kme_cceip1_ob_out_pre[48], \kme_cceip1_ob_out_pre.tdata [48]);
tran (kme_cceip1_ob_out_pre[47], \kme_cceip1_ob_out_pre.tdata [47]);
tran (kme_cceip1_ob_out_pre[46], \kme_cceip1_ob_out_pre.tdata [46]);
tran (kme_cceip1_ob_out_pre[45], \kme_cceip1_ob_out_pre.tdata [45]);
tran (kme_cceip1_ob_out_pre[44], \kme_cceip1_ob_out_pre.tdata [44]);
tran (kme_cceip1_ob_out_pre[43], \kme_cceip1_ob_out_pre.tdata [43]);
tran (kme_cceip1_ob_out_pre[42], \kme_cceip1_ob_out_pre.tdata [42]);
tran (kme_cceip1_ob_out_pre[41], \kme_cceip1_ob_out_pre.tdata [41]);
tran (kme_cceip1_ob_out_pre[40], \kme_cceip1_ob_out_pre.tdata [40]);
tran (kme_cceip1_ob_out_pre[39], \kme_cceip1_ob_out_pre.tdata [39]);
tran (kme_cceip1_ob_out_pre[38], \kme_cceip1_ob_out_pre.tdata [38]);
tran (kme_cceip1_ob_out_pre[37], \kme_cceip1_ob_out_pre.tdata [37]);
tran (kme_cceip1_ob_out_pre[36], \kme_cceip1_ob_out_pre.tdata [36]);
tran (kme_cceip1_ob_out_pre[35], \kme_cceip1_ob_out_pre.tdata [35]);
tran (kme_cceip1_ob_out_pre[34], \kme_cceip1_ob_out_pre.tdata [34]);
tran (kme_cceip1_ob_out_pre[33], \kme_cceip1_ob_out_pre.tdata [33]);
tran (kme_cceip1_ob_out_pre[32], \kme_cceip1_ob_out_pre.tdata [32]);
tran (kme_cceip1_ob_out_pre[31], \kme_cceip1_ob_out_pre.tdata [31]);
tran (kme_cceip1_ob_out_pre[30], \kme_cceip1_ob_out_pre.tdata [30]);
tran (kme_cceip1_ob_out_pre[29], \kme_cceip1_ob_out_pre.tdata [29]);
tran (kme_cceip1_ob_out_pre[28], \kme_cceip1_ob_out_pre.tdata [28]);
tran (kme_cceip1_ob_out_pre[27], \kme_cceip1_ob_out_pre.tdata [27]);
tran (kme_cceip1_ob_out_pre[26], \kme_cceip1_ob_out_pre.tdata [26]);
tran (kme_cceip1_ob_out_pre[25], \kme_cceip1_ob_out_pre.tdata [25]);
tran (kme_cceip1_ob_out_pre[24], \kme_cceip1_ob_out_pre.tdata [24]);
tran (kme_cceip1_ob_out_pre[23], \kme_cceip1_ob_out_pre.tdata [23]);
tran (kme_cceip1_ob_out_pre[22], \kme_cceip1_ob_out_pre.tdata [22]);
tran (kme_cceip1_ob_out_pre[21], \kme_cceip1_ob_out_pre.tdata [21]);
tran (kme_cceip1_ob_out_pre[20], \kme_cceip1_ob_out_pre.tdata [20]);
tran (kme_cceip1_ob_out_pre[19], \kme_cceip1_ob_out_pre.tdata [19]);
tran (kme_cceip1_ob_out_pre[18], \kme_cceip1_ob_out_pre.tdata [18]);
tran (kme_cceip1_ob_out_pre[17], \kme_cceip1_ob_out_pre.tdata [17]);
tran (kme_cceip1_ob_out_pre[16], \kme_cceip1_ob_out_pre.tdata [16]);
tran (kme_cceip1_ob_out_pre[15], \kme_cceip1_ob_out_pre.tdata [15]);
tran (kme_cceip1_ob_out_pre[14], \kme_cceip1_ob_out_pre.tdata [14]);
tran (kme_cceip1_ob_out_pre[13], \kme_cceip1_ob_out_pre.tdata [13]);
tran (kme_cceip1_ob_out_pre[12], \kme_cceip1_ob_out_pre.tdata [12]);
tran (kme_cceip1_ob_out_pre[11], \kme_cceip1_ob_out_pre.tdata [11]);
tran (kme_cceip1_ob_out_pre[10], \kme_cceip1_ob_out_pre.tdata [10]);
tran (kme_cceip1_ob_out_pre[9], \kme_cceip1_ob_out_pre.tdata [9]);
tran (kme_cceip1_ob_out_pre[8], \kme_cceip1_ob_out_pre.tdata [8]);
tran (kme_cceip1_ob_out_pre[7], \kme_cceip1_ob_out_pre.tdata [7]);
tran (kme_cceip1_ob_out_pre[6], \kme_cceip1_ob_out_pre.tdata [6]);
tran (kme_cceip1_ob_out_pre[5], \kme_cceip1_ob_out_pre.tdata [5]);
tran (kme_cceip1_ob_out_pre[4], \kme_cceip1_ob_out_pre.tdata [4]);
tran (kme_cceip1_ob_out_pre[3], \kme_cceip1_ob_out_pre.tdata [3]);
tran (kme_cceip1_ob_out_pre[2], \kme_cceip1_ob_out_pre.tdata [2]);
tran (kme_cceip1_ob_out_pre[1], \kme_cceip1_ob_out_pre.tdata [1]);
tran (kme_cceip1_ob_out_pre[0], \kme_cceip1_ob_out_pre.tdata [0]);
tran (kme_cceip1_ob_in[0], \kme_cceip1_ob_in.tready );
tran (kme_cceip2_ob_out_pre[82], \kme_cceip2_ob_out_pre.tvalid );
tran (kme_cceip2_ob_out_pre[81], \kme_cceip2_ob_out_pre.tlast );
tran (kme_cceip2_ob_out_pre[80], \kme_cceip2_ob_out_pre.tid [0]);
tran (kme_cceip2_ob_out_pre[79], \kme_cceip2_ob_out_pre.tstrb [7]);
tran (kme_cceip2_ob_out_pre[78], \kme_cceip2_ob_out_pre.tstrb [6]);
tran (kme_cceip2_ob_out_pre[77], \kme_cceip2_ob_out_pre.tstrb [5]);
tran (kme_cceip2_ob_out_pre[76], \kme_cceip2_ob_out_pre.tstrb [4]);
tran (kme_cceip2_ob_out_pre[75], \kme_cceip2_ob_out_pre.tstrb [3]);
tran (kme_cceip2_ob_out_pre[74], \kme_cceip2_ob_out_pre.tstrb [2]);
tran (kme_cceip2_ob_out_pre[73], \kme_cceip2_ob_out_pre.tstrb [1]);
tran (kme_cceip2_ob_out_pre[72], \kme_cceip2_ob_out_pre.tstrb [0]);
tran (kme_cceip2_ob_out_pre[71], \kme_cceip2_ob_out_pre.tuser [7]);
tran (kme_cceip2_ob_out_pre[70], \kme_cceip2_ob_out_pre.tuser [6]);
tran (kme_cceip2_ob_out_pre[69], \kme_cceip2_ob_out_pre.tuser [5]);
tran (kme_cceip2_ob_out_pre[68], \kme_cceip2_ob_out_pre.tuser [4]);
tran (kme_cceip2_ob_out_pre[67], \kme_cceip2_ob_out_pre.tuser [3]);
tran (kme_cceip2_ob_out_pre[66], \kme_cceip2_ob_out_pre.tuser [2]);
tran (kme_cceip2_ob_out_pre[65], \kme_cceip2_ob_out_pre.tuser [1]);
tran (kme_cceip2_ob_out_pre[64], \kme_cceip2_ob_out_pre.tuser [0]);
tran (kme_cceip2_ob_out_pre[63], \kme_cceip2_ob_out_pre.tdata [63]);
tran (kme_cceip2_ob_out_pre[62], \kme_cceip2_ob_out_pre.tdata [62]);
tran (kme_cceip2_ob_out_pre[61], \kme_cceip2_ob_out_pre.tdata [61]);
tran (kme_cceip2_ob_out_pre[60], \kme_cceip2_ob_out_pre.tdata [60]);
tran (kme_cceip2_ob_out_pre[59], \kme_cceip2_ob_out_pre.tdata [59]);
tran (kme_cceip2_ob_out_pre[58], \kme_cceip2_ob_out_pre.tdata [58]);
tran (kme_cceip2_ob_out_pre[57], \kme_cceip2_ob_out_pre.tdata [57]);
tran (kme_cceip2_ob_out_pre[56], \kme_cceip2_ob_out_pre.tdata [56]);
tran (kme_cceip2_ob_out_pre[55], \kme_cceip2_ob_out_pre.tdata [55]);
tran (kme_cceip2_ob_out_pre[54], \kme_cceip2_ob_out_pre.tdata [54]);
tran (kme_cceip2_ob_out_pre[53], \kme_cceip2_ob_out_pre.tdata [53]);
tran (kme_cceip2_ob_out_pre[52], \kme_cceip2_ob_out_pre.tdata [52]);
tran (kme_cceip2_ob_out_pre[51], \kme_cceip2_ob_out_pre.tdata [51]);
tran (kme_cceip2_ob_out_pre[50], \kme_cceip2_ob_out_pre.tdata [50]);
tran (kme_cceip2_ob_out_pre[49], \kme_cceip2_ob_out_pre.tdata [49]);
tran (kme_cceip2_ob_out_pre[48], \kme_cceip2_ob_out_pre.tdata [48]);
tran (kme_cceip2_ob_out_pre[47], \kme_cceip2_ob_out_pre.tdata [47]);
tran (kme_cceip2_ob_out_pre[46], \kme_cceip2_ob_out_pre.tdata [46]);
tran (kme_cceip2_ob_out_pre[45], \kme_cceip2_ob_out_pre.tdata [45]);
tran (kme_cceip2_ob_out_pre[44], \kme_cceip2_ob_out_pre.tdata [44]);
tran (kme_cceip2_ob_out_pre[43], \kme_cceip2_ob_out_pre.tdata [43]);
tran (kme_cceip2_ob_out_pre[42], \kme_cceip2_ob_out_pre.tdata [42]);
tran (kme_cceip2_ob_out_pre[41], \kme_cceip2_ob_out_pre.tdata [41]);
tran (kme_cceip2_ob_out_pre[40], \kme_cceip2_ob_out_pre.tdata [40]);
tran (kme_cceip2_ob_out_pre[39], \kme_cceip2_ob_out_pre.tdata [39]);
tran (kme_cceip2_ob_out_pre[38], \kme_cceip2_ob_out_pre.tdata [38]);
tran (kme_cceip2_ob_out_pre[37], \kme_cceip2_ob_out_pre.tdata [37]);
tran (kme_cceip2_ob_out_pre[36], \kme_cceip2_ob_out_pre.tdata [36]);
tran (kme_cceip2_ob_out_pre[35], \kme_cceip2_ob_out_pre.tdata [35]);
tran (kme_cceip2_ob_out_pre[34], \kme_cceip2_ob_out_pre.tdata [34]);
tran (kme_cceip2_ob_out_pre[33], \kme_cceip2_ob_out_pre.tdata [33]);
tran (kme_cceip2_ob_out_pre[32], \kme_cceip2_ob_out_pre.tdata [32]);
tran (kme_cceip2_ob_out_pre[31], \kme_cceip2_ob_out_pre.tdata [31]);
tran (kme_cceip2_ob_out_pre[30], \kme_cceip2_ob_out_pre.tdata [30]);
tran (kme_cceip2_ob_out_pre[29], \kme_cceip2_ob_out_pre.tdata [29]);
tran (kme_cceip2_ob_out_pre[28], \kme_cceip2_ob_out_pre.tdata [28]);
tran (kme_cceip2_ob_out_pre[27], \kme_cceip2_ob_out_pre.tdata [27]);
tran (kme_cceip2_ob_out_pre[26], \kme_cceip2_ob_out_pre.tdata [26]);
tran (kme_cceip2_ob_out_pre[25], \kme_cceip2_ob_out_pre.tdata [25]);
tran (kme_cceip2_ob_out_pre[24], \kme_cceip2_ob_out_pre.tdata [24]);
tran (kme_cceip2_ob_out_pre[23], \kme_cceip2_ob_out_pre.tdata [23]);
tran (kme_cceip2_ob_out_pre[22], \kme_cceip2_ob_out_pre.tdata [22]);
tran (kme_cceip2_ob_out_pre[21], \kme_cceip2_ob_out_pre.tdata [21]);
tran (kme_cceip2_ob_out_pre[20], \kme_cceip2_ob_out_pre.tdata [20]);
tran (kme_cceip2_ob_out_pre[19], \kme_cceip2_ob_out_pre.tdata [19]);
tran (kme_cceip2_ob_out_pre[18], \kme_cceip2_ob_out_pre.tdata [18]);
tran (kme_cceip2_ob_out_pre[17], \kme_cceip2_ob_out_pre.tdata [17]);
tran (kme_cceip2_ob_out_pre[16], \kme_cceip2_ob_out_pre.tdata [16]);
tran (kme_cceip2_ob_out_pre[15], \kme_cceip2_ob_out_pre.tdata [15]);
tran (kme_cceip2_ob_out_pre[14], \kme_cceip2_ob_out_pre.tdata [14]);
tran (kme_cceip2_ob_out_pre[13], \kme_cceip2_ob_out_pre.tdata [13]);
tran (kme_cceip2_ob_out_pre[12], \kme_cceip2_ob_out_pre.tdata [12]);
tran (kme_cceip2_ob_out_pre[11], \kme_cceip2_ob_out_pre.tdata [11]);
tran (kme_cceip2_ob_out_pre[10], \kme_cceip2_ob_out_pre.tdata [10]);
tran (kme_cceip2_ob_out_pre[9], \kme_cceip2_ob_out_pre.tdata [9]);
tran (kme_cceip2_ob_out_pre[8], \kme_cceip2_ob_out_pre.tdata [8]);
tran (kme_cceip2_ob_out_pre[7], \kme_cceip2_ob_out_pre.tdata [7]);
tran (kme_cceip2_ob_out_pre[6], \kme_cceip2_ob_out_pre.tdata [6]);
tran (kme_cceip2_ob_out_pre[5], \kme_cceip2_ob_out_pre.tdata [5]);
tran (kme_cceip2_ob_out_pre[4], \kme_cceip2_ob_out_pre.tdata [4]);
tran (kme_cceip2_ob_out_pre[3], \kme_cceip2_ob_out_pre.tdata [3]);
tran (kme_cceip2_ob_out_pre[2], \kme_cceip2_ob_out_pre.tdata [2]);
tran (kme_cceip2_ob_out_pre[1], \kme_cceip2_ob_out_pre.tdata [1]);
tran (kme_cceip2_ob_out_pre[0], \kme_cceip2_ob_out_pre.tdata [0]);
tran (kme_cceip2_ob_in[0], \kme_cceip2_ob_in.tready );
tran (kme_cceip3_ob_out_pre[82], \kme_cceip3_ob_out_pre.tvalid );
tran (kme_cceip3_ob_out_pre[81], \kme_cceip3_ob_out_pre.tlast );
tran (kme_cceip3_ob_out_pre[80], \kme_cceip3_ob_out_pre.tid [0]);
tran (kme_cceip3_ob_out_pre[79], \kme_cceip3_ob_out_pre.tstrb [7]);
tran (kme_cceip3_ob_out_pre[78], \kme_cceip3_ob_out_pre.tstrb [6]);
tran (kme_cceip3_ob_out_pre[77], \kme_cceip3_ob_out_pre.tstrb [5]);
tran (kme_cceip3_ob_out_pre[76], \kme_cceip3_ob_out_pre.tstrb [4]);
tran (kme_cceip3_ob_out_pre[75], \kme_cceip3_ob_out_pre.tstrb [3]);
tran (kme_cceip3_ob_out_pre[74], \kme_cceip3_ob_out_pre.tstrb [2]);
tran (kme_cceip3_ob_out_pre[73], \kme_cceip3_ob_out_pre.tstrb [1]);
tran (kme_cceip3_ob_out_pre[72], \kme_cceip3_ob_out_pre.tstrb [0]);
tran (kme_cceip3_ob_out_pre[71], \kme_cceip3_ob_out_pre.tuser [7]);
tran (kme_cceip3_ob_out_pre[70], \kme_cceip3_ob_out_pre.tuser [6]);
tran (kme_cceip3_ob_out_pre[69], \kme_cceip3_ob_out_pre.tuser [5]);
tran (kme_cceip3_ob_out_pre[68], \kme_cceip3_ob_out_pre.tuser [4]);
tran (kme_cceip3_ob_out_pre[67], \kme_cceip3_ob_out_pre.tuser [3]);
tran (kme_cceip3_ob_out_pre[66], \kme_cceip3_ob_out_pre.tuser [2]);
tran (kme_cceip3_ob_out_pre[65], \kme_cceip3_ob_out_pre.tuser [1]);
tran (kme_cceip3_ob_out_pre[64], \kme_cceip3_ob_out_pre.tuser [0]);
tran (kme_cceip3_ob_out_pre[63], \kme_cceip3_ob_out_pre.tdata [63]);
tran (kme_cceip3_ob_out_pre[62], \kme_cceip3_ob_out_pre.tdata [62]);
tran (kme_cceip3_ob_out_pre[61], \kme_cceip3_ob_out_pre.tdata [61]);
tran (kme_cceip3_ob_out_pre[60], \kme_cceip3_ob_out_pre.tdata [60]);
tran (kme_cceip3_ob_out_pre[59], \kme_cceip3_ob_out_pre.tdata [59]);
tran (kme_cceip3_ob_out_pre[58], \kme_cceip3_ob_out_pre.tdata [58]);
tran (kme_cceip3_ob_out_pre[57], \kme_cceip3_ob_out_pre.tdata [57]);
tran (kme_cceip3_ob_out_pre[56], \kme_cceip3_ob_out_pre.tdata [56]);
tran (kme_cceip3_ob_out_pre[55], \kme_cceip3_ob_out_pre.tdata [55]);
tran (kme_cceip3_ob_out_pre[54], \kme_cceip3_ob_out_pre.tdata [54]);
tran (kme_cceip3_ob_out_pre[53], \kme_cceip3_ob_out_pre.tdata [53]);
tran (kme_cceip3_ob_out_pre[52], \kme_cceip3_ob_out_pre.tdata [52]);
tran (kme_cceip3_ob_out_pre[51], \kme_cceip3_ob_out_pre.tdata [51]);
tran (kme_cceip3_ob_out_pre[50], \kme_cceip3_ob_out_pre.tdata [50]);
tran (kme_cceip3_ob_out_pre[49], \kme_cceip3_ob_out_pre.tdata [49]);
tran (kme_cceip3_ob_out_pre[48], \kme_cceip3_ob_out_pre.tdata [48]);
tran (kme_cceip3_ob_out_pre[47], \kme_cceip3_ob_out_pre.tdata [47]);
tran (kme_cceip3_ob_out_pre[46], \kme_cceip3_ob_out_pre.tdata [46]);
tran (kme_cceip3_ob_out_pre[45], \kme_cceip3_ob_out_pre.tdata [45]);
tran (kme_cceip3_ob_out_pre[44], \kme_cceip3_ob_out_pre.tdata [44]);
tran (kme_cceip3_ob_out_pre[43], \kme_cceip3_ob_out_pre.tdata [43]);
tran (kme_cceip3_ob_out_pre[42], \kme_cceip3_ob_out_pre.tdata [42]);
tran (kme_cceip3_ob_out_pre[41], \kme_cceip3_ob_out_pre.tdata [41]);
tran (kme_cceip3_ob_out_pre[40], \kme_cceip3_ob_out_pre.tdata [40]);
tran (kme_cceip3_ob_out_pre[39], \kme_cceip3_ob_out_pre.tdata [39]);
tran (kme_cceip3_ob_out_pre[38], \kme_cceip3_ob_out_pre.tdata [38]);
tran (kme_cceip3_ob_out_pre[37], \kme_cceip3_ob_out_pre.tdata [37]);
tran (kme_cceip3_ob_out_pre[36], \kme_cceip3_ob_out_pre.tdata [36]);
tran (kme_cceip3_ob_out_pre[35], \kme_cceip3_ob_out_pre.tdata [35]);
tran (kme_cceip3_ob_out_pre[34], \kme_cceip3_ob_out_pre.tdata [34]);
tran (kme_cceip3_ob_out_pre[33], \kme_cceip3_ob_out_pre.tdata [33]);
tran (kme_cceip3_ob_out_pre[32], \kme_cceip3_ob_out_pre.tdata [32]);
tran (kme_cceip3_ob_out_pre[31], \kme_cceip3_ob_out_pre.tdata [31]);
tran (kme_cceip3_ob_out_pre[30], \kme_cceip3_ob_out_pre.tdata [30]);
tran (kme_cceip3_ob_out_pre[29], \kme_cceip3_ob_out_pre.tdata [29]);
tran (kme_cceip3_ob_out_pre[28], \kme_cceip3_ob_out_pre.tdata [28]);
tran (kme_cceip3_ob_out_pre[27], \kme_cceip3_ob_out_pre.tdata [27]);
tran (kme_cceip3_ob_out_pre[26], \kme_cceip3_ob_out_pre.tdata [26]);
tran (kme_cceip3_ob_out_pre[25], \kme_cceip3_ob_out_pre.tdata [25]);
tran (kme_cceip3_ob_out_pre[24], \kme_cceip3_ob_out_pre.tdata [24]);
tran (kme_cceip3_ob_out_pre[23], \kme_cceip3_ob_out_pre.tdata [23]);
tran (kme_cceip3_ob_out_pre[22], \kme_cceip3_ob_out_pre.tdata [22]);
tran (kme_cceip3_ob_out_pre[21], \kme_cceip3_ob_out_pre.tdata [21]);
tran (kme_cceip3_ob_out_pre[20], \kme_cceip3_ob_out_pre.tdata [20]);
tran (kme_cceip3_ob_out_pre[19], \kme_cceip3_ob_out_pre.tdata [19]);
tran (kme_cceip3_ob_out_pre[18], \kme_cceip3_ob_out_pre.tdata [18]);
tran (kme_cceip3_ob_out_pre[17], \kme_cceip3_ob_out_pre.tdata [17]);
tran (kme_cceip3_ob_out_pre[16], \kme_cceip3_ob_out_pre.tdata [16]);
tran (kme_cceip3_ob_out_pre[15], \kme_cceip3_ob_out_pre.tdata [15]);
tran (kme_cceip3_ob_out_pre[14], \kme_cceip3_ob_out_pre.tdata [14]);
tran (kme_cceip3_ob_out_pre[13], \kme_cceip3_ob_out_pre.tdata [13]);
tran (kme_cceip3_ob_out_pre[12], \kme_cceip3_ob_out_pre.tdata [12]);
tran (kme_cceip3_ob_out_pre[11], \kme_cceip3_ob_out_pre.tdata [11]);
tran (kme_cceip3_ob_out_pre[10], \kme_cceip3_ob_out_pre.tdata [10]);
tran (kme_cceip3_ob_out_pre[9], \kme_cceip3_ob_out_pre.tdata [9]);
tran (kme_cceip3_ob_out_pre[8], \kme_cceip3_ob_out_pre.tdata [8]);
tran (kme_cceip3_ob_out_pre[7], \kme_cceip3_ob_out_pre.tdata [7]);
tran (kme_cceip3_ob_out_pre[6], \kme_cceip3_ob_out_pre.tdata [6]);
tran (kme_cceip3_ob_out_pre[5], \kme_cceip3_ob_out_pre.tdata [5]);
tran (kme_cceip3_ob_out_pre[4], \kme_cceip3_ob_out_pre.tdata [4]);
tran (kme_cceip3_ob_out_pre[3], \kme_cceip3_ob_out_pre.tdata [3]);
tran (kme_cceip3_ob_out_pre[2], \kme_cceip3_ob_out_pre.tdata [2]);
tran (kme_cceip3_ob_out_pre[1], \kme_cceip3_ob_out_pre.tdata [1]);
tran (kme_cceip3_ob_out_pre[0], \kme_cceip3_ob_out_pre.tdata [0]);
tran (kme_cceip3_ob_in[0], \kme_cceip3_ob_in.tready );
tran (kme_cddip0_ob_out_pre[82], \kme_cddip0_ob_out_pre.tvalid );
tran (kme_cddip0_ob_out_pre[81], \kme_cddip0_ob_out_pre.tlast );
tran (kme_cddip0_ob_out_pre[80], \kme_cddip0_ob_out_pre.tid [0]);
tran (kme_cddip0_ob_out_pre[79], \kme_cddip0_ob_out_pre.tstrb [7]);
tran (kme_cddip0_ob_out_pre[78], \kme_cddip0_ob_out_pre.tstrb [6]);
tran (kme_cddip0_ob_out_pre[77], \kme_cddip0_ob_out_pre.tstrb [5]);
tran (kme_cddip0_ob_out_pre[76], \kme_cddip0_ob_out_pre.tstrb [4]);
tran (kme_cddip0_ob_out_pre[75], \kme_cddip0_ob_out_pre.tstrb [3]);
tran (kme_cddip0_ob_out_pre[74], \kme_cddip0_ob_out_pre.tstrb [2]);
tran (kme_cddip0_ob_out_pre[73], \kme_cddip0_ob_out_pre.tstrb [1]);
tran (kme_cddip0_ob_out_pre[72], \kme_cddip0_ob_out_pre.tstrb [0]);
tran (kme_cddip0_ob_out_pre[71], \kme_cddip0_ob_out_pre.tuser [7]);
tran (kme_cddip0_ob_out_pre[70], \kme_cddip0_ob_out_pre.tuser [6]);
tran (kme_cddip0_ob_out_pre[69], \kme_cddip0_ob_out_pre.tuser [5]);
tran (kme_cddip0_ob_out_pre[68], \kme_cddip0_ob_out_pre.tuser [4]);
tran (kme_cddip0_ob_out_pre[67], \kme_cddip0_ob_out_pre.tuser [3]);
tran (kme_cddip0_ob_out_pre[66], \kme_cddip0_ob_out_pre.tuser [2]);
tran (kme_cddip0_ob_out_pre[65], \kme_cddip0_ob_out_pre.tuser [1]);
tran (kme_cddip0_ob_out_pre[64], \kme_cddip0_ob_out_pre.tuser [0]);
tran (kme_cddip0_ob_out_pre[63], \kme_cddip0_ob_out_pre.tdata [63]);
tran (kme_cddip0_ob_out_pre[62], \kme_cddip0_ob_out_pre.tdata [62]);
tran (kme_cddip0_ob_out_pre[61], \kme_cddip0_ob_out_pre.tdata [61]);
tran (kme_cddip0_ob_out_pre[60], \kme_cddip0_ob_out_pre.tdata [60]);
tran (kme_cddip0_ob_out_pre[59], \kme_cddip0_ob_out_pre.tdata [59]);
tran (kme_cddip0_ob_out_pre[58], \kme_cddip0_ob_out_pre.tdata [58]);
tran (kme_cddip0_ob_out_pre[57], \kme_cddip0_ob_out_pre.tdata [57]);
tran (kme_cddip0_ob_out_pre[56], \kme_cddip0_ob_out_pre.tdata [56]);
tran (kme_cddip0_ob_out_pre[55], \kme_cddip0_ob_out_pre.tdata [55]);
tran (kme_cddip0_ob_out_pre[54], \kme_cddip0_ob_out_pre.tdata [54]);
tran (kme_cddip0_ob_out_pre[53], \kme_cddip0_ob_out_pre.tdata [53]);
tran (kme_cddip0_ob_out_pre[52], \kme_cddip0_ob_out_pre.tdata [52]);
tran (kme_cddip0_ob_out_pre[51], \kme_cddip0_ob_out_pre.tdata [51]);
tran (kme_cddip0_ob_out_pre[50], \kme_cddip0_ob_out_pre.tdata [50]);
tran (kme_cddip0_ob_out_pre[49], \kme_cddip0_ob_out_pre.tdata [49]);
tran (kme_cddip0_ob_out_pre[48], \kme_cddip0_ob_out_pre.tdata [48]);
tran (kme_cddip0_ob_out_pre[47], \kme_cddip0_ob_out_pre.tdata [47]);
tran (kme_cddip0_ob_out_pre[46], \kme_cddip0_ob_out_pre.tdata [46]);
tran (kme_cddip0_ob_out_pre[45], \kme_cddip0_ob_out_pre.tdata [45]);
tran (kme_cddip0_ob_out_pre[44], \kme_cddip0_ob_out_pre.tdata [44]);
tran (kme_cddip0_ob_out_pre[43], \kme_cddip0_ob_out_pre.tdata [43]);
tran (kme_cddip0_ob_out_pre[42], \kme_cddip0_ob_out_pre.tdata [42]);
tran (kme_cddip0_ob_out_pre[41], \kme_cddip0_ob_out_pre.tdata [41]);
tran (kme_cddip0_ob_out_pre[40], \kme_cddip0_ob_out_pre.tdata [40]);
tran (kme_cddip0_ob_out_pre[39], \kme_cddip0_ob_out_pre.tdata [39]);
tran (kme_cddip0_ob_out_pre[38], \kme_cddip0_ob_out_pre.tdata [38]);
tran (kme_cddip0_ob_out_pre[37], \kme_cddip0_ob_out_pre.tdata [37]);
tran (kme_cddip0_ob_out_pre[36], \kme_cddip0_ob_out_pre.tdata [36]);
tran (kme_cddip0_ob_out_pre[35], \kme_cddip0_ob_out_pre.tdata [35]);
tran (kme_cddip0_ob_out_pre[34], \kme_cddip0_ob_out_pre.tdata [34]);
tran (kme_cddip0_ob_out_pre[33], \kme_cddip0_ob_out_pre.tdata [33]);
tran (kme_cddip0_ob_out_pre[32], \kme_cddip0_ob_out_pre.tdata [32]);
tran (kme_cddip0_ob_out_pre[31], \kme_cddip0_ob_out_pre.tdata [31]);
tran (kme_cddip0_ob_out_pre[30], \kme_cddip0_ob_out_pre.tdata [30]);
tran (kme_cddip0_ob_out_pre[29], \kme_cddip0_ob_out_pre.tdata [29]);
tran (kme_cddip0_ob_out_pre[28], \kme_cddip0_ob_out_pre.tdata [28]);
tran (kme_cddip0_ob_out_pre[27], \kme_cddip0_ob_out_pre.tdata [27]);
tran (kme_cddip0_ob_out_pre[26], \kme_cddip0_ob_out_pre.tdata [26]);
tran (kme_cddip0_ob_out_pre[25], \kme_cddip0_ob_out_pre.tdata [25]);
tran (kme_cddip0_ob_out_pre[24], \kme_cddip0_ob_out_pre.tdata [24]);
tran (kme_cddip0_ob_out_pre[23], \kme_cddip0_ob_out_pre.tdata [23]);
tran (kme_cddip0_ob_out_pre[22], \kme_cddip0_ob_out_pre.tdata [22]);
tran (kme_cddip0_ob_out_pre[21], \kme_cddip0_ob_out_pre.tdata [21]);
tran (kme_cddip0_ob_out_pre[20], \kme_cddip0_ob_out_pre.tdata [20]);
tran (kme_cddip0_ob_out_pre[19], \kme_cddip0_ob_out_pre.tdata [19]);
tran (kme_cddip0_ob_out_pre[18], \kme_cddip0_ob_out_pre.tdata [18]);
tran (kme_cddip0_ob_out_pre[17], \kme_cddip0_ob_out_pre.tdata [17]);
tran (kme_cddip0_ob_out_pre[16], \kme_cddip0_ob_out_pre.tdata [16]);
tran (kme_cddip0_ob_out_pre[15], \kme_cddip0_ob_out_pre.tdata [15]);
tran (kme_cddip0_ob_out_pre[14], \kme_cddip0_ob_out_pre.tdata [14]);
tran (kme_cddip0_ob_out_pre[13], \kme_cddip0_ob_out_pre.tdata [13]);
tran (kme_cddip0_ob_out_pre[12], \kme_cddip0_ob_out_pre.tdata [12]);
tran (kme_cddip0_ob_out_pre[11], \kme_cddip0_ob_out_pre.tdata [11]);
tran (kme_cddip0_ob_out_pre[10], \kme_cddip0_ob_out_pre.tdata [10]);
tran (kme_cddip0_ob_out_pre[9], \kme_cddip0_ob_out_pre.tdata [9]);
tran (kme_cddip0_ob_out_pre[8], \kme_cddip0_ob_out_pre.tdata [8]);
tran (kme_cddip0_ob_out_pre[7], \kme_cddip0_ob_out_pre.tdata [7]);
tran (kme_cddip0_ob_out_pre[6], \kme_cddip0_ob_out_pre.tdata [6]);
tran (kme_cddip0_ob_out_pre[5], \kme_cddip0_ob_out_pre.tdata [5]);
tran (kme_cddip0_ob_out_pre[4], \kme_cddip0_ob_out_pre.tdata [4]);
tran (kme_cddip0_ob_out_pre[3], \kme_cddip0_ob_out_pre.tdata [3]);
tran (kme_cddip0_ob_out_pre[2], \kme_cddip0_ob_out_pre.tdata [2]);
tran (kme_cddip0_ob_out_pre[1], \kme_cddip0_ob_out_pre.tdata [1]);
tran (kme_cddip0_ob_out_pre[0], \kme_cddip0_ob_out_pre.tdata [0]);
tran (kme_cddip0_ob_in[0], \kme_cddip0_ob_in.tready );
tran (kme_cddip1_ob_out_pre[82], \kme_cddip1_ob_out_pre.tvalid );
tran (kme_cddip1_ob_out_pre[81], \kme_cddip1_ob_out_pre.tlast );
tran (kme_cddip1_ob_out_pre[80], \kme_cddip1_ob_out_pre.tid [0]);
tran (kme_cddip1_ob_out_pre[79], \kme_cddip1_ob_out_pre.tstrb [7]);
tran (kme_cddip1_ob_out_pre[78], \kme_cddip1_ob_out_pre.tstrb [6]);
tran (kme_cddip1_ob_out_pre[77], \kme_cddip1_ob_out_pre.tstrb [5]);
tran (kme_cddip1_ob_out_pre[76], \kme_cddip1_ob_out_pre.tstrb [4]);
tran (kme_cddip1_ob_out_pre[75], \kme_cddip1_ob_out_pre.tstrb [3]);
tran (kme_cddip1_ob_out_pre[74], \kme_cddip1_ob_out_pre.tstrb [2]);
tran (kme_cddip1_ob_out_pre[73], \kme_cddip1_ob_out_pre.tstrb [1]);
tran (kme_cddip1_ob_out_pre[72], \kme_cddip1_ob_out_pre.tstrb [0]);
tran (kme_cddip1_ob_out_pre[71], \kme_cddip1_ob_out_pre.tuser [7]);
tran (kme_cddip1_ob_out_pre[70], \kme_cddip1_ob_out_pre.tuser [6]);
tran (kme_cddip1_ob_out_pre[69], \kme_cddip1_ob_out_pre.tuser [5]);
tran (kme_cddip1_ob_out_pre[68], \kme_cddip1_ob_out_pre.tuser [4]);
tran (kme_cddip1_ob_out_pre[67], \kme_cddip1_ob_out_pre.tuser [3]);
tran (kme_cddip1_ob_out_pre[66], \kme_cddip1_ob_out_pre.tuser [2]);
tran (kme_cddip1_ob_out_pre[65], \kme_cddip1_ob_out_pre.tuser [1]);
tran (kme_cddip1_ob_out_pre[64], \kme_cddip1_ob_out_pre.tuser [0]);
tran (kme_cddip1_ob_out_pre[63], \kme_cddip1_ob_out_pre.tdata [63]);
tran (kme_cddip1_ob_out_pre[62], \kme_cddip1_ob_out_pre.tdata [62]);
tran (kme_cddip1_ob_out_pre[61], \kme_cddip1_ob_out_pre.tdata [61]);
tran (kme_cddip1_ob_out_pre[60], \kme_cddip1_ob_out_pre.tdata [60]);
tran (kme_cddip1_ob_out_pre[59], \kme_cddip1_ob_out_pre.tdata [59]);
tran (kme_cddip1_ob_out_pre[58], \kme_cddip1_ob_out_pre.tdata [58]);
tran (kme_cddip1_ob_out_pre[57], \kme_cddip1_ob_out_pre.tdata [57]);
tran (kme_cddip1_ob_out_pre[56], \kme_cddip1_ob_out_pre.tdata [56]);
tran (kme_cddip1_ob_out_pre[55], \kme_cddip1_ob_out_pre.tdata [55]);
tran (kme_cddip1_ob_out_pre[54], \kme_cddip1_ob_out_pre.tdata [54]);
tran (kme_cddip1_ob_out_pre[53], \kme_cddip1_ob_out_pre.tdata [53]);
tran (kme_cddip1_ob_out_pre[52], \kme_cddip1_ob_out_pre.tdata [52]);
tran (kme_cddip1_ob_out_pre[51], \kme_cddip1_ob_out_pre.tdata [51]);
tran (kme_cddip1_ob_out_pre[50], \kme_cddip1_ob_out_pre.tdata [50]);
tran (kme_cddip1_ob_out_pre[49], \kme_cddip1_ob_out_pre.tdata [49]);
tran (kme_cddip1_ob_out_pre[48], \kme_cddip1_ob_out_pre.tdata [48]);
tran (kme_cddip1_ob_out_pre[47], \kme_cddip1_ob_out_pre.tdata [47]);
tran (kme_cddip1_ob_out_pre[46], \kme_cddip1_ob_out_pre.tdata [46]);
tran (kme_cddip1_ob_out_pre[45], \kme_cddip1_ob_out_pre.tdata [45]);
tran (kme_cddip1_ob_out_pre[44], \kme_cddip1_ob_out_pre.tdata [44]);
tran (kme_cddip1_ob_out_pre[43], \kme_cddip1_ob_out_pre.tdata [43]);
tran (kme_cddip1_ob_out_pre[42], \kme_cddip1_ob_out_pre.tdata [42]);
tran (kme_cddip1_ob_out_pre[41], \kme_cddip1_ob_out_pre.tdata [41]);
tran (kme_cddip1_ob_out_pre[40], \kme_cddip1_ob_out_pre.tdata [40]);
tran (kme_cddip1_ob_out_pre[39], \kme_cddip1_ob_out_pre.tdata [39]);
tran (kme_cddip1_ob_out_pre[38], \kme_cddip1_ob_out_pre.tdata [38]);
tran (kme_cddip1_ob_out_pre[37], \kme_cddip1_ob_out_pre.tdata [37]);
tran (kme_cddip1_ob_out_pre[36], \kme_cddip1_ob_out_pre.tdata [36]);
tran (kme_cddip1_ob_out_pre[35], \kme_cddip1_ob_out_pre.tdata [35]);
tran (kme_cddip1_ob_out_pre[34], \kme_cddip1_ob_out_pre.tdata [34]);
tran (kme_cddip1_ob_out_pre[33], \kme_cddip1_ob_out_pre.tdata [33]);
tran (kme_cddip1_ob_out_pre[32], \kme_cddip1_ob_out_pre.tdata [32]);
tran (kme_cddip1_ob_out_pre[31], \kme_cddip1_ob_out_pre.tdata [31]);
tran (kme_cddip1_ob_out_pre[30], \kme_cddip1_ob_out_pre.tdata [30]);
tran (kme_cddip1_ob_out_pre[29], \kme_cddip1_ob_out_pre.tdata [29]);
tran (kme_cddip1_ob_out_pre[28], \kme_cddip1_ob_out_pre.tdata [28]);
tran (kme_cddip1_ob_out_pre[27], \kme_cddip1_ob_out_pre.tdata [27]);
tran (kme_cddip1_ob_out_pre[26], \kme_cddip1_ob_out_pre.tdata [26]);
tran (kme_cddip1_ob_out_pre[25], \kme_cddip1_ob_out_pre.tdata [25]);
tran (kme_cddip1_ob_out_pre[24], \kme_cddip1_ob_out_pre.tdata [24]);
tran (kme_cddip1_ob_out_pre[23], \kme_cddip1_ob_out_pre.tdata [23]);
tran (kme_cddip1_ob_out_pre[22], \kme_cddip1_ob_out_pre.tdata [22]);
tran (kme_cddip1_ob_out_pre[21], \kme_cddip1_ob_out_pre.tdata [21]);
tran (kme_cddip1_ob_out_pre[20], \kme_cddip1_ob_out_pre.tdata [20]);
tran (kme_cddip1_ob_out_pre[19], \kme_cddip1_ob_out_pre.tdata [19]);
tran (kme_cddip1_ob_out_pre[18], \kme_cddip1_ob_out_pre.tdata [18]);
tran (kme_cddip1_ob_out_pre[17], \kme_cddip1_ob_out_pre.tdata [17]);
tran (kme_cddip1_ob_out_pre[16], \kme_cddip1_ob_out_pre.tdata [16]);
tran (kme_cddip1_ob_out_pre[15], \kme_cddip1_ob_out_pre.tdata [15]);
tran (kme_cddip1_ob_out_pre[14], \kme_cddip1_ob_out_pre.tdata [14]);
tran (kme_cddip1_ob_out_pre[13], \kme_cddip1_ob_out_pre.tdata [13]);
tran (kme_cddip1_ob_out_pre[12], \kme_cddip1_ob_out_pre.tdata [12]);
tran (kme_cddip1_ob_out_pre[11], \kme_cddip1_ob_out_pre.tdata [11]);
tran (kme_cddip1_ob_out_pre[10], \kme_cddip1_ob_out_pre.tdata [10]);
tran (kme_cddip1_ob_out_pre[9], \kme_cddip1_ob_out_pre.tdata [9]);
tran (kme_cddip1_ob_out_pre[8], \kme_cddip1_ob_out_pre.tdata [8]);
tran (kme_cddip1_ob_out_pre[7], \kme_cddip1_ob_out_pre.tdata [7]);
tran (kme_cddip1_ob_out_pre[6], \kme_cddip1_ob_out_pre.tdata [6]);
tran (kme_cddip1_ob_out_pre[5], \kme_cddip1_ob_out_pre.tdata [5]);
tran (kme_cddip1_ob_out_pre[4], \kme_cddip1_ob_out_pre.tdata [4]);
tran (kme_cddip1_ob_out_pre[3], \kme_cddip1_ob_out_pre.tdata [3]);
tran (kme_cddip1_ob_out_pre[2], \kme_cddip1_ob_out_pre.tdata [2]);
tran (kme_cddip1_ob_out_pre[1], \kme_cddip1_ob_out_pre.tdata [1]);
tran (kme_cddip1_ob_out_pre[0], \kme_cddip1_ob_out_pre.tdata [0]);
tran (kme_cddip1_ob_in[0], \kme_cddip1_ob_in.tready );
tran (kme_cddip2_ob_out_pre[82], \kme_cddip2_ob_out_pre.tvalid );
tran (kme_cddip2_ob_out_pre[81], \kme_cddip2_ob_out_pre.tlast );
tran (kme_cddip2_ob_out_pre[80], \kme_cddip2_ob_out_pre.tid [0]);
tran (kme_cddip2_ob_out_pre[79], \kme_cddip2_ob_out_pre.tstrb [7]);
tran (kme_cddip2_ob_out_pre[78], \kme_cddip2_ob_out_pre.tstrb [6]);
tran (kme_cddip2_ob_out_pre[77], \kme_cddip2_ob_out_pre.tstrb [5]);
tran (kme_cddip2_ob_out_pre[76], \kme_cddip2_ob_out_pre.tstrb [4]);
tran (kme_cddip2_ob_out_pre[75], \kme_cddip2_ob_out_pre.tstrb [3]);
tran (kme_cddip2_ob_out_pre[74], \kme_cddip2_ob_out_pre.tstrb [2]);
tran (kme_cddip2_ob_out_pre[73], \kme_cddip2_ob_out_pre.tstrb [1]);
tran (kme_cddip2_ob_out_pre[72], \kme_cddip2_ob_out_pre.tstrb [0]);
tran (kme_cddip2_ob_out_pre[71], \kme_cddip2_ob_out_pre.tuser [7]);
tran (kme_cddip2_ob_out_pre[70], \kme_cddip2_ob_out_pre.tuser [6]);
tran (kme_cddip2_ob_out_pre[69], \kme_cddip2_ob_out_pre.tuser [5]);
tran (kme_cddip2_ob_out_pre[68], \kme_cddip2_ob_out_pre.tuser [4]);
tran (kme_cddip2_ob_out_pre[67], \kme_cddip2_ob_out_pre.tuser [3]);
tran (kme_cddip2_ob_out_pre[66], \kme_cddip2_ob_out_pre.tuser [2]);
tran (kme_cddip2_ob_out_pre[65], \kme_cddip2_ob_out_pre.tuser [1]);
tran (kme_cddip2_ob_out_pre[64], \kme_cddip2_ob_out_pre.tuser [0]);
tran (kme_cddip2_ob_out_pre[63], \kme_cddip2_ob_out_pre.tdata [63]);
tran (kme_cddip2_ob_out_pre[62], \kme_cddip2_ob_out_pre.tdata [62]);
tran (kme_cddip2_ob_out_pre[61], \kme_cddip2_ob_out_pre.tdata [61]);
tran (kme_cddip2_ob_out_pre[60], \kme_cddip2_ob_out_pre.tdata [60]);
tran (kme_cddip2_ob_out_pre[59], \kme_cddip2_ob_out_pre.tdata [59]);
tran (kme_cddip2_ob_out_pre[58], \kme_cddip2_ob_out_pre.tdata [58]);
tran (kme_cddip2_ob_out_pre[57], \kme_cddip2_ob_out_pre.tdata [57]);
tran (kme_cddip2_ob_out_pre[56], \kme_cddip2_ob_out_pre.tdata [56]);
tran (kme_cddip2_ob_out_pre[55], \kme_cddip2_ob_out_pre.tdata [55]);
tran (kme_cddip2_ob_out_pre[54], \kme_cddip2_ob_out_pre.tdata [54]);
tran (kme_cddip2_ob_out_pre[53], \kme_cddip2_ob_out_pre.tdata [53]);
tran (kme_cddip2_ob_out_pre[52], \kme_cddip2_ob_out_pre.tdata [52]);
tran (kme_cddip2_ob_out_pre[51], \kme_cddip2_ob_out_pre.tdata [51]);
tran (kme_cddip2_ob_out_pre[50], \kme_cddip2_ob_out_pre.tdata [50]);
tran (kme_cddip2_ob_out_pre[49], \kme_cddip2_ob_out_pre.tdata [49]);
tran (kme_cddip2_ob_out_pre[48], \kme_cddip2_ob_out_pre.tdata [48]);
tran (kme_cddip2_ob_out_pre[47], \kme_cddip2_ob_out_pre.tdata [47]);
tran (kme_cddip2_ob_out_pre[46], \kme_cddip2_ob_out_pre.tdata [46]);
tran (kme_cddip2_ob_out_pre[45], \kme_cddip2_ob_out_pre.tdata [45]);
tran (kme_cddip2_ob_out_pre[44], \kme_cddip2_ob_out_pre.tdata [44]);
tran (kme_cddip2_ob_out_pre[43], \kme_cddip2_ob_out_pre.tdata [43]);
tran (kme_cddip2_ob_out_pre[42], \kme_cddip2_ob_out_pre.tdata [42]);
tran (kme_cddip2_ob_out_pre[41], \kme_cddip2_ob_out_pre.tdata [41]);
tran (kme_cddip2_ob_out_pre[40], \kme_cddip2_ob_out_pre.tdata [40]);
tran (kme_cddip2_ob_out_pre[39], \kme_cddip2_ob_out_pre.tdata [39]);
tran (kme_cddip2_ob_out_pre[38], \kme_cddip2_ob_out_pre.tdata [38]);
tran (kme_cddip2_ob_out_pre[37], \kme_cddip2_ob_out_pre.tdata [37]);
tran (kme_cddip2_ob_out_pre[36], \kme_cddip2_ob_out_pre.tdata [36]);
tran (kme_cddip2_ob_out_pre[35], \kme_cddip2_ob_out_pre.tdata [35]);
tran (kme_cddip2_ob_out_pre[34], \kme_cddip2_ob_out_pre.tdata [34]);
tran (kme_cddip2_ob_out_pre[33], \kme_cddip2_ob_out_pre.tdata [33]);
tran (kme_cddip2_ob_out_pre[32], \kme_cddip2_ob_out_pre.tdata [32]);
tran (kme_cddip2_ob_out_pre[31], \kme_cddip2_ob_out_pre.tdata [31]);
tran (kme_cddip2_ob_out_pre[30], \kme_cddip2_ob_out_pre.tdata [30]);
tran (kme_cddip2_ob_out_pre[29], \kme_cddip2_ob_out_pre.tdata [29]);
tran (kme_cddip2_ob_out_pre[28], \kme_cddip2_ob_out_pre.tdata [28]);
tran (kme_cddip2_ob_out_pre[27], \kme_cddip2_ob_out_pre.tdata [27]);
tran (kme_cddip2_ob_out_pre[26], \kme_cddip2_ob_out_pre.tdata [26]);
tran (kme_cddip2_ob_out_pre[25], \kme_cddip2_ob_out_pre.tdata [25]);
tran (kme_cddip2_ob_out_pre[24], \kme_cddip2_ob_out_pre.tdata [24]);
tran (kme_cddip2_ob_out_pre[23], \kme_cddip2_ob_out_pre.tdata [23]);
tran (kme_cddip2_ob_out_pre[22], \kme_cddip2_ob_out_pre.tdata [22]);
tran (kme_cddip2_ob_out_pre[21], \kme_cddip2_ob_out_pre.tdata [21]);
tran (kme_cddip2_ob_out_pre[20], \kme_cddip2_ob_out_pre.tdata [20]);
tran (kme_cddip2_ob_out_pre[19], \kme_cddip2_ob_out_pre.tdata [19]);
tran (kme_cddip2_ob_out_pre[18], \kme_cddip2_ob_out_pre.tdata [18]);
tran (kme_cddip2_ob_out_pre[17], \kme_cddip2_ob_out_pre.tdata [17]);
tran (kme_cddip2_ob_out_pre[16], \kme_cddip2_ob_out_pre.tdata [16]);
tran (kme_cddip2_ob_out_pre[15], \kme_cddip2_ob_out_pre.tdata [15]);
tran (kme_cddip2_ob_out_pre[14], \kme_cddip2_ob_out_pre.tdata [14]);
tran (kme_cddip2_ob_out_pre[13], \kme_cddip2_ob_out_pre.tdata [13]);
tran (kme_cddip2_ob_out_pre[12], \kme_cddip2_ob_out_pre.tdata [12]);
tran (kme_cddip2_ob_out_pre[11], \kme_cddip2_ob_out_pre.tdata [11]);
tran (kme_cddip2_ob_out_pre[10], \kme_cddip2_ob_out_pre.tdata [10]);
tran (kme_cddip2_ob_out_pre[9], \kme_cddip2_ob_out_pre.tdata [9]);
tran (kme_cddip2_ob_out_pre[8], \kme_cddip2_ob_out_pre.tdata [8]);
tran (kme_cddip2_ob_out_pre[7], \kme_cddip2_ob_out_pre.tdata [7]);
tran (kme_cddip2_ob_out_pre[6], \kme_cddip2_ob_out_pre.tdata [6]);
tran (kme_cddip2_ob_out_pre[5], \kme_cddip2_ob_out_pre.tdata [5]);
tran (kme_cddip2_ob_out_pre[4], \kme_cddip2_ob_out_pre.tdata [4]);
tran (kme_cddip2_ob_out_pre[3], \kme_cddip2_ob_out_pre.tdata [3]);
tran (kme_cddip2_ob_out_pre[2], \kme_cddip2_ob_out_pre.tdata [2]);
tran (kme_cddip2_ob_out_pre[1], \kme_cddip2_ob_out_pre.tdata [1]);
tran (kme_cddip2_ob_out_pre[0], \kme_cddip2_ob_out_pre.tdata [0]);
tran (kme_cddip2_ob_in[0], \kme_cddip2_ob_in.tready );
tran (kme_cddip3_ob_out_pre[82], \kme_cddip3_ob_out_pre.tvalid );
tran (kme_cddip3_ob_out_pre[81], \kme_cddip3_ob_out_pre.tlast );
tran (kme_cddip3_ob_out_pre[80], \kme_cddip3_ob_out_pre.tid [0]);
tran (kme_cddip3_ob_out_pre[79], \kme_cddip3_ob_out_pre.tstrb [7]);
tran (kme_cddip3_ob_out_pre[78], \kme_cddip3_ob_out_pre.tstrb [6]);
tran (kme_cddip3_ob_out_pre[77], \kme_cddip3_ob_out_pre.tstrb [5]);
tran (kme_cddip3_ob_out_pre[76], \kme_cddip3_ob_out_pre.tstrb [4]);
tran (kme_cddip3_ob_out_pre[75], \kme_cddip3_ob_out_pre.tstrb [3]);
tran (kme_cddip3_ob_out_pre[74], \kme_cddip3_ob_out_pre.tstrb [2]);
tran (kme_cddip3_ob_out_pre[73], \kme_cddip3_ob_out_pre.tstrb [1]);
tran (kme_cddip3_ob_out_pre[72], \kme_cddip3_ob_out_pre.tstrb [0]);
tran (kme_cddip3_ob_out_pre[71], \kme_cddip3_ob_out_pre.tuser [7]);
tran (kme_cddip3_ob_out_pre[70], \kme_cddip3_ob_out_pre.tuser [6]);
tran (kme_cddip3_ob_out_pre[69], \kme_cddip3_ob_out_pre.tuser [5]);
tran (kme_cddip3_ob_out_pre[68], \kme_cddip3_ob_out_pre.tuser [4]);
tran (kme_cddip3_ob_out_pre[67], \kme_cddip3_ob_out_pre.tuser [3]);
tran (kme_cddip3_ob_out_pre[66], \kme_cddip3_ob_out_pre.tuser [2]);
tran (kme_cddip3_ob_out_pre[65], \kme_cddip3_ob_out_pre.tuser [1]);
tran (kme_cddip3_ob_out_pre[64], \kme_cddip3_ob_out_pre.tuser [0]);
tran (kme_cddip3_ob_out_pre[63], \kme_cddip3_ob_out_pre.tdata [63]);
tran (kme_cddip3_ob_out_pre[62], \kme_cddip3_ob_out_pre.tdata [62]);
tran (kme_cddip3_ob_out_pre[61], \kme_cddip3_ob_out_pre.tdata [61]);
tran (kme_cddip3_ob_out_pre[60], \kme_cddip3_ob_out_pre.tdata [60]);
tran (kme_cddip3_ob_out_pre[59], \kme_cddip3_ob_out_pre.tdata [59]);
tran (kme_cddip3_ob_out_pre[58], \kme_cddip3_ob_out_pre.tdata [58]);
tran (kme_cddip3_ob_out_pre[57], \kme_cddip3_ob_out_pre.tdata [57]);
tran (kme_cddip3_ob_out_pre[56], \kme_cddip3_ob_out_pre.tdata [56]);
tran (kme_cddip3_ob_out_pre[55], \kme_cddip3_ob_out_pre.tdata [55]);
tran (kme_cddip3_ob_out_pre[54], \kme_cddip3_ob_out_pre.tdata [54]);
tran (kme_cddip3_ob_out_pre[53], \kme_cddip3_ob_out_pre.tdata [53]);
tran (kme_cddip3_ob_out_pre[52], \kme_cddip3_ob_out_pre.tdata [52]);
tran (kme_cddip3_ob_out_pre[51], \kme_cddip3_ob_out_pre.tdata [51]);
tran (kme_cddip3_ob_out_pre[50], \kme_cddip3_ob_out_pre.tdata [50]);
tran (kme_cddip3_ob_out_pre[49], \kme_cddip3_ob_out_pre.tdata [49]);
tran (kme_cddip3_ob_out_pre[48], \kme_cddip3_ob_out_pre.tdata [48]);
tran (kme_cddip3_ob_out_pre[47], \kme_cddip3_ob_out_pre.tdata [47]);
tran (kme_cddip3_ob_out_pre[46], \kme_cddip3_ob_out_pre.tdata [46]);
tran (kme_cddip3_ob_out_pre[45], \kme_cddip3_ob_out_pre.tdata [45]);
tran (kme_cddip3_ob_out_pre[44], \kme_cddip3_ob_out_pre.tdata [44]);
tran (kme_cddip3_ob_out_pre[43], \kme_cddip3_ob_out_pre.tdata [43]);
tran (kme_cddip3_ob_out_pre[42], \kme_cddip3_ob_out_pre.tdata [42]);
tran (kme_cddip3_ob_out_pre[41], \kme_cddip3_ob_out_pre.tdata [41]);
tran (kme_cddip3_ob_out_pre[40], \kme_cddip3_ob_out_pre.tdata [40]);
tran (kme_cddip3_ob_out_pre[39], \kme_cddip3_ob_out_pre.tdata [39]);
tran (kme_cddip3_ob_out_pre[38], \kme_cddip3_ob_out_pre.tdata [38]);
tran (kme_cddip3_ob_out_pre[37], \kme_cddip3_ob_out_pre.tdata [37]);
tran (kme_cddip3_ob_out_pre[36], \kme_cddip3_ob_out_pre.tdata [36]);
tran (kme_cddip3_ob_out_pre[35], \kme_cddip3_ob_out_pre.tdata [35]);
tran (kme_cddip3_ob_out_pre[34], \kme_cddip3_ob_out_pre.tdata [34]);
tran (kme_cddip3_ob_out_pre[33], \kme_cddip3_ob_out_pre.tdata [33]);
tran (kme_cddip3_ob_out_pre[32], \kme_cddip3_ob_out_pre.tdata [32]);
tran (kme_cddip3_ob_out_pre[31], \kme_cddip3_ob_out_pre.tdata [31]);
tran (kme_cddip3_ob_out_pre[30], \kme_cddip3_ob_out_pre.tdata [30]);
tran (kme_cddip3_ob_out_pre[29], \kme_cddip3_ob_out_pre.tdata [29]);
tran (kme_cddip3_ob_out_pre[28], \kme_cddip3_ob_out_pre.tdata [28]);
tran (kme_cddip3_ob_out_pre[27], \kme_cddip3_ob_out_pre.tdata [27]);
tran (kme_cddip3_ob_out_pre[26], \kme_cddip3_ob_out_pre.tdata [26]);
tran (kme_cddip3_ob_out_pre[25], \kme_cddip3_ob_out_pre.tdata [25]);
tran (kme_cddip3_ob_out_pre[24], \kme_cddip3_ob_out_pre.tdata [24]);
tran (kme_cddip3_ob_out_pre[23], \kme_cddip3_ob_out_pre.tdata [23]);
tran (kme_cddip3_ob_out_pre[22], \kme_cddip3_ob_out_pre.tdata [22]);
tran (kme_cddip3_ob_out_pre[21], \kme_cddip3_ob_out_pre.tdata [21]);
tran (kme_cddip3_ob_out_pre[20], \kme_cddip3_ob_out_pre.tdata [20]);
tran (kme_cddip3_ob_out_pre[19], \kme_cddip3_ob_out_pre.tdata [19]);
tran (kme_cddip3_ob_out_pre[18], \kme_cddip3_ob_out_pre.tdata [18]);
tran (kme_cddip3_ob_out_pre[17], \kme_cddip3_ob_out_pre.tdata [17]);
tran (kme_cddip3_ob_out_pre[16], \kme_cddip3_ob_out_pre.tdata [16]);
tran (kme_cddip3_ob_out_pre[15], \kme_cddip3_ob_out_pre.tdata [15]);
tran (kme_cddip3_ob_out_pre[14], \kme_cddip3_ob_out_pre.tdata [14]);
tran (kme_cddip3_ob_out_pre[13], \kme_cddip3_ob_out_pre.tdata [13]);
tran (kme_cddip3_ob_out_pre[12], \kme_cddip3_ob_out_pre.tdata [12]);
tran (kme_cddip3_ob_out_pre[11], \kme_cddip3_ob_out_pre.tdata [11]);
tran (kme_cddip3_ob_out_pre[10], \kme_cddip3_ob_out_pre.tdata [10]);
tran (kme_cddip3_ob_out_pre[9], \kme_cddip3_ob_out_pre.tdata [9]);
tran (kme_cddip3_ob_out_pre[8], \kme_cddip3_ob_out_pre.tdata [8]);
tran (kme_cddip3_ob_out_pre[7], \kme_cddip3_ob_out_pre.tdata [7]);
tran (kme_cddip3_ob_out_pre[6], \kme_cddip3_ob_out_pre.tdata [6]);
tran (kme_cddip3_ob_out_pre[5], \kme_cddip3_ob_out_pre.tdata [5]);
tran (kme_cddip3_ob_out_pre[4], \kme_cddip3_ob_out_pre.tdata [4]);
tran (kme_cddip3_ob_out_pre[3], \kme_cddip3_ob_out_pre.tdata [3]);
tran (kme_cddip3_ob_out_pre[2], \kme_cddip3_ob_out_pre.tdata [2]);
tran (kme_cddip3_ob_out_pre[1], \kme_cddip3_ob_out_pre.tdata [1]);
tran (kme_cddip3_ob_out_pre[0], \kme_cddip3_ob_out_pre.tdata [0]);
tran (kme_cddip3_ob_in[0], \kme_cddip3_ob_in.tready );
tran (idle_components[31], \idle_components.r.part0 [31]);
tran (idle_components[31], \idle_components.f.num_key_tlvs_in_flight [19]);
tran (idle_components[30], \idle_components.r.part0 [30]);
tran (idle_components[30], \idle_components.f.num_key_tlvs_in_flight [18]);
tran (idle_components[29], \idle_components.r.part0 [29]);
tran (idle_components[29], \idle_components.f.num_key_tlvs_in_flight [17]);
tran (idle_components[28], \idle_components.r.part0 [28]);
tran (idle_components[28], \idle_components.f.num_key_tlvs_in_flight [16]);
tran (idle_components[27], \idle_components.r.part0 [27]);
tran (idle_components[27], \idle_components.f.num_key_tlvs_in_flight [15]);
tran (idle_components[26], \idle_components.r.part0 [26]);
tran (idle_components[26], \idle_components.f.num_key_tlvs_in_flight [14]);
tran (idle_components[25], \idle_components.r.part0 [25]);
tran (idle_components[25], \idle_components.f.num_key_tlvs_in_flight [13]);
tran (idle_components[24], \idle_components.r.part0 [24]);
tran (idle_components[24], \idle_components.f.num_key_tlvs_in_flight [12]);
tran (idle_components[23], \idle_components.r.part0 [23]);
tran (idle_components[23], \idle_components.f.num_key_tlvs_in_flight [11]);
tran (idle_components[22], \idle_components.r.part0 [22]);
tran (idle_components[22], \idle_components.f.num_key_tlvs_in_flight [10]);
tran (idle_components[21], \idle_components.r.part0 [21]);
tran (idle_components[21], \idle_components.f.num_key_tlvs_in_flight [9]);
tran (idle_components[20], \idle_components.r.part0 [20]);
tran (idle_components[20], \idle_components.f.num_key_tlvs_in_flight [8]);
tran (idle_components[19], \idle_components.r.part0 [19]);
tran (idle_components[19], \idle_components.f.num_key_tlvs_in_flight [7]);
tran (idle_components[18], \idle_components.r.part0 [18]);
tran (idle_components[18], \idle_components.f.num_key_tlvs_in_flight [6]);
tran (idle_components[17], \idle_components.r.part0 [17]);
tran (idle_components[17], \idle_components.f.num_key_tlvs_in_flight [5]);
tran (idle_components[16], \idle_components.r.part0 [16]);
tran (idle_components[16], \idle_components.f.num_key_tlvs_in_flight [4]);
tran (idle_components[15], \idle_components.r.part0 [15]);
tran (idle_components[15], \idle_components.f.num_key_tlvs_in_flight [3]);
tran (idle_components[14], \idle_components.r.part0 [14]);
tran (idle_components[14], \idle_components.f.num_key_tlvs_in_flight [2]);
tran (idle_components[13], \idle_components.r.part0 [13]);
tran (idle_components[13], \idle_components.f.num_key_tlvs_in_flight [1]);
tran (idle_components[12], \idle_components.r.part0 [12]);
tran (idle_components[12], \idle_components.f.num_key_tlvs_in_flight [0]);
tran (idle_components[11], \idle_components.r.part0 [11]);
tran (idle_components[11], \idle_components.f.cddip0_key_tlv_rsm_idle );
tran (idle_components[10], \idle_components.r.part0 [10]);
tran (idle_components[10], \idle_components.f.cddip1_key_tlv_rsm_idle );
tran (idle_components[9], \idle_components.r.part0 [9]);
tran (idle_components[9], \idle_components.f.cddip2_key_tlv_rsm_idle );
tran (idle_components[8], \idle_components.r.part0 [8]);
tran (idle_components[8], \idle_components.f.cddip3_key_tlv_rsm_idle );
tran (idle_components[7], \idle_components.r.part0 [7]);
tran (idle_components[7], \idle_components.f.cceip0_key_tlv_rsm_idle );
tran (idle_components[6], \idle_components.r.part0 [6]);
tran (idle_components[6], \idle_components.f.cceip1_key_tlv_rsm_idle );
tran (idle_components[5], \idle_components.r.part0 [5]);
tran (idle_components[5], \idle_components.f.cceip2_key_tlv_rsm_idle );
tran (idle_components[4], \idle_components.r.part0 [4]);
tran (idle_components[4], \idle_components.f.cceip3_key_tlv_rsm_idle );
tran (idle_components[3], \idle_components.r.part0 [3]);
tran (idle_components[3], \idle_components.f.no_key_tlv_in_flight );
tran (idle_components[2], \idle_components.r.part0 [2]);
tran (idle_components[2], \idle_components.f.tlv_parser_idle );
tran (idle_components[1], \idle_components.r.part0 [1]);
tran (idle_components[1], \idle_components.f.drng_idle );
tran (idle_components[0], \idle_components.r.part0 [0]);
tran (idle_components[0], \idle_components.f.kme_slv_empty );
tran (\sa_snapshot[0][0] , \sa_snapshot[0].r.part0[0] );
tran (\sa_snapshot[0][0] , \sa_snapshot[0].f.lower[0] );
tran (\sa_snapshot[0][1] , \sa_snapshot[0].r.part0[1] );
tran (\sa_snapshot[0][1] , \sa_snapshot[0].f.lower[1] );
tran (\sa_snapshot[0][2] , \sa_snapshot[0].r.part0[2] );
tran (\sa_snapshot[0][2] , \sa_snapshot[0].f.lower[2] );
tran (\sa_snapshot[0][3] , \sa_snapshot[0].r.part0[3] );
tran (\sa_snapshot[0][3] , \sa_snapshot[0].f.lower[3] );
tran (\sa_snapshot[0][4] , \sa_snapshot[0].r.part0[4] );
tran (\sa_snapshot[0][4] , \sa_snapshot[0].f.lower[4] );
tran (\sa_snapshot[0][5] , \sa_snapshot[0].r.part0[5] );
tran (\sa_snapshot[0][5] , \sa_snapshot[0].f.lower[5] );
tran (\sa_snapshot[0][6] , \sa_snapshot[0].r.part0[6] );
tran (\sa_snapshot[0][6] , \sa_snapshot[0].f.lower[6] );
tran (\sa_snapshot[0][7] , \sa_snapshot[0].r.part0[7] );
tran (\sa_snapshot[0][7] , \sa_snapshot[0].f.lower[7] );
tran (\sa_snapshot[0][8] , \sa_snapshot[0].r.part0[8] );
tran (\sa_snapshot[0][8] , \sa_snapshot[0].f.lower[8] );
tran (\sa_snapshot[0][9] , \sa_snapshot[0].r.part0[9] );
tran (\sa_snapshot[0][9] , \sa_snapshot[0].f.lower[9] );
tran (\sa_snapshot[0][10] , \sa_snapshot[0].r.part0[10] );
tran (\sa_snapshot[0][10] , \sa_snapshot[0].f.lower[10] );
tran (\sa_snapshot[0][11] , \sa_snapshot[0].r.part0[11] );
tran (\sa_snapshot[0][11] , \sa_snapshot[0].f.lower[11] );
tran (\sa_snapshot[0][12] , \sa_snapshot[0].r.part0[12] );
tran (\sa_snapshot[0][12] , \sa_snapshot[0].f.lower[12] );
tran (\sa_snapshot[0][13] , \sa_snapshot[0].r.part0[13] );
tran (\sa_snapshot[0][13] , \sa_snapshot[0].f.lower[13] );
tran (\sa_snapshot[0][14] , \sa_snapshot[0].r.part0[14] );
tran (\sa_snapshot[0][14] , \sa_snapshot[0].f.lower[14] );
tran (\sa_snapshot[0][15] , \sa_snapshot[0].r.part0[15] );
tran (\sa_snapshot[0][15] , \sa_snapshot[0].f.lower[15] );
tran (\sa_snapshot[0][16] , \sa_snapshot[0].r.part0[16] );
tran (\sa_snapshot[0][16] , \sa_snapshot[0].f.lower[16] );
tran (\sa_snapshot[0][17] , \sa_snapshot[0].r.part0[17] );
tran (\sa_snapshot[0][17] , \sa_snapshot[0].f.lower[17] );
tran (\sa_snapshot[0][18] , \sa_snapshot[0].r.part0[18] );
tran (\sa_snapshot[0][18] , \sa_snapshot[0].f.lower[18] );
tran (\sa_snapshot[0][19] , \sa_snapshot[0].r.part0[19] );
tran (\sa_snapshot[0][19] , \sa_snapshot[0].f.lower[19] );
tran (\sa_snapshot[0][20] , \sa_snapshot[0].r.part0[20] );
tran (\sa_snapshot[0][20] , \sa_snapshot[0].f.lower[20] );
tran (\sa_snapshot[0][21] , \sa_snapshot[0].r.part0[21] );
tran (\sa_snapshot[0][21] , \sa_snapshot[0].f.lower[21] );
tran (\sa_snapshot[0][22] , \sa_snapshot[0].r.part0[22] );
tran (\sa_snapshot[0][22] , \sa_snapshot[0].f.lower[22] );
tran (\sa_snapshot[0][23] , \sa_snapshot[0].r.part0[23] );
tran (\sa_snapshot[0][23] , \sa_snapshot[0].f.lower[23] );
tran (\sa_snapshot[0][24] , \sa_snapshot[0].r.part0[24] );
tran (\sa_snapshot[0][24] , \sa_snapshot[0].f.lower[24] );
tran (\sa_snapshot[0][25] , \sa_snapshot[0].r.part0[25] );
tran (\sa_snapshot[0][25] , \sa_snapshot[0].f.lower[25] );
tran (\sa_snapshot[0][26] , \sa_snapshot[0].r.part0[26] );
tran (\sa_snapshot[0][26] , \sa_snapshot[0].f.lower[26] );
tran (\sa_snapshot[0][27] , \sa_snapshot[0].r.part0[27] );
tran (\sa_snapshot[0][27] , \sa_snapshot[0].f.lower[27] );
tran (\sa_snapshot[0][28] , \sa_snapshot[0].r.part0[28] );
tran (\sa_snapshot[0][28] , \sa_snapshot[0].f.lower[28] );
tran (\sa_snapshot[0][29] , \sa_snapshot[0].r.part0[29] );
tran (\sa_snapshot[0][29] , \sa_snapshot[0].f.lower[29] );
tran (\sa_snapshot[0][30] , \sa_snapshot[0].r.part0[30] );
tran (\sa_snapshot[0][30] , \sa_snapshot[0].f.lower[30] );
tran (\sa_snapshot[0][31] , \sa_snapshot[0].r.part0[31] );
tran (\sa_snapshot[0][31] , \sa_snapshot[0].f.lower[31] );
tran (\sa_snapshot[0][32] , \sa_snapshot[0].r.part1[0] );
tran (\sa_snapshot[0][32] , \sa_snapshot[0].f.upper[0] );
tran (\sa_snapshot[0][33] , \sa_snapshot[0].r.part1[1] );
tran (\sa_snapshot[0][33] , \sa_snapshot[0].f.upper[1] );
tran (\sa_snapshot[0][34] , \sa_snapshot[0].r.part1[2] );
tran (\sa_snapshot[0][34] , \sa_snapshot[0].f.upper[2] );
tran (\sa_snapshot[0][35] , \sa_snapshot[0].r.part1[3] );
tran (\sa_snapshot[0][35] , \sa_snapshot[0].f.upper[3] );
tran (\sa_snapshot[0][36] , \sa_snapshot[0].r.part1[4] );
tran (\sa_snapshot[0][36] , \sa_snapshot[0].f.upper[4] );
tran (\sa_snapshot[0][37] , \sa_snapshot[0].r.part1[5] );
tran (\sa_snapshot[0][37] , \sa_snapshot[0].f.upper[5] );
tran (\sa_snapshot[0][38] , \sa_snapshot[0].r.part1[6] );
tran (\sa_snapshot[0][38] , \sa_snapshot[0].f.upper[6] );
tran (\sa_snapshot[0][39] , \sa_snapshot[0].r.part1[7] );
tran (\sa_snapshot[0][39] , \sa_snapshot[0].f.upper[7] );
tran (\sa_snapshot[0][40] , \sa_snapshot[0].r.part1[8] );
tran (\sa_snapshot[0][40] , \sa_snapshot[0].f.upper[8] );
tran (\sa_snapshot[0][41] , \sa_snapshot[0].r.part1[9] );
tran (\sa_snapshot[0][41] , \sa_snapshot[0].f.upper[9] );
tran (\sa_snapshot[0][42] , \sa_snapshot[0].r.part1[10] );
tran (\sa_snapshot[0][42] , \sa_snapshot[0].f.upper[10] );
tran (\sa_snapshot[0][43] , \sa_snapshot[0].r.part1[11] );
tran (\sa_snapshot[0][43] , \sa_snapshot[0].f.upper[11] );
tran (\sa_snapshot[0][44] , \sa_snapshot[0].r.part1[12] );
tran (\sa_snapshot[0][44] , \sa_snapshot[0].f.upper[12] );
tran (\sa_snapshot[0][45] , \sa_snapshot[0].r.part1[13] );
tran (\sa_snapshot[0][45] , \sa_snapshot[0].f.upper[13] );
tran (\sa_snapshot[0][46] , \sa_snapshot[0].r.part1[14] );
tran (\sa_snapshot[0][46] , \sa_snapshot[0].f.upper[14] );
tran (\sa_snapshot[0][47] , \sa_snapshot[0].r.part1[15] );
tran (\sa_snapshot[0][47] , \sa_snapshot[0].f.upper[15] );
tran (\sa_snapshot[0][48] , \sa_snapshot[0].r.part1[16] );
tran (\sa_snapshot[0][48] , \sa_snapshot[0].f.upper[16] );
tran (\sa_snapshot[0][49] , \sa_snapshot[0].r.part1[17] );
tran (\sa_snapshot[0][49] , \sa_snapshot[0].f.upper[17] );
tran (\sa_snapshot[0][50] , \sa_snapshot[0].r.part1[18] );
tran (\sa_snapshot[0][50] , \sa_snapshot[0].f.unused[0] );
tran (\sa_snapshot[0][51] , \sa_snapshot[0].r.part1[19] );
tran (\sa_snapshot[0][51] , \sa_snapshot[0].f.unused[1] );
tran (\sa_snapshot[0][52] , \sa_snapshot[0].r.part1[20] );
tran (\sa_snapshot[0][52] , \sa_snapshot[0].f.unused[2] );
tran (\sa_snapshot[0][53] , \sa_snapshot[0].r.part1[21] );
tran (\sa_snapshot[0][53] , \sa_snapshot[0].f.unused[3] );
tran (\sa_snapshot[0][54] , \sa_snapshot[0].r.part1[22] );
tran (\sa_snapshot[0][54] , \sa_snapshot[0].f.unused[4] );
tran (\sa_snapshot[0][55] , \sa_snapshot[0].r.part1[23] );
tran (\sa_snapshot[0][55] , \sa_snapshot[0].f.unused[5] );
tran (\sa_snapshot[0][56] , \sa_snapshot[0].r.part1[24] );
tran (\sa_snapshot[0][56] , \sa_snapshot[0].f.unused[6] );
tran (\sa_snapshot[0][57] , \sa_snapshot[0].r.part1[25] );
tran (\sa_snapshot[0][57] , \sa_snapshot[0].f.unused[7] );
tran (\sa_snapshot[0][58] , \sa_snapshot[0].r.part1[26] );
tran (\sa_snapshot[0][58] , \sa_snapshot[0].f.unused[8] );
tran (\sa_snapshot[0][59] , \sa_snapshot[0].r.part1[27] );
tran (\sa_snapshot[0][59] , \sa_snapshot[0].f.unused[9] );
tran (\sa_snapshot[0][60] , \sa_snapshot[0].r.part1[28] );
tran (\sa_snapshot[0][60] , \sa_snapshot[0].f.unused[10] );
tran (\sa_snapshot[0][61] , \sa_snapshot[0].r.part1[29] );
tran (\sa_snapshot[0][61] , \sa_snapshot[0].f.unused[11] );
tran (\sa_snapshot[0][62] , \sa_snapshot[0].r.part1[30] );
tran (\sa_snapshot[0][62] , \sa_snapshot[0].f.unused[12] );
tran (\sa_snapshot[0][63] , \sa_snapshot[0].r.part1[31] );
tran (\sa_snapshot[0][63] , \sa_snapshot[0].f.unused[13] );
tran (\sa_snapshot[1][0] , \sa_snapshot[1].r.part0[0] );
tran (\sa_snapshot[1][0] , \sa_snapshot[1].f.lower[0] );
tran (\sa_snapshot[1][1] , \sa_snapshot[1].r.part0[1] );
tran (\sa_snapshot[1][1] , \sa_snapshot[1].f.lower[1] );
tran (\sa_snapshot[1][2] , \sa_snapshot[1].r.part0[2] );
tran (\sa_snapshot[1][2] , \sa_snapshot[1].f.lower[2] );
tran (\sa_snapshot[1][3] , \sa_snapshot[1].r.part0[3] );
tran (\sa_snapshot[1][3] , \sa_snapshot[1].f.lower[3] );
tran (\sa_snapshot[1][4] , \sa_snapshot[1].r.part0[4] );
tran (\sa_snapshot[1][4] , \sa_snapshot[1].f.lower[4] );
tran (\sa_snapshot[1][5] , \sa_snapshot[1].r.part0[5] );
tran (\sa_snapshot[1][5] , \sa_snapshot[1].f.lower[5] );
tran (\sa_snapshot[1][6] , \sa_snapshot[1].r.part0[6] );
tran (\sa_snapshot[1][6] , \sa_snapshot[1].f.lower[6] );
tran (\sa_snapshot[1][7] , \sa_snapshot[1].r.part0[7] );
tran (\sa_snapshot[1][7] , \sa_snapshot[1].f.lower[7] );
tran (\sa_snapshot[1][8] , \sa_snapshot[1].r.part0[8] );
tran (\sa_snapshot[1][8] , \sa_snapshot[1].f.lower[8] );
tran (\sa_snapshot[1][9] , \sa_snapshot[1].r.part0[9] );
tran (\sa_snapshot[1][9] , \sa_snapshot[1].f.lower[9] );
tran (\sa_snapshot[1][10] , \sa_snapshot[1].r.part0[10] );
tran (\sa_snapshot[1][10] , \sa_snapshot[1].f.lower[10] );
tran (\sa_snapshot[1][11] , \sa_snapshot[1].r.part0[11] );
tran (\sa_snapshot[1][11] , \sa_snapshot[1].f.lower[11] );
tran (\sa_snapshot[1][12] , \sa_snapshot[1].r.part0[12] );
tran (\sa_snapshot[1][12] , \sa_snapshot[1].f.lower[12] );
tran (\sa_snapshot[1][13] , \sa_snapshot[1].r.part0[13] );
tran (\sa_snapshot[1][13] , \sa_snapshot[1].f.lower[13] );
tran (\sa_snapshot[1][14] , \sa_snapshot[1].r.part0[14] );
tran (\sa_snapshot[1][14] , \sa_snapshot[1].f.lower[14] );
tran (\sa_snapshot[1][15] , \sa_snapshot[1].r.part0[15] );
tran (\sa_snapshot[1][15] , \sa_snapshot[1].f.lower[15] );
tran (\sa_snapshot[1][16] , \sa_snapshot[1].r.part0[16] );
tran (\sa_snapshot[1][16] , \sa_snapshot[1].f.lower[16] );
tran (\sa_snapshot[1][17] , \sa_snapshot[1].r.part0[17] );
tran (\sa_snapshot[1][17] , \sa_snapshot[1].f.lower[17] );
tran (\sa_snapshot[1][18] , \sa_snapshot[1].r.part0[18] );
tran (\sa_snapshot[1][18] , \sa_snapshot[1].f.lower[18] );
tran (\sa_snapshot[1][19] , \sa_snapshot[1].r.part0[19] );
tran (\sa_snapshot[1][19] , \sa_snapshot[1].f.lower[19] );
tran (\sa_snapshot[1][20] , \sa_snapshot[1].r.part0[20] );
tran (\sa_snapshot[1][20] , \sa_snapshot[1].f.lower[20] );
tran (\sa_snapshot[1][21] , \sa_snapshot[1].r.part0[21] );
tran (\sa_snapshot[1][21] , \sa_snapshot[1].f.lower[21] );
tran (\sa_snapshot[1][22] , \sa_snapshot[1].r.part0[22] );
tran (\sa_snapshot[1][22] , \sa_snapshot[1].f.lower[22] );
tran (\sa_snapshot[1][23] , \sa_snapshot[1].r.part0[23] );
tran (\sa_snapshot[1][23] , \sa_snapshot[1].f.lower[23] );
tran (\sa_snapshot[1][24] , \sa_snapshot[1].r.part0[24] );
tran (\sa_snapshot[1][24] , \sa_snapshot[1].f.lower[24] );
tran (\sa_snapshot[1][25] , \sa_snapshot[1].r.part0[25] );
tran (\sa_snapshot[1][25] , \sa_snapshot[1].f.lower[25] );
tran (\sa_snapshot[1][26] , \sa_snapshot[1].r.part0[26] );
tran (\sa_snapshot[1][26] , \sa_snapshot[1].f.lower[26] );
tran (\sa_snapshot[1][27] , \sa_snapshot[1].r.part0[27] );
tran (\sa_snapshot[1][27] , \sa_snapshot[1].f.lower[27] );
tran (\sa_snapshot[1][28] , \sa_snapshot[1].r.part0[28] );
tran (\sa_snapshot[1][28] , \sa_snapshot[1].f.lower[28] );
tran (\sa_snapshot[1][29] , \sa_snapshot[1].r.part0[29] );
tran (\sa_snapshot[1][29] , \sa_snapshot[1].f.lower[29] );
tran (\sa_snapshot[1][30] , \sa_snapshot[1].r.part0[30] );
tran (\sa_snapshot[1][30] , \sa_snapshot[1].f.lower[30] );
tran (\sa_snapshot[1][31] , \sa_snapshot[1].r.part0[31] );
tran (\sa_snapshot[1][31] , \sa_snapshot[1].f.lower[31] );
tran (\sa_snapshot[1][32] , \sa_snapshot[1].r.part1[0] );
tran (\sa_snapshot[1][32] , \sa_snapshot[1].f.upper[0] );
tran (\sa_snapshot[1][33] , \sa_snapshot[1].r.part1[1] );
tran (\sa_snapshot[1][33] , \sa_snapshot[1].f.upper[1] );
tran (\sa_snapshot[1][34] , \sa_snapshot[1].r.part1[2] );
tran (\sa_snapshot[1][34] , \sa_snapshot[1].f.upper[2] );
tran (\sa_snapshot[1][35] , \sa_snapshot[1].r.part1[3] );
tran (\sa_snapshot[1][35] , \sa_snapshot[1].f.upper[3] );
tran (\sa_snapshot[1][36] , \sa_snapshot[1].r.part1[4] );
tran (\sa_snapshot[1][36] , \sa_snapshot[1].f.upper[4] );
tran (\sa_snapshot[1][37] , \sa_snapshot[1].r.part1[5] );
tran (\sa_snapshot[1][37] , \sa_snapshot[1].f.upper[5] );
tran (\sa_snapshot[1][38] , \sa_snapshot[1].r.part1[6] );
tran (\sa_snapshot[1][38] , \sa_snapshot[1].f.upper[6] );
tran (\sa_snapshot[1][39] , \sa_snapshot[1].r.part1[7] );
tran (\sa_snapshot[1][39] , \sa_snapshot[1].f.upper[7] );
tran (\sa_snapshot[1][40] , \sa_snapshot[1].r.part1[8] );
tran (\sa_snapshot[1][40] , \sa_snapshot[1].f.upper[8] );
tran (\sa_snapshot[1][41] , \sa_snapshot[1].r.part1[9] );
tran (\sa_snapshot[1][41] , \sa_snapshot[1].f.upper[9] );
tran (\sa_snapshot[1][42] , \sa_snapshot[1].r.part1[10] );
tran (\sa_snapshot[1][42] , \sa_snapshot[1].f.upper[10] );
tran (\sa_snapshot[1][43] , \sa_snapshot[1].r.part1[11] );
tran (\sa_snapshot[1][43] , \sa_snapshot[1].f.upper[11] );
tran (\sa_snapshot[1][44] , \sa_snapshot[1].r.part1[12] );
tran (\sa_snapshot[1][44] , \sa_snapshot[1].f.upper[12] );
tran (\sa_snapshot[1][45] , \sa_snapshot[1].r.part1[13] );
tran (\sa_snapshot[1][45] , \sa_snapshot[1].f.upper[13] );
tran (\sa_snapshot[1][46] , \sa_snapshot[1].r.part1[14] );
tran (\sa_snapshot[1][46] , \sa_snapshot[1].f.upper[14] );
tran (\sa_snapshot[1][47] , \sa_snapshot[1].r.part1[15] );
tran (\sa_snapshot[1][47] , \sa_snapshot[1].f.upper[15] );
tran (\sa_snapshot[1][48] , \sa_snapshot[1].r.part1[16] );
tran (\sa_snapshot[1][48] , \sa_snapshot[1].f.upper[16] );
tran (\sa_snapshot[1][49] , \sa_snapshot[1].r.part1[17] );
tran (\sa_snapshot[1][49] , \sa_snapshot[1].f.upper[17] );
tran (\sa_snapshot[1][50] , \sa_snapshot[1].r.part1[18] );
tran (\sa_snapshot[1][50] , \sa_snapshot[1].f.unused[0] );
tran (\sa_snapshot[1][51] , \sa_snapshot[1].r.part1[19] );
tran (\sa_snapshot[1][51] , \sa_snapshot[1].f.unused[1] );
tran (\sa_snapshot[1][52] , \sa_snapshot[1].r.part1[20] );
tran (\sa_snapshot[1][52] , \sa_snapshot[1].f.unused[2] );
tran (\sa_snapshot[1][53] , \sa_snapshot[1].r.part1[21] );
tran (\sa_snapshot[1][53] , \sa_snapshot[1].f.unused[3] );
tran (\sa_snapshot[1][54] , \sa_snapshot[1].r.part1[22] );
tran (\sa_snapshot[1][54] , \sa_snapshot[1].f.unused[4] );
tran (\sa_snapshot[1][55] , \sa_snapshot[1].r.part1[23] );
tran (\sa_snapshot[1][55] , \sa_snapshot[1].f.unused[5] );
tran (\sa_snapshot[1][56] , \sa_snapshot[1].r.part1[24] );
tran (\sa_snapshot[1][56] , \sa_snapshot[1].f.unused[6] );
tran (\sa_snapshot[1][57] , \sa_snapshot[1].r.part1[25] );
tran (\sa_snapshot[1][57] , \sa_snapshot[1].f.unused[7] );
tran (\sa_snapshot[1][58] , \sa_snapshot[1].r.part1[26] );
tran (\sa_snapshot[1][58] , \sa_snapshot[1].f.unused[8] );
tran (\sa_snapshot[1][59] , \sa_snapshot[1].r.part1[27] );
tran (\sa_snapshot[1][59] , \sa_snapshot[1].f.unused[9] );
tran (\sa_snapshot[1][60] , \sa_snapshot[1].r.part1[28] );
tran (\sa_snapshot[1][60] , \sa_snapshot[1].f.unused[10] );
tran (\sa_snapshot[1][61] , \sa_snapshot[1].r.part1[29] );
tran (\sa_snapshot[1][61] , \sa_snapshot[1].f.unused[11] );
tran (\sa_snapshot[1][62] , \sa_snapshot[1].r.part1[30] );
tran (\sa_snapshot[1][62] , \sa_snapshot[1].f.unused[12] );
tran (\sa_snapshot[1][63] , \sa_snapshot[1].r.part1[31] );
tran (\sa_snapshot[1][63] , \sa_snapshot[1].f.unused[13] );
tran (\sa_snapshot[2][0] , \sa_snapshot[2].r.part0[0] );
tran (\sa_snapshot[2][0] , \sa_snapshot[2].f.lower[0] );
tran (\sa_snapshot[2][1] , \sa_snapshot[2].r.part0[1] );
tran (\sa_snapshot[2][1] , \sa_snapshot[2].f.lower[1] );
tran (\sa_snapshot[2][2] , \sa_snapshot[2].r.part0[2] );
tran (\sa_snapshot[2][2] , \sa_snapshot[2].f.lower[2] );
tran (\sa_snapshot[2][3] , \sa_snapshot[2].r.part0[3] );
tran (\sa_snapshot[2][3] , \sa_snapshot[2].f.lower[3] );
tran (\sa_snapshot[2][4] , \sa_snapshot[2].r.part0[4] );
tran (\sa_snapshot[2][4] , \sa_snapshot[2].f.lower[4] );
tran (\sa_snapshot[2][5] , \sa_snapshot[2].r.part0[5] );
tran (\sa_snapshot[2][5] , \sa_snapshot[2].f.lower[5] );
tran (\sa_snapshot[2][6] , \sa_snapshot[2].r.part0[6] );
tran (\sa_snapshot[2][6] , \sa_snapshot[2].f.lower[6] );
tran (\sa_snapshot[2][7] , \sa_snapshot[2].r.part0[7] );
tran (\sa_snapshot[2][7] , \sa_snapshot[2].f.lower[7] );
tran (\sa_snapshot[2][8] , \sa_snapshot[2].r.part0[8] );
tran (\sa_snapshot[2][8] , \sa_snapshot[2].f.lower[8] );
tran (\sa_snapshot[2][9] , \sa_snapshot[2].r.part0[9] );
tran (\sa_snapshot[2][9] , \sa_snapshot[2].f.lower[9] );
tran (\sa_snapshot[2][10] , \sa_snapshot[2].r.part0[10] );
tran (\sa_snapshot[2][10] , \sa_snapshot[2].f.lower[10] );
tran (\sa_snapshot[2][11] , \sa_snapshot[2].r.part0[11] );
tran (\sa_snapshot[2][11] , \sa_snapshot[2].f.lower[11] );
tran (\sa_snapshot[2][12] , \sa_snapshot[2].r.part0[12] );
tran (\sa_snapshot[2][12] , \sa_snapshot[2].f.lower[12] );
tran (\sa_snapshot[2][13] , \sa_snapshot[2].r.part0[13] );
tran (\sa_snapshot[2][13] , \sa_snapshot[2].f.lower[13] );
tran (\sa_snapshot[2][14] , \sa_snapshot[2].r.part0[14] );
tran (\sa_snapshot[2][14] , \sa_snapshot[2].f.lower[14] );
tran (\sa_snapshot[2][15] , \sa_snapshot[2].r.part0[15] );
tran (\sa_snapshot[2][15] , \sa_snapshot[2].f.lower[15] );
tran (\sa_snapshot[2][16] , \sa_snapshot[2].r.part0[16] );
tran (\sa_snapshot[2][16] , \sa_snapshot[2].f.lower[16] );
tran (\sa_snapshot[2][17] , \sa_snapshot[2].r.part0[17] );
tran (\sa_snapshot[2][17] , \sa_snapshot[2].f.lower[17] );
tran (\sa_snapshot[2][18] , \sa_snapshot[2].r.part0[18] );
tran (\sa_snapshot[2][18] , \sa_snapshot[2].f.lower[18] );
tran (\sa_snapshot[2][19] , \sa_snapshot[2].r.part0[19] );
tran (\sa_snapshot[2][19] , \sa_snapshot[2].f.lower[19] );
tran (\sa_snapshot[2][20] , \sa_snapshot[2].r.part0[20] );
tran (\sa_snapshot[2][20] , \sa_snapshot[2].f.lower[20] );
tran (\sa_snapshot[2][21] , \sa_snapshot[2].r.part0[21] );
tran (\sa_snapshot[2][21] , \sa_snapshot[2].f.lower[21] );
tran (\sa_snapshot[2][22] , \sa_snapshot[2].r.part0[22] );
tran (\sa_snapshot[2][22] , \sa_snapshot[2].f.lower[22] );
tran (\sa_snapshot[2][23] , \sa_snapshot[2].r.part0[23] );
tran (\sa_snapshot[2][23] , \sa_snapshot[2].f.lower[23] );
tran (\sa_snapshot[2][24] , \sa_snapshot[2].r.part0[24] );
tran (\sa_snapshot[2][24] , \sa_snapshot[2].f.lower[24] );
tran (\sa_snapshot[2][25] , \sa_snapshot[2].r.part0[25] );
tran (\sa_snapshot[2][25] , \sa_snapshot[2].f.lower[25] );
tran (\sa_snapshot[2][26] , \sa_snapshot[2].r.part0[26] );
tran (\sa_snapshot[2][26] , \sa_snapshot[2].f.lower[26] );
tran (\sa_snapshot[2][27] , \sa_snapshot[2].r.part0[27] );
tran (\sa_snapshot[2][27] , \sa_snapshot[2].f.lower[27] );
tran (\sa_snapshot[2][28] , \sa_snapshot[2].r.part0[28] );
tran (\sa_snapshot[2][28] , \sa_snapshot[2].f.lower[28] );
tran (\sa_snapshot[2][29] , \sa_snapshot[2].r.part0[29] );
tran (\sa_snapshot[2][29] , \sa_snapshot[2].f.lower[29] );
tran (\sa_snapshot[2][30] , \sa_snapshot[2].r.part0[30] );
tran (\sa_snapshot[2][30] , \sa_snapshot[2].f.lower[30] );
tran (\sa_snapshot[2][31] , \sa_snapshot[2].r.part0[31] );
tran (\sa_snapshot[2][31] , \sa_snapshot[2].f.lower[31] );
tran (\sa_snapshot[2][32] , \sa_snapshot[2].r.part1[0] );
tran (\sa_snapshot[2][32] , \sa_snapshot[2].f.upper[0] );
tran (\sa_snapshot[2][33] , \sa_snapshot[2].r.part1[1] );
tran (\sa_snapshot[2][33] , \sa_snapshot[2].f.upper[1] );
tran (\sa_snapshot[2][34] , \sa_snapshot[2].r.part1[2] );
tran (\sa_snapshot[2][34] , \sa_snapshot[2].f.upper[2] );
tran (\sa_snapshot[2][35] , \sa_snapshot[2].r.part1[3] );
tran (\sa_snapshot[2][35] , \sa_snapshot[2].f.upper[3] );
tran (\sa_snapshot[2][36] , \sa_snapshot[2].r.part1[4] );
tran (\sa_snapshot[2][36] , \sa_snapshot[2].f.upper[4] );
tran (\sa_snapshot[2][37] , \sa_snapshot[2].r.part1[5] );
tran (\sa_snapshot[2][37] , \sa_snapshot[2].f.upper[5] );
tran (\sa_snapshot[2][38] , \sa_snapshot[2].r.part1[6] );
tran (\sa_snapshot[2][38] , \sa_snapshot[2].f.upper[6] );
tran (\sa_snapshot[2][39] , \sa_snapshot[2].r.part1[7] );
tran (\sa_snapshot[2][39] , \sa_snapshot[2].f.upper[7] );
tran (\sa_snapshot[2][40] , \sa_snapshot[2].r.part1[8] );
tran (\sa_snapshot[2][40] , \sa_snapshot[2].f.upper[8] );
tran (\sa_snapshot[2][41] , \sa_snapshot[2].r.part1[9] );
tran (\sa_snapshot[2][41] , \sa_snapshot[2].f.upper[9] );
tran (\sa_snapshot[2][42] , \sa_snapshot[2].r.part1[10] );
tran (\sa_snapshot[2][42] , \sa_snapshot[2].f.upper[10] );
tran (\sa_snapshot[2][43] , \sa_snapshot[2].r.part1[11] );
tran (\sa_snapshot[2][43] , \sa_snapshot[2].f.upper[11] );
tran (\sa_snapshot[2][44] , \sa_snapshot[2].r.part1[12] );
tran (\sa_snapshot[2][44] , \sa_snapshot[2].f.upper[12] );
tran (\sa_snapshot[2][45] , \sa_snapshot[2].r.part1[13] );
tran (\sa_snapshot[2][45] , \sa_snapshot[2].f.upper[13] );
tran (\sa_snapshot[2][46] , \sa_snapshot[2].r.part1[14] );
tran (\sa_snapshot[2][46] , \sa_snapshot[2].f.upper[14] );
tran (\sa_snapshot[2][47] , \sa_snapshot[2].r.part1[15] );
tran (\sa_snapshot[2][47] , \sa_snapshot[2].f.upper[15] );
tran (\sa_snapshot[2][48] , \sa_snapshot[2].r.part1[16] );
tran (\sa_snapshot[2][48] , \sa_snapshot[2].f.upper[16] );
tran (\sa_snapshot[2][49] , \sa_snapshot[2].r.part1[17] );
tran (\sa_snapshot[2][49] , \sa_snapshot[2].f.upper[17] );
tran (\sa_snapshot[2][50] , \sa_snapshot[2].r.part1[18] );
tran (\sa_snapshot[2][50] , \sa_snapshot[2].f.unused[0] );
tran (\sa_snapshot[2][51] , \sa_snapshot[2].r.part1[19] );
tran (\sa_snapshot[2][51] , \sa_snapshot[2].f.unused[1] );
tran (\sa_snapshot[2][52] , \sa_snapshot[2].r.part1[20] );
tran (\sa_snapshot[2][52] , \sa_snapshot[2].f.unused[2] );
tran (\sa_snapshot[2][53] , \sa_snapshot[2].r.part1[21] );
tran (\sa_snapshot[2][53] , \sa_snapshot[2].f.unused[3] );
tran (\sa_snapshot[2][54] , \sa_snapshot[2].r.part1[22] );
tran (\sa_snapshot[2][54] , \sa_snapshot[2].f.unused[4] );
tran (\sa_snapshot[2][55] , \sa_snapshot[2].r.part1[23] );
tran (\sa_snapshot[2][55] , \sa_snapshot[2].f.unused[5] );
tran (\sa_snapshot[2][56] , \sa_snapshot[2].r.part1[24] );
tran (\sa_snapshot[2][56] , \sa_snapshot[2].f.unused[6] );
tran (\sa_snapshot[2][57] , \sa_snapshot[2].r.part1[25] );
tran (\sa_snapshot[2][57] , \sa_snapshot[2].f.unused[7] );
tran (\sa_snapshot[2][58] , \sa_snapshot[2].r.part1[26] );
tran (\sa_snapshot[2][58] , \sa_snapshot[2].f.unused[8] );
tran (\sa_snapshot[2][59] , \sa_snapshot[2].r.part1[27] );
tran (\sa_snapshot[2][59] , \sa_snapshot[2].f.unused[9] );
tran (\sa_snapshot[2][60] , \sa_snapshot[2].r.part1[28] );
tran (\sa_snapshot[2][60] , \sa_snapshot[2].f.unused[10] );
tran (\sa_snapshot[2][61] , \sa_snapshot[2].r.part1[29] );
tran (\sa_snapshot[2][61] , \sa_snapshot[2].f.unused[11] );
tran (\sa_snapshot[2][62] , \sa_snapshot[2].r.part1[30] );
tran (\sa_snapshot[2][62] , \sa_snapshot[2].f.unused[12] );
tran (\sa_snapshot[2][63] , \sa_snapshot[2].r.part1[31] );
tran (\sa_snapshot[2][63] , \sa_snapshot[2].f.unused[13] );
tran (\sa_snapshot[3][0] , \sa_snapshot[3].r.part0[0] );
tran (\sa_snapshot[3][0] , \sa_snapshot[3].f.lower[0] );
tran (\sa_snapshot[3][1] , \sa_snapshot[3].r.part0[1] );
tran (\sa_snapshot[3][1] , \sa_snapshot[3].f.lower[1] );
tran (\sa_snapshot[3][2] , \sa_snapshot[3].r.part0[2] );
tran (\sa_snapshot[3][2] , \sa_snapshot[3].f.lower[2] );
tran (\sa_snapshot[3][3] , \sa_snapshot[3].r.part0[3] );
tran (\sa_snapshot[3][3] , \sa_snapshot[3].f.lower[3] );
tran (\sa_snapshot[3][4] , \sa_snapshot[3].r.part0[4] );
tran (\sa_snapshot[3][4] , \sa_snapshot[3].f.lower[4] );
tran (\sa_snapshot[3][5] , \sa_snapshot[3].r.part0[5] );
tran (\sa_snapshot[3][5] , \sa_snapshot[3].f.lower[5] );
tran (\sa_snapshot[3][6] , \sa_snapshot[3].r.part0[6] );
tran (\sa_snapshot[3][6] , \sa_snapshot[3].f.lower[6] );
tran (\sa_snapshot[3][7] , \sa_snapshot[3].r.part0[7] );
tran (\sa_snapshot[3][7] , \sa_snapshot[3].f.lower[7] );
tran (\sa_snapshot[3][8] , \sa_snapshot[3].r.part0[8] );
tran (\sa_snapshot[3][8] , \sa_snapshot[3].f.lower[8] );
tran (\sa_snapshot[3][9] , \sa_snapshot[3].r.part0[9] );
tran (\sa_snapshot[3][9] , \sa_snapshot[3].f.lower[9] );
tran (\sa_snapshot[3][10] , \sa_snapshot[3].r.part0[10] );
tran (\sa_snapshot[3][10] , \sa_snapshot[3].f.lower[10] );
tran (\sa_snapshot[3][11] , \sa_snapshot[3].r.part0[11] );
tran (\sa_snapshot[3][11] , \sa_snapshot[3].f.lower[11] );
tran (\sa_snapshot[3][12] , \sa_snapshot[3].r.part0[12] );
tran (\sa_snapshot[3][12] , \sa_snapshot[3].f.lower[12] );
tran (\sa_snapshot[3][13] , \sa_snapshot[3].r.part0[13] );
tran (\sa_snapshot[3][13] , \sa_snapshot[3].f.lower[13] );
tran (\sa_snapshot[3][14] , \sa_snapshot[3].r.part0[14] );
tran (\sa_snapshot[3][14] , \sa_snapshot[3].f.lower[14] );
tran (\sa_snapshot[3][15] , \sa_snapshot[3].r.part0[15] );
tran (\sa_snapshot[3][15] , \sa_snapshot[3].f.lower[15] );
tran (\sa_snapshot[3][16] , \sa_snapshot[3].r.part0[16] );
tran (\sa_snapshot[3][16] , \sa_snapshot[3].f.lower[16] );
tran (\sa_snapshot[3][17] , \sa_snapshot[3].r.part0[17] );
tran (\sa_snapshot[3][17] , \sa_snapshot[3].f.lower[17] );
tran (\sa_snapshot[3][18] , \sa_snapshot[3].r.part0[18] );
tran (\sa_snapshot[3][18] , \sa_snapshot[3].f.lower[18] );
tran (\sa_snapshot[3][19] , \sa_snapshot[3].r.part0[19] );
tran (\sa_snapshot[3][19] , \sa_snapshot[3].f.lower[19] );
tran (\sa_snapshot[3][20] , \sa_snapshot[3].r.part0[20] );
tran (\sa_snapshot[3][20] , \sa_snapshot[3].f.lower[20] );
tran (\sa_snapshot[3][21] , \sa_snapshot[3].r.part0[21] );
tran (\sa_snapshot[3][21] , \sa_snapshot[3].f.lower[21] );
tran (\sa_snapshot[3][22] , \sa_snapshot[3].r.part0[22] );
tran (\sa_snapshot[3][22] , \sa_snapshot[3].f.lower[22] );
tran (\sa_snapshot[3][23] , \sa_snapshot[3].r.part0[23] );
tran (\sa_snapshot[3][23] , \sa_snapshot[3].f.lower[23] );
tran (\sa_snapshot[3][24] , \sa_snapshot[3].r.part0[24] );
tran (\sa_snapshot[3][24] , \sa_snapshot[3].f.lower[24] );
tran (\sa_snapshot[3][25] , \sa_snapshot[3].r.part0[25] );
tran (\sa_snapshot[3][25] , \sa_snapshot[3].f.lower[25] );
tran (\sa_snapshot[3][26] , \sa_snapshot[3].r.part0[26] );
tran (\sa_snapshot[3][26] , \sa_snapshot[3].f.lower[26] );
tran (\sa_snapshot[3][27] , \sa_snapshot[3].r.part0[27] );
tran (\sa_snapshot[3][27] , \sa_snapshot[3].f.lower[27] );
tran (\sa_snapshot[3][28] , \sa_snapshot[3].r.part0[28] );
tran (\sa_snapshot[3][28] , \sa_snapshot[3].f.lower[28] );
tran (\sa_snapshot[3][29] , \sa_snapshot[3].r.part0[29] );
tran (\sa_snapshot[3][29] , \sa_snapshot[3].f.lower[29] );
tran (\sa_snapshot[3][30] , \sa_snapshot[3].r.part0[30] );
tran (\sa_snapshot[3][30] , \sa_snapshot[3].f.lower[30] );
tran (\sa_snapshot[3][31] , \sa_snapshot[3].r.part0[31] );
tran (\sa_snapshot[3][31] , \sa_snapshot[3].f.lower[31] );
tran (\sa_snapshot[3][32] , \sa_snapshot[3].r.part1[0] );
tran (\sa_snapshot[3][32] , \sa_snapshot[3].f.upper[0] );
tran (\sa_snapshot[3][33] , \sa_snapshot[3].r.part1[1] );
tran (\sa_snapshot[3][33] , \sa_snapshot[3].f.upper[1] );
tran (\sa_snapshot[3][34] , \sa_snapshot[3].r.part1[2] );
tran (\sa_snapshot[3][34] , \sa_snapshot[3].f.upper[2] );
tran (\sa_snapshot[3][35] , \sa_snapshot[3].r.part1[3] );
tran (\sa_snapshot[3][35] , \sa_snapshot[3].f.upper[3] );
tran (\sa_snapshot[3][36] , \sa_snapshot[3].r.part1[4] );
tran (\sa_snapshot[3][36] , \sa_snapshot[3].f.upper[4] );
tran (\sa_snapshot[3][37] , \sa_snapshot[3].r.part1[5] );
tran (\sa_snapshot[3][37] , \sa_snapshot[3].f.upper[5] );
tran (\sa_snapshot[3][38] , \sa_snapshot[3].r.part1[6] );
tran (\sa_snapshot[3][38] , \sa_snapshot[3].f.upper[6] );
tran (\sa_snapshot[3][39] , \sa_snapshot[3].r.part1[7] );
tran (\sa_snapshot[3][39] , \sa_snapshot[3].f.upper[7] );
tran (\sa_snapshot[3][40] , \sa_snapshot[3].r.part1[8] );
tran (\sa_snapshot[3][40] , \sa_snapshot[3].f.upper[8] );
tran (\sa_snapshot[3][41] , \sa_snapshot[3].r.part1[9] );
tran (\sa_snapshot[3][41] , \sa_snapshot[3].f.upper[9] );
tran (\sa_snapshot[3][42] , \sa_snapshot[3].r.part1[10] );
tran (\sa_snapshot[3][42] , \sa_snapshot[3].f.upper[10] );
tran (\sa_snapshot[3][43] , \sa_snapshot[3].r.part1[11] );
tran (\sa_snapshot[3][43] , \sa_snapshot[3].f.upper[11] );
tran (\sa_snapshot[3][44] , \sa_snapshot[3].r.part1[12] );
tran (\sa_snapshot[3][44] , \sa_snapshot[3].f.upper[12] );
tran (\sa_snapshot[3][45] , \sa_snapshot[3].r.part1[13] );
tran (\sa_snapshot[3][45] , \sa_snapshot[3].f.upper[13] );
tran (\sa_snapshot[3][46] , \sa_snapshot[3].r.part1[14] );
tran (\sa_snapshot[3][46] , \sa_snapshot[3].f.upper[14] );
tran (\sa_snapshot[3][47] , \sa_snapshot[3].r.part1[15] );
tran (\sa_snapshot[3][47] , \sa_snapshot[3].f.upper[15] );
tran (\sa_snapshot[3][48] , \sa_snapshot[3].r.part1[16] );
tran (\sa_snapshot[3][48] , \sa_snapshot[3].f.upper[16] );
tran (\sa_snapshot[3][49] , \sa_snapshot[3].r.part1[17] );
tran (\sa_snapshot[3][49] , \sa_snapshot[3].f.upper[17] );
tran (\sa_snapshot[3][50] , \sa_snapshot[3].r.part1[18] );
tran (\sa_snapshot[3][50] , \sa_snapshot[3].f.unused[0] );
tran (\sa_snapshot[3][51] , \sa_snapshot[3].r.part1[19] );
tran (\sa_snapshot[3][51] , \sa_snapshot[3].f.unused[1] );
tran (\sa_snapshot[3][52] , \sa_snapshot[3].r.part1[20] );
tran (\sa_snapshot[3][52] , \sa_snapshot[3].f.unused[2] );
tran (\sa_snapshot[3][53] , \sa_snapshot[3].r.part1[21] );
tran (\sa_snapshot[3][53] , \sa_snapshot[3].f.unused[3] );
tran (\sa_snapshot[3][54] , \sa_snapshot[3].r.part1[22] );
tran (\sa_snapshot[3][54] , \sa_snapshot[3].f.unused[4] );
tran (\sa_snapshot[3][55] , \sa_snapshot[3].r.part1[23] );
tran (\sa_snapshot[3][55] , \sa_snapshot[3].f.unused[5] );
tran (\sa_snapshot[3][56] , \sa_snapshot[3].r.part1[24] );
tran (\sa_snapshot[3][56] , \sa_snapshot[3].f.unused[6] );
tran (\sa_snapshot[3][57] , \sa_snapshot[3].r.part1[25] );
tran (\sa_snapshot[3][57] , \sa_snapshot[3].f.unused[7] );
tran (\sa_snapshot[3][58] , \sa_snapshot[3].r.part1[26] );
tran (\sa_snapshot[3][58] , \sa_snapshot[3].f.unused[8] );
tran (\sa_snapshot[3][59] , \sa_snapshot[3].r.part1[27] );
tran (\sa_snapshot[3][59] , \sa_snapshot[3].f.unused[9] );
tran (\sa_snapshot[3][60] , \sa_snapshot[3].r.part1[28] );
tran (\sa_snapshot[3][60] , \sa_snapshot[3].f.unused[10] );
tran (\sa_snapshot[3][61] , \sa_snapshot[3].r.part1[29] );
tran (\sa_snapshot[3][61] , \sa_snapshot[3].f.unused[11] );
tran (\sa_snapshot[3][62] , \sa_snapshot[3].r.part1[30] );
tran (\sa_snapshot[3][62] , \sa_snapshot[3].f.unused[12] );
tran (\sa_snapshot[3][63] , \sa_snapshot[3].r.part1[31] );
tran (\sa_snapshot[3][63] , \sa_snapshot[3].f.unused[13] );
tran (\sa_snapshot[4][0] , \sa_snapshot[4].r.part0[0] );
tran (\sa_snapshot[4][0] , \sa_snapshot[4].f.lower[0] );
tran (\sa_snapshot[4][1] , \sa_snapshot[4].r.part0[1] );
tran (\sa_snapshot[4][1] , \sa_snapshot[4].f.lower[1] );
tran (\sa_snapshot[4][2] , \sa_snapshot[4].r.part0[2] );
tran (\sa_snapshot[4][2] , \sa_snapshot[4].f.lower[2] );
tran (\sa_snapshot[4][3] , \sa_snapshot[4].r.part0[3] );
tran (\sa_snapshot[4][3] , \sa_snapshot[4].f.lower[3] );
tran (\sa_snapshot[4][4] , \sa_snapshot[4].r.part0[4] );
tran (\sa_snapshot[4][4] , \sa_snapshot[4].f.lower[4] );
tran (\sa_snapshot[4][5] , \sa_snapshot[4].r.part0[5] );
tran (\sa_snapshot[4][5] , \sa_snapshot[4].f.lower[5] );
tran (\sa_snapshot[4][6] , \sa_snapshot[4].r.part0[6] );
tran (\sa_snapshot[4][6] , \sa_snapshot[4].f.lower[6] );
tran (\sa_snapshot[4][7] , \sa_snapshot[4].r.part0[7] );
tran (\sa_snapshot[4][7] , \sa_snapshot[4].f.lower[7] );
tran (\sa_snapshot[4][8] , \sa_snapshot[4].r.part0[8] );
tran (\sa_snapshot[4][8] , \sa_snapshot[4].f.lower[8] );
tran (\sa_snapshot[4][9] , \sa_snapshot[4].r.part0[9] );
tran (\sa_snapshot[4][9] , \sa_snapshot[4].f.lower[9] );
tran (\sa_snapshot[4][10] , \sa_snapshot[4].r.part0[10] );
tran (\sa_snapshot[4][10] , \sa_snapshot[4].f.lower[10] );
tran (\sa_snapshot[4][11] , \sa_snapshot[4].r.part0[11] );
tran (\sa_snapshot[4][11] , \sa_snapshot[4].f.lower[11] );
tran (\sa_snapshot[4][12] , \sa_snapshot[4].r.part0[12] );
tran (\sa_snapshot[4][12] , \sa_snapshot[4].f.lower[12] );
tran (\sa_snapshot[4][13] , \sa_snapshot[4].r.part0[13] );
tran (\sa_snapshot[4][13] , \sa_snapshot[4].f.lower[13] );
tran (\sa_snapshot[4][14] , \sa_snapshot[4].r.part0[14] );
tran (\sa_snapshot[4][14] , \sa_snapshot[4].f.lower[14] );
tran (\sa_snapshot[4][15] , \sa_snapshot[4].r.part0[15] );
tran (\sa_snapshot[4][15] , \sa_snapshot[4].f.lower[15] );
tran (\sa_snapshot[4][16] , \sa_snapshot[4].r.part0[16] );
tran (\sa_snapshot[4][16] , \sa_snapshot[4].f.lower[16] );
tran (\sa_snapshot[4][17] , \sa_snapshot[4].r.part0[17] );
tran (\sa_snapshot[4][17] , \sa_snapshot[4].f.lower[17] );
tran (\sa_snapshot[4][18] , \sa_snapshot[4].r.part0[18] );
tran (\sa_snapshot[4][18] , \sa_snapshot[4].f.lower[18] );
tran (\sa_snapshot[4][19] , \sa_snapshot[4].r.part0[19] );
tran (\sa_snapshot[4][19] , \sa_snapshot[4].f.lower[19] );
tran (\sa_snapshot[4][20] , \sa_snapshot[4].r.part0[20] );
tran (\sa_snapshot[4][20] , \sa_snapshot[4].f.lower[20] );
tran (\sa_snapshot[4][21] , \sa_snapshot[4].r.part0[21] );
tran (\sa_snapshot[4][21] , \sa_snapshot[4].f.lower[21] );
tran (\sa_snapshot[4][22] , \sa_snapshot[4].r.part0[22] );
tran (\sa_snapshot[4][22] , \sa_snapshot[4].f.lower[22] );
tran (\sa_snapshot[4][23] , \sa_snapshot[4].r.part0[23] );
tran (\sa_snapshot[4][23] , \sa_snapshot[4].f.lower[23] );
tran (\sa_snapshot[4][24] , \sa_snapshot[4].r.part0[24] );
tran (\sa_snapshot[4][24] , \sa_snapshot[4].f.lower[24] );
tran (\sa_snapshot[4][25] , \sa_snapshot[4].r.part0[25] );
tran (\sa_snapshot[4][25] , \sa_snapshot[4].f.lower[25] );
tran (\sa_snapshot[4][26] , \sa_snapshot[4].r.part0[26] );
tran (\sa_snapshot[4][26] , \sa_snapshot[4].f.lower[26] );
tran (\sa_snapshot[4][27] , \sa_snapshot[4].r.part0[27] );
tran (\sa_snapshot[4][27] , \sa_snapshot[4].f.lower[27] );
tran (\sa_snapshot[4][28] , \sa_snapshot[4].r.part0[28] );
tran (\sa_snapshot[4][28] , \sa_snapshot[4].f.lower[28] );
tran (\sa_snapshot[4][29] , \sa_snapshot[4].r.part0[29] );
tran (\sa_snapshot[4][29] , \sa_snapshot[4].f.lower[29] );
tran (\sa_snapshot[4][30] , \sa_snapshot[4].r.part0[30] );
tran (\sa_snapshot[4][30] , \sa_snapshot[4].f.lower[30] );
tran (\sa_snapshot[4][31] , \sa_snapshot[4].r.part0[31] );
tran (\sa_snapshot[4][31] , \sa_snapshot[4].f.lower[31] );
tran (\sa_snapshot[4][32] , \sa_snapshot[4].r.part1[0] );
tran (\sa_snapshot[4][32] , \sa_snapshot[4].f.upper[0] );
tran (\sa_snapshot[4][33] , \sa_snapshot[4].r.part1[1] );
tran (\sa_snapshot[4][33] , \sa_snapshot[4].f.upper[1] );
tran (\sa_snapshot[4][34] , \sa_snapshot[4].r.part1[2] );
tran (\sa_snapshot[4][34] , \sa_snapshot[4].f.upper[2] );
tran (\sa_snapshot[4][35] , \sa_snapshot[4].r.part1[3] );
tran (\sa_snapshot[4][35] , \sa_snapshot[4].f.upper[3] );
tran (\sa_snapshot[4][36] , \sa_snapshot[4].r.part1[4] );
tran (\sa_snapshot[4][36] , \sa_snapshot[4].f.upper[4] );
tran (\sa_snapshot[4][37] , \sa_snapshot[4].r.part1[5] );
tran (\sa_snapshot[4][37] , \sa_snapshot[4].f.upper[5] );
tran (\sa_snapshot[4][38] , \sa_snapshot[4].r.part1[6] );
tran (\sa_snapshot[4][38] , \sa_snapshot[4].f.upper[6] );
tran (\sa_snapshot[4][39] , \sa_snapshot[4].r.part1[7] );
tran (\sa_snapshot[4][39] , \sa_snapshot[4].f.upper[7] );
tran (\sa_snapshot[4][40] , \sa_snapshot[4].r.part1[8] );
tran (\sa_snapshot[4][40] , \sa_snapshot[4].f.upper[8] );
tran (\sa_snapshot[4][41] , \sa_snapshot[4].r.part1[9] );
tran (\sa_snapshot[4][41] , \sa_snapshot[4].f.upper[9] );
tran (\sa_snapshot[4][42] , \sa_snapshot[4].r.part1[10] );
tran (\sa_snapshot[4][42] , \sa_snapshot[4].f.upper[10] );
tran (\sa_snapshot[4][43] , \sa_snapshot[4].r.part1[11] );
tran (\sa_snapshot[4][43] , \sa_snapshot[4].f.upper[11] );
tran (\sa_snapshot[4][44] , \sa_snapshot[4].r.part1[12] );
tran (\sa_snapshot[4][44] , \sa_snapshot[4].f.upper[12] );
tran (\sa_snapshot[4][45] , \sa_snapshot[4].r.part1[13] );
tran (\sa_snapshot[4][45] , \sa_snapshot[4].f.upper[13] );
tran (\sa_snapshot[4][46] , \sa_snapshot[4].r.part1[14] );
tran (\sa_snapshot[4][46] , \sa_snapshot[4].f.upper[14] );
tran (\sa_snapshot[4][47] , \sa_snapshot[4].r.part1[15] );
tran (\sa_snapshot[4][47] , \sa_snapshot[4].f.upper[15] );
tran (\sa_snapshot[4][48] , \sa_snapshot[4].r.part1[16] );
tran (\sa_snapshot[4][48] , \sa_snapshot[4].f.upper[16] );
tran (\sa_snapshot[4][49] , \sa_snapshot[4].r.part1[17] );
tran (\sa_snapshot[4][49] , \sa_snapshot[4].f.upper[17] );
tran (\sa_snapshot[4][50] , \sa_snapshot[4].r.part1[18] );
tran (\sa_snapshot[4][50] , \sa_snapshot[4].f.unused[0] );
tran (\sa_snapshot[4][51] , \sa_snapshot[4].r.part1[19] );
tran (\sa_snapshot[4][51] , \sa_snapshot[4].f.unused[1] );
tran (\sa_snapshot[4][52] , \sa_snapshot[4].r.part1[20] );
tran (\sa_snapshot[4][52] , \sa_snapshot[4].f.unused[2] );
tran (\sa_snapshot[4][53] , \sa_snapshot[4].r.part1[21] );
tran (\sa_snapshot[4][53] , \sa_snapshot[4].f.unused[3] );
tran (\sa_snapshot[4][54] , \sa_snapshot[4].r.part1[22] );
tran (\sa_snapshot[4][54] , \sa_snapshot[4].f.unused[4] );
tran (\sa_snapshot[4][55] , \sa_snapshot[4].r.part1[23] );
tran (\sa_snapshot[4][55] , \sa_snapshot[4].f.unused[5] );
tran (\sa_snapshot[4][56] , \sa_snapshot[4].r.part1[24] );
tran (\sa_snapshot[4][56] , \sa_snapshot[4].f.unused[6] );
tran (\sa_snapshot[4][57] , \sa_snapshot[4].r.part1[25] );
tran (\sa_snapshot[4][57] , \sa_snapshot[4].f.unused[7] );
tran (\sa_snapshot[4][58] , \sa_snapshot[4].r.part1[26] );
tran (\sa_snapshot[4][58] , \sa_snapshot[4].f.unused[8] );
tran (\sa_snapshot[4][59] , \sa_snapshot[4].r.part1[27] );
tran (\sa_snapshot[4][59] , \sa_snapshot[4].f.unused[9] );
tran (\sa_snapshot[4][60] , \sa_snapshot[4].r.part1[28] );
tran (\sa_snapshot[4][60] , \sa_snapshot[4].f.unused[10] );
tran (\sa_snapshot[4][61] , \sa_snapshot[4].r.part1[29] );
tran (\sa_snapshot[4][61] , \sa_snapshot[4].f.unused[11] );
tran (\sa_snapshot[4][62] , \sa_snapshot[4].r.part1[30] );
tran (\sa_snapshot[4][62] , \sa_snapshot[4].f.unused[12] );
tran (\sa_snapshot[4][63] , \sa_snapshot[4].r.part1[31] );
tran (\sa_snapshot[4][63] , \sa_snapshot[4].f.unused[13] );
tran (\sa_snapshot[5][0] , \sa_snapshot[5].r.part0[0] );
tran (\sa_snapshot[5][0] , \sa_snapshot[5].f.lower[0] );
tran (\sa_snapshot[5][1] , \sa_snapshot[5].r.part0[1] );
tran (\sa_snapshot[5][1] , \sa_snapshot[5].f.lower[1] );
tran (\sa_snapshot[5][2] , \sa_snapshot[5].r.part0[2] );
tran (\sa_snapshot[5][2] , \sa_snapshot[5].f.lower[2] );
tran (\sa_snapshot[5][3] , \sa_snapshot[5].r.part0[3] );
tran (\sa_snapshot[5][3] , \sa_snapshot[5].f.lower[3] );
tran (\sa_snapshot[5][4] , \sa_snapshot[5].r.part0[4] );
tran (\sa_snapshot[5][4] , \sa_snapshot[5].f.lower[4] );
tran (\sa_snapshot[5][5] , \sa_snapshot[5].r.part0[5] );
tran (\sa_snapshot[5][5] , \sa_snapshot[5].f.lower[5] );
tran (\sa_snapshot[5][6] , \sa_snapshot[5].r.part0[6] );
tran (\sa_snapshot[5][6] , \sa_snapshot[5].f.lower[6] );
tran (\sa_snapshot[5][7] , \sa_snapshot[5].r.part0[7] );
tran (\sa_snapshot[5][7] , \sa_snapshot[5].f.lower[7] );
tran (\sa_snapshot[5][8] , \sa_snapshot[5].r.part0[8] );
tran (\sa_snapshot[5][8] , \sa_snapshot[5].f.lower[8] );
tran (\sa_snapshot[5][9] , \sa_snapshot[5].r.part0[9] );
tran (\sa_snapshot[5][9] , \sa_snapshot[5].f.lower[9] );
tran (\sa_snapshot[5][10] , \sa_snapshot[5].r.part0[10] );
tran (\sa_snapshot[5][10] , \sa_snapshot[5].f.lower[10] );
tran (\sa_snapshot[5][11] , \sa_snapshot[5].r.part0[11] );
tran (\sa_snapshot[5][11] , \sa_snapshot[5].f.lower[11] );
tran (\sa_snapshot[5][12] , \sa_snapshot[5].r.part0[12] );
tran (\sa_snapshot[5][12] , \sa_snapshot[5].f.lower[12] );
tran (\sa_snapshot[5][13] , \sa_snapshot[5].r.part0[13] );
tran (\sa_snapshot[5][13] , \sa_snapshot[5].f.lower[13] );
tran (\sa_snapshot[5][14] , \sa_snapshot[5].r.part0[14] );
tran (\sa_snapshot[5][14] , \sa_snapshot[5].f.lower[14] );
tran (\sa_snapshot[5][15] , \sa_snapshot[5].r.part0[15] );
tran (\sa_snapshot[5][15] , \sa_snapshot[5].f.lower[15] );
tran (\sa_snapshot[5][16] , \sa_snapshot[5].r.part0[16] );
tran (\sa_snapshot[5][16] , \sa_snapshot[5].f.lower[16] );
tran (\sa_snapshot[5][17] , \sa_snapshot[5].r.part0[17] );
tran (\sa_snapshot[5][17] , \sa_snapshot[5].f.lower[17] );
tran (\sa_snapshot[5][18] , \sa_snapshot[5].r.part0[18] );
tran (\sa_snapshot[5][18] , \sa_snapshot[5].f.lower[18] );
tran (\sa_snapshot[5][19] , \sa_snapshot[5].r.part0[19] );
tran (\sa_snapshot[5][19] , \sa_snapshot[5].f.lower[19] );
tran (\sa_snapshot[5][20] , \sa_snapshot[5].r.part0[20] );
tran (\sa_snapshot[5][20] , \sa_snapshot[5].f.lower[20] );
tran (\sa_snapshot[5][21] , \sa_snapshot[5].r.part0[21] );
tran (\sa_snapshot[5][21] , \sa_snapshot[5].f.lower[21] );
tran (\sa_snapshot[5][22] , \sa_snapshot[5].r.part0[22] );
tran (\sa_snapshot[5][22] , \sa_snapshot[5].f.lower[22] );
tran (\sa_snapshot[5][23] , \sa_snapshot[5].r.part0[23] );
tran (\sa_snapshot[5][23] , \sa_snapshot[5].f.lower[23] );
tran (\sa_snapshot[5][24] , \sa_snapshot[5].r.part0[24] );
tran (\sa_snapshot[5][24] , \sa_snapshot[5].f.lower[24] );
tran (\sa_snapshot[5][25] , \sa_snapshot[5].r.part0[25] );
tran (\sa_snapshot[5][25] , \sa_snapshot[5].f.lower[25] );
tran (\sa_snapshot[5][26] , \sa_snapshot[5].r.part0[26] );
tran (\sa_snapshot[5][26] , \sa_snapshot[5].f.lower[26] );
tran (\sa_snapshot[5][27] , \sa_snapshot[5].r.part0[27] );
tran (\sa_snapshot[5][27] , \sa_snapshot[5].f.lower[27] );
tran (\sa_snapshot[5][28] , \sa_snapshot[5].r.part0[28] );
tran (\sa_snapshot[5][28] , \sa_snapshot[5].f.lower[28] );
tran (\sa_snapshot[5][29] , \sa_snapshot[5].r.part0[29] );
tran (\sa_snapshot[5][29] , \sa_snapshot[5].f.lower[29] );
tran (\sa_snapshot[5][30] , \sa_snapshot[5].r.part0[30] );
tran (\sa_snapshot[5][30] , \sa_snapshot[5].f.lower[30] );
tran (\sa_snapshot[5][31] , \sa_snapshot[5].r.part0[31] );
tran (\sa_snapshot[5][31] , \sa_snapshot[5].f.lower[31] );
tran (\sa_snapshot[5][32] , \sa_snapshot[5].r.part1[0] );
tran (\sa_snapshot[5][32] , \sa_snapshot[5].f.upper[0] );
tran (\sa_snapshot[5][33] , \sa_snapshot[5].r.part1[1] );
tran (\sa_snapshot[5][33] , \sa_snapshot[5].f.upper[1] );
tran (\sa_snapshot[5][34] , \sa_snapshot[5].r.part1[2] );
tran (\sa_snapshot[5][34] , \sa_snapshot[5].f.upper[2] );
tran (\sa_snapshot[5][35] , \sa_snapshot[5].r.part1[3] );
tran (\sa_snapshot[5][35] , \sa_snapshot[5].f.upper[3] );
tran (\sa_snapshot[5][36] , \sa_snapshot[5].r.part1[4] );
tran (\sa_snapshot[5][36] , \sa_snapshot[5].f.upper[4] );
tran (\sa_snapshot[5][37] , \sa_snapshot[5].r.part1[5] );
tran (\sa_snapshot[5][37] , \sa_snapshot[5].f.upper[5] );
tran (\sa_snapshot[5][38] , \sa_snapshot[5].r.part1[6] );
tran (\sa_snapshot[5][38] , \sa_snapshot[5].f.upper[6] );
tran (\sa_snapshot[5][39] , \sa_snapshot[5].r.part1[7] );
tran (\sa_snapshot[5][39] , \sa_snapshot[5].f.upper[7] );
tran (\sa_snapshot[5][40] , \sa_snapshot[5].r.part1[8] );
tran (\sa_snapshot[5][40] , \sa_snapshot[5].f.upper[8] );
tran (\sa_snapshot[5][41] , \sa_snapshot[5].r.part1[9] );
tran (\sa_snapshot[5][41] , \sa_snapshot[5].f.upper[9] );
tran (\sa_snapshot[5][42] , \sa_snapshot[5].r.part1[10] );
tran (\sa_snapshot[5][42] , \sa_snapshot[5].f.upper[10] );
tran (\sa_snapshot[5][43] , \sa_snapshot[5].r.part1[11] );
tran (\sa_snapshot[5][43] , \sa_snapshot[5].f.upper[11] );
tran (\sa_snapshot[5][44] , \sa_snapshot[5].r.part1[12] );
tran (\sa_snapshot[5][44] , \sa_snapshot[5].f.upper[12] );
tran (\sa_snapshot[5][45] , \sa_snapshot[5].r.part1[13] );
tran (\sa_snapshot[5][45] , \sa_snapshot[5].f.upper[13] );
tran (\sa_snapshot[5][46] , \sa_snapshot[5].r.part1[14] );
tran (\sa_snapshot[5][46] , \sa_snapshot[5].f.upper[14] );
tran (\sa_snapshot[5][47] , \sa_snapshot[5].r.part1[15] );
tran (\sa_snapshot[5][47] , \sa_snapshot[5].f.upper[15] );
tran (\sa_snapshot[5][48] , \sa_snapshot[5].r.part1[16] );
tran (\sa_snapshot[5][48] , \sa_snapshot[5].f.upper[16] );
tran (\sa_snapshot[5][49] , \sa_snapshot[5].r.part1[17] );
tran (\sa_snapshot[5][49] , \sa_snapshot[5].f.upper[17] );
tran (\sa_snapshot[5][50] , \sa_snapshot[5].r.part1[18] );
tran (\sa_snapshot[5][50] , \sa_snapshot[5].f.unused[0] );
tran (\sa_snapshot[5][51] , \sa_snapshot[5].r.part1[19] );
tran (\sa_snapshot[5][51] , \sa_snapshot[5].f.unused[1] );
tran (\sa_snapshot[5][52] , \sa_snapshot[5].r.part1[20] );
tran (\sa_snapshot[5][52] , \sa_snapshot[5].f.unused[2] );
tran (\sa_snapshot[5][53] , \sa_snapshot[5].r.part1[21] );
tran (\sa_snapshot[5][53] , \sa_snapshot[5].f.unused[3] );
tran (\sa_snapshot[5][54] , \sa_snapshot[5].r.part1[22] );
tran (\sa_snapshot[5][54] , \sa_snapshot[5].f.unused[4] );
tran (\sa_snapshot[5][55] , \sa_snapshot[5].r.part1[23] );
tran (\sa_snapshot[5][55] , \sa_snapshot[5].f.unused[5] );
tran (\sa_snapshot[5][56] , \sa_snapshot[5].r.part1[24] );
tran (\sa_snapshot[5][56] , \sa_snapshot[5].f.unused[6] );
tran (\sa_snapshot[5][57] , \sa_snapshot[5].r.part1[25] );
tran (\sa_snapshot[5][57] , \sa_snapshot[5].f.unused[7] );
tran (\sa_snapshot[5][58] , \sa_snapshot[5].r.part1[26] );
tran (\sa_snapshot[5][58] , \sa_snapshot[5].f.unused[8] );
tran (\sa_snapshot[5][59] , \sa_snapshot[5].r.part1[27] );
tran (\sa_snapshot[5][59] , \sa_snapshot[5].f.unused[9] );
tran (\sa_snapshot[5][60] , \sa_snapshot[5].r.part1[28] );
tran (\sa_snapshot[5][60] , \sa_snapshot[5].f.unused[10] );
tran (\sa_snapshot[5][61] , \sa_snapshot[5].r.part1[29] );
tran (\sa_snapshot[5][61] , \sa_snapshot[5].f.unused[11] );
tran (\sa_snapshot[5][62] , \sa_snapshot[5].r.part1[30] );
tran (\sa_snapshot[5][62] , \sa_snapshot[5].f.unused[12] );
tran (\sa_snapshot[5][63] , \sa_snapshot[5].r.part1[31] );
tran (\sa_snapshot[5][63] , \sa_snapshot[5].f.unused[13] );
tran (\sa_snapshot[6][0] , \sa_snapshot[6].r.part0[0] );
tran (\sa_snapshot[6][0] , \sa_snapshot[6].f.lower[0] );
tran (\sa_snapshot[6][1] , \sa_snapshot[6].r.part0[1] );
tran (\sa_snapshot[6][1] , \sa_snapshot[6].f.lower[1] );
tran (\sa_snapshot[6][2] , \sa_snapshot[6].r.part0[2] );
tran (\sa_snapshot[6][2] , \sa_snapshot[6].f.lower[2] );
tran (\sa_snapshot[6][3] , \sa_snapshot[6].r.part0[3] );
tran (\sa_snapshot[6][3] , \sa_snapshot[6].f.lower[3] );
tran (\sa_snapshot[6][4] , \sa_snapshot[6].r.part0[4] );
tran (\sa_snapshot[6][4] , \sa_snapshot[6].f.lower[4] );
tran (\sa_snapshot[6][5] , \sa_snapshot[6].r.part0[5] );
tran (\sa_snapshot[6][5] , \sa_snapshot[6].f.lower[5] );
tran (\sa_snapshot[6][6] , \sa_snapshot[6].r.part0[6] );
tran (\sa_snapshot[6][6] , \sa_snapshot[6].f.lower[6] );
tran (\sa_snapshot[6][7] , \sa_snapshot[6].r.part0[7] );
tran (\sa_snapshot[6][7] , \sa_snapshot[6].f.lower[7] );
tran (\sa_snapshot[6][8] , \sa_snapshot[6].r.part0[8] );
tran (\sa_snapshot[6][8] , \sa_snapshot[6].f.lower[8] );
tran (\sa_snapshot[6][9] , \sa_snapshot[6].r.part0[9] );
tran (\sa_snapshot[6][9] , \sa_snapshot[6].f.lower[9] );
tran (\sa_snapshot[6][10] , \sa_snapshot[6].r.part0[10] );
tran (\sa_snapshot[6][10] , \sa_snapshot[6].f.lower[10] );
tran (\sa_snapshot[6][11] , \sa_snapshot[6].r.part0[11] );
tran (\sa_snapshot[6][11] , \sa_snapshot[6].f.lower[11] );
tran (\sa_snapshot[6][12] , \sa_snapshot[6].r.part0[12] );
tran (\sa_snapshot[6][12] , \sa_snapshot[6].f.lower[12] );
tran (\sa_snapshot[6][13] , \sa_snapshot[6].r.part0[13] );
tran (\sa_snapshot[6][13] , \sa_snapshot[6].f.lower[13] );
tran (\sa_snapshot[6][14] , \sa_snapshot[6].r.part0[14] );
tran (\sa_snapshot[6][14] , \sa_snapshot[6].f.lower[14] );
tran (\sa_snapshot[6][15] , \sa_snapshot[6].r.part0[15] );
tran (\sa_snapshot[6][15] , \sa_snapshot[6].f.lower[15] );
tran (\sa_snapshot[6][16] , \sa_snapshot[6].r.part0[16] );
tran (\sa_snapshot[6][16] , \sa_snapshot[6].f.lower[16] );
tran (\sa_snapshot[6][17] , \sa_snapshot[6].r.part0[17] );
tran (\sa_snapshot[6][17] , \sa_snapshot[6].f.lower[17] );
tran (\sa_snapshot[6][18] , \sa_snapshot[6].r.part0[18] );
tran (\sa_snapshot[6][18] , \sa_snapshot[6].f.lower[18] );
tran (\sa_snapshot[6][19] , \sa_snapshot[6].r.part0[19] );
tran (\sa_snapshot[6][19] , \sa_snapshot[6].f.lower[19] );
tran (\sa_snapshot[6][20] , \sa_snapshot[6].r.part0[20] );
tran (\sa_snapshot[6][20] , \sa_snapshot[6].f.lower[20] );
tran (\sa_snapshot[6][21] , \sa_snapshot[6].r.part0[21] );
tran (\sa_snapshot[6][21] , \sa_snapshot[6].f.lower[21] );
tran (\sa_snapshot[6][22] , \sa_snapshot[6].r.part0[22] );
tran (\sa_snapshot[6][22] , \sa_snapshot[6].f.lower[22] );
tran (\sa_snapshot[6][23] , \sa_snapshot[6].r.part0[23] );
tran (\sa_snapshot[6][23] , \sa_snapshot[6].f.lower[23] );
tran (\sa_snapshot[6][24] , \sa_snapshot[6].r.part0[24] );
tran (\sa_snapshot[6][24] , \sa_snapshot[6].f.lower[24] );
tran (\sa_snapshot[6][25] , \sa_snapshot[6].r.part0[25] );
tran (\sa_snapshot[6][25] , \sa_snapshot[6].f.lower[25] );
tran (\sa_snapshot[6][26] , \sa_snapshot[6].r.part0[26] );
tran (\sa_snapshot[6][26] , \sa_snapshot[6].f.lower[26] );
tran (\sa_snapshot[6][27] , \sa_snapshot[6].r.part0[27] );
tran (\sa_snapshot[6][27] , \sa_snapshot[6].f.lower[27] );
tran (\sa_snapshot[6][28] , \sa_snapshot[6].r.part0[28] );
tran (\sa_snapshot[6][28] , \sa_snapshot[6].f.lower[28] );
tran (\sa_snapshot[6][29] , \sa_snapshot[6].r.part0[29] );
tran (\sa_snapshot[6][29] , \sa_snapshot[6].f.lower[29] );
tran (\sa_snapshot[6][30] , \sa_snapshot[6].r.part0[30] );
tran (\sa_snapshot[6][30] , \sa_snapshot[6].f.lower[30] );
tran (\sa_snapshot[6][31] , \sa_snapshot[6].r.part0[31] );
tran (\sa_snapshot[6][31] , \sa_snapshot[6].f.lower[31] );
tran (\sa_snapshot[6][32] , \sa_snapshot[6].r.part1[0] );
tran (\sa_snapshot[6][32] , \sa_snapshot[6].f.upper[0] );
tran (\sa_snapshot[6][33] , \sa_snapshot[6].r.part1[1] );
tran (\sa_snapshot[6][33] , \sa_snapshot[6].f.upper[1] );
tran (\sa_snapshot[6][34] , \sa_snapshot[6].r.part1[2] );
tran (\sa_snapshot[6][34] , \sa_snapshot[6].f.upper[2] );
tran (\sa_snapshot[6][35] , \sa_snapshot[6].r.part1[3] );
tran (\sa_snapshot[6][35] , \sa_snapshot[6].f.upper[3] );
tran (\sa_snapshot[6][36] , \sa_snapshot[6].r.part1[4] );
tran (\sa_snapshot[6][36] , \sa_snapshot[6].f.upper[4] );
tran (\sa_snapshot[6][37] , \sa_snapshot[6].r.part1[5] );
tran (\sa_snapshot[6][37] , \sa_snapshot[6].f.upper[5] );
tran (\sa_snapshot[6][38] , \sa_snapshot[6].r.part1[6] );
tran (\sa_snapshot[6][38] , \sa_snapshot[6].f.upper[6] );
tran (\sa_snapshot[6][39] , \sa_snapshot[6].r.part1[7] );
tran (\sa_snapshot[6][39] , \sa_snapshot[6].f.upper[7] );
tran (\sa_snapshot[6][40] , \sa_snapshot[6].r.part1[8] );
tran (\sa_snapshot[6][40] , \sa_snapshot[6].f.upper[8] );
tran (\sa_snapshot[6][41] , \sa_snapshot[6].r.part1[9] );
tran (\sa_snapshot[6][41] , \sa_snapshot[6].f.upper[9] );
tran (\sa_snapshot[6][42] , \sa_snapshot[6].r.part1[10] );
tran (\sa_snapshot[6][42] , \sa_snapshot[6].f.upper[10] );
tran (\sa_snapshot[6][43] , \sa_snapshot[6].r.part1[11] );
tran (\sa_snapshot[6][43] , \sa_snapshot[6].f.upper[11] );
tran (\sa_snapshot[6][44] , \sa_snapshot[6].r.part1[12] );
tran (\sa_snapshot[6][44] , \sa_snapshot[6].f.upper[12] );
tran (\sa_snapshot[6][45] , \sa_snapshot[6].r.part1[13] );
tran (\sa_snapshot[6][45] , \sa_snapshot[6].f.upper[13] );
tran (\sa_snapshot[6][46] , \sa_snapshot[6].r.part1[14] );
tran (\sa_snapshot[6][46] , \sa_snapshot[6].f.upper[14] );
tran (\sa_snapshot[6][47] , \sa_snapshot[6].r.part1[15] );
tran (\sa_snapshot[6][47] , \sa_snapshot[6].f.upper[15] );
tran (\sa_snapshot[6][48] , \sa_snapshot[6].r.part1[16] );
tran (\sa_snapshot[6][48] , \sa_snapshot[6].f.upper[16] );
tran (\sa_snapshot[6][49] , \sa_snapshot[6].r.part1[17] );
tran (\sa_snapshot[6][49] , \sa_snapshot[6].f.upper[17] );
tran (\sa_snapshot[6][50] , \sa_snapshot[6].r.part1[18] );
tran (\sa_snapshot[6][50] , \sa_snapshot[6].f.unused[0] );
tran (\sa_snapshot[6][51] , \sa_snapshot[6].r.part1[19] );
tran (\sa_snapshot[6][51] , \sa_snapshot[6].f.unused[1] );
tran (\sa_snapshot[6][52] , \sa_snapshot[6].r.part1[20] );
tran (\sa_snapshot[6][52] , \sa_snapshot[6].f.unused[2] );
tran (\sa_snapshot[6][53] , \sa_snapshot[6].r.part1[21] );
tran (\sa_snapshot[6][53] , \sa_snapshot[6].f.unused[3] );
tran (\sa_snapshot[6][54] , \sa_snapshot[6].r.part1[22] );
tran (\sa_snapshot[6][54] , \sa_snapshot[6].f.unused[4] );
tran (\sa_snapshot[6][55] , \sa_snapshot[6].r.part1[23] );
tran (\sa_snapshot[6][55] , \sa_snapshot[6].f.unused[5] );
tran (\sa_snapshot[6][56] , \sa_snapshot[6].r.part1[24] );
tran (\sa_snapshot[6][56] , \sa_snapshot[6].f.unused[6] );
tran (\sa_snapshot[6][57] , \sa_snapshot[6].r.part1[25] );
tran (\sa_snapshot[6][57] , \sa_snapshot[6].f.unused[7] );
tran (\sa_snapshot[6][58] , \sa_snapshot[6].r.part1[26] );
tran (\sa_snapshot[6][58] , \sa_snapshot[6].f.unused[8] );
tran (\sa_snapshot[6][59] , \sa_snapshot[6].r.part1[27] );
tran (\sa_snapshot[6][59] , \sa_snapshot[6].f.unused[9] );
tran (\sa_snapshot[6][60] , \sa_snapshot[6].r.part1[28] );
tran (\sa_snapshot[6][60] , \sa_snapshot[6].f.unused[10] );
tran (\sa_snapshot[6][61] , \sa_snapshot[6].r.part1[29] );
tran (\sa_snapshot[6][61] , \sa_snapshot[6].f.unused[11] );
tran (\sa_snapshot[6][62] , \sa_snapshot[6].r.part1[30] );
tran (\sa_snapshot[6][62] , \sa_snapshot[6].f.unused[12] );
tran (\sa_snapshot[6][63] , \sa_snapshot[6].r.part1[31] );
tran (\sa_snapshot[6][63] , \sa_snapshot[6].f.unused[13] );
tran (\sa_snapshot[7][0] , \sa_snapshot[7].r.part0[0] );
tran (\sa_snapshot[7][0] , \sa_snapshot[7].f.lower[0] );
tran (\sa_snapshot[7][1] , \sa_snapshot[7].r.part0[1] );
tran (\sa_snapshot[7][1] , \sa_snapshot[7].f.lower[1] );
tran (\sa_snapshot[7][2] , \sa_snapshot[7].r.part0[2] );
tran (\sa_snapshot[7][2] , \sa_snapshot[7].f.lower[2] );
tran (\sa_snapshot[7][3] , \sa_snapshot[7].r.part0[3] );
tran (\sa_snapshot[7][3] , \sa_snapshot[7].f.lower[3] );
tran (\sa_snapshot[7][4] , \sa_snapshot[7].r.part0[4] );
tran (\sa_snapshot[7][4] , \sa_snapshot[7].f.lower[4] );
tran (\sa_snapshot[7][5] , \sa_snapshot[7].r.part0[5] );
tran (\sa_snapshot[7][5] , \sa_snapshot[7].f.lower[5] );
tran (\sa_snapshot[7][6] , \sa_snapshot[7].r.part0[6] );
tran (\sa_snapshot[7][6] , \sa_snapshot[7].f.lower[6] );
tran (\sa_snapshot[7][7] , \sa_snapshot[7].r.part0[7] );
tran (\sa_snapshot[7][7] , \sa_snapshot[7].f.lower[7] );
tran (\sa_snapshot[7][8] , \sa_snapshot[7].r.part0[8] );
tran (\sa_snapshot[7][8] , \sa_snapshot[7].f.lower[8] );
tran (\sa_snapshot[7][9] , \sa_snapshot[7].r.part0[9] );
tran (\sa_snapshot[7][9] , \sa_snapshot[7].f.lower[9] );
tran (\sa_snapshot[7][10] , \sa_snapshot[7].r.part0[10] );
tran (\sa_snapshot[7][10] , \sa_snapshot[7].f.lower[10] );
tran (\sa_snapshot[7][11] , \sa_snapshot[7].r.part0[11] );
tran (\sa_snapshot[7][11] , \sa_snapshot[7].f.lower[11] );
tran (\sa_snapshot[7][12] , \sa_snapshot[7].r.part0[12] );
tran (\sa_snapshot[7][12] , \sa_snapshot[7].f.lower[12] );
tran (\sa_snapshot[7][13] , \sa_snapshot[7].r.part0[13] );
tran (\sa_snapshot[7][13] , \sa_snapshot[7].f.lower[13] );
tran (\sa_snapshot[7][14] , \sa_snapshot[7].r.part0[14] );
tran (\sa_snapshot[7][14] , \sa_snapshot[7].f.lower[14] );
tran (\sa_snapshot[7][15] , \sa_snapshot[7].r.part0[15] );
tran (\sa_snapshot[7][15] , \sa_snapshot[7].f.lower[15] );
tran (\sa_snapshot[7][16] , \sa_snapshot[7].r.part0[16] );
tran (\sa_snapshot[7][16] , \sa_snapshot[7].f.lower[16] );
tran (\sa_snapshot[7][17] , \sa_snapshot[7].r.part0[17] );
tran (\sa_snapshot[7][17] , \sa_snapshot[7].f.lower[17] );
tran (\sa_snapshot[7][18] , \sa_snapshot[7].r.part0[18] );
tran (\sa_snapshot[7][18] , \sa_snapshot[7].f.lower[18] );
tran (\sa_snapshot[7][19] , \sa_snapshot[7].r.part0[19] );
tran (\sa_snapshot[7][19] , \sa_snapshot[7].f.lower[19] );
tran (\sa_snapshot[7][20] , \sa_snapshot[7].r.part0[20] );
tran (\sa_snapshot[7][20] , \sa_snapshot[7].f.lower[20] );
tran (\sa_snapshot[7][21] , \sa_snapshot[7].r.part0[21] );
tran (\sa_snapshot[7][21] , \sa_snapshot[7].f.lower[21] );
tran (\sa_snapshot[7][22] , \sa_snapshot[7].r.part0[22] );
tran (\sa_snapshot[7][22] , \sa_snapshot[7].f.lower[22] );
tran (\sa_snapshot[7][23] , \sa_snapshot[7].r.part0[23] );
tran (\sa_snapshot[7][23] , \sa_snapshot[7].f.lower[23] );
tran (\sa_snapshot[7][24] , \sa_snapshot[7].r.part0[24] );
tran (\sa_snapshot[7][24] , \sa_snapshot[7].f.lower[24] );
tran (\sa_snapshot[7][25] , \sa_snapshot[7].r.part0[25] );
tran (\sa_snapshot[7][25] , \sa_snapshot[7].f.lower[25] );
tran (\sa_snapshot[7][26] , \sa_snapshot[7].r.part0[26] );
tran (\sa_snapshot[7][26] , \sa_snapshot[7].f.lower[26] );
tran (\sa_snapshot[7][27] , \sa_snapshot[7].r.part0[27] );
tran (\sa_snapshot[7][27] , \sa_snapshot[7].f.lower[27] );
tran (\sa_snapshot[7][28] , \sa_snapshot[7].r.part0[28] );
tran (\sa_snapshot[7][28] , \sa_snapshot[7].f.lower[28] );
tran (\sa_snapshot[7][29] , \sa_snapshot[7].r.part0[29] );
tran (\sa_snapshot[7][29] , \sa_snapshot[7].f.lower[29] );
tran (\sa_snapshot[7][30] , \sa_snapshot[7].r.part0[30] );
tran (\sa_snapshot[7][30] , \sa_snapshot[7].f.lower[30] );
tran (\sa_snapshot[7][31] , \sa_snapshot[7].r.part0[31] );
tran (\sa_snapshot[7][31] , \sa_snapshot[7].f.lower[31] );
tran (\sa_snapshot[7][32] , \sa_snapshot[7].r.part1[0] );
tran (\sa_snapshot[7][32] , \sa_snapshot[7].f.upper[0] );
tran (\sa_snapshot[7][33] , \sa_snapshot[7].r.part1[1] );
tran (\sa_snapshot[7][33] , \sa_snapshot[7].f.upper[1] );
tran (\sa_snapshot[7][34] , \sa_snapshot[7].r.part1[2] );
tran (\sa_snapshot[7][34] , \sa_snapshot[7].f.upper[2] );
tran (\sa_snapshot[7][35] , \sa_snapshot[7].r.part1[3] );
tran (\sa_snapshot[7][35] , \sa_snapshot[7].f.upper[3] );
tran (\sa_snapshot[7][36] , \sa_snapshot[7].r.part1[4] );
tran (\sa_snapshot[7][36] , \sa_snapshot[7].f.upper[4] );
tran (\sa_snapshot[7][37] , \sa_snapshot[7].r.part1[5] );
tran (\sa_snapshot[7][37] , \sa_snapshot[7].f.upper[5] );
tran (\sa_snapshot[7][38] , \sa_snapshot[7].r.part1[6] );
tran (\sa_snapshot[7][38] , \sa_snapshot[7].f.upper[6] );
tran (\sa_snapshot[7][39] , \sa_snapshot[7].r.part1[7] );
tran (\sa_snapshot[7][39] , \sa_snapshot[7].f.upper[7] );
tran (\sa_snapshot[7][40] , \sa_snapshot[7].r.part1[8] );
tran (\sa_snapshot[7][40] , \sa_snapshot[7].f.upper[8] );
tran (\sa_snapshot[7][41] , \sa_snapshot[7].r.part1[9] );
tran (\sa_snapshot[7][41] , \sa_snapshot[7].f.upper[9] );
tran (\sa_snapshot[7][42] , \sa_snapshot[7].r.part1[10] );
tran (\sa_snapshot[7][42] , \sa_snapshot[7].f.upper[10] );
tran (\sa_snapshot[7][43] , \sa_snapshot[7].r.part1[11] );
tran (\sa_snapshot[7][43] , \sa_snapshot[7].f.upper[11] );
tran (\sa_snapshot[7][44] , \sa_snapshot[7].r.part1[12] );
tran (\sa_snapshot[7][44] , \sa_snapshot[7].f.upper[12] );
tran (\sa_snapshot[7][45] , \sa_snapshot[7].r.part1[13] );
tran (\sa_snapshot[7][45] , \sa_snapshot[7].f.upper[13] );
tran (\sa_snapshot[7][46] , \sa_snapshot[7].r.part1[14] );
tran (\sa_snapshot[7][46] , \sa_snapshot[7].f.upper[14] );
tran (\sa_snapshot[7][47] , \sa_snapshot[7].r.part1[15] );
tran (\sa_snapshot[7][47] , \sa_snapshot[7].f.upper[15] );
tran (\sa_snapshot[7][48] , \sa_snapshot[7].r.part1[16] );
tran (\sa_snapshot[7][48] , \sa_snapshot[7].f.upper[16] );
tran (\sa_snapshot[7][49] , \sa_snapshot[7].r.part1[17] );
tran (\sa_snapshot[7][49] , \sa_snapshot[7].f.upper[17] );
tran (\sa_snapshot[7][50] , \sa_snapshot[7].r.part1[18] );
tran (\sa_snapshot[7][50] , \sa_snapshot[7].f.unused[0] );
tran (\sa_snapshot[7][51] , \sa_snapshot[7].r.part1[19] );
tran (\sa_snapshot[7][51] , \sa_snapshot[7].f.unused[1] );
tran (\sa_snapshot[7][52] , \sa_snapshot[7].r.part1[20] );
tran (\sa_snapshot[7][52] , \sa_snapshot[7].f.unused[2] );
tran (\sa_snapshot[7][53] , \sa_snapshot[7].r.part1[21] );
tran (\sa_snapshot[7][53] , \sa_snapshot[7].f.unused[3] );
tran (\sa_snapshot[7][54] , \sa_snapshot[7].r.part1[22] );
tran (\sa_snapshot[7][54] , \sa_snapshot[7].f.unused[4] );
tran (\sa_snapshot[7][55] , \sa_snapshot[7].r.part1[23] );
tran (\sa_snapshot[7][55] , \sa_snapshot[7].f.unused[5] );
tran (\sa_snapshot[7][56] , \sa_snapshot[7].r.part1[24] );
tran (\sa_snapshot[7][56] , \sa_snapshot[7].f.unused[6] );
tran (\sa_snapshot[7][57] , \sa_snapshot[7].r.part1[25] );
tran (\sa_snapshot[7][57] , \sa_snapshot[7].f.unused[7] );
tran (\sa_snapshot[7][58] , \sa_snapshot[7].r.part1[26] );
tran (\sa_snapshot[7][58] , \sa_snapshot[7].f.unused[8] );
tran (\sa_snapshot[7][59] , \sa_snapshot[7].r.part1[27] );
tran (\sa_snapshot[7][59] , \sa_snapshot[7].f.unused[9] );
tran (\sa_snapshot[7][60] , \sa_snapshot[7].r.part1[28] );
tran (\sa_snapshot[7][60] , \sa_snapshot[7].f.unused[10] );
tran (\sa_snapshot[7][61] , \sa_snapshot[7].r.part1[29] );
tran (\sa_snapshot[7][61] , \sa_snapshot[7].f.unused[11] );
tran (\sa_snapshot[7][62] , \sa_snapshot[7].r.part1[30] );
tran (\sa_snapshot[7][62] , \sa_snapshot[7].f.unused[12] );
tran (\sa_snapshot[7][63] , \sa_snapshot[7].r.part1[31] );
tran (\sa_snapshot[7][63] , \sa_snapshot[7].f.unused[13] );
tran (\sa_snapshot[8][0] , \sa_snapshot[8].r.part0[0] );
tran (\sa_snapshot[8][0] , \sa_snapshot[8].f.lower[0] );
tran (\sa_snapshot[8][1] , \sa_snapshot[8].r.part0[1] );
tran (\sa_snapshot[8][1] , \sa_snapshot[8].f.lower[1] );
tran (\sa_snapshot[8][2] , \sa_snapshot[8].r.part0[2] );
tran (\sa_snapshot[8][2] , \sa_snapshot[8].f.lower[2] );
tran (\sa_snapshot[8][3] , \sa_snapshot[8].r.part0[3] );
tran (\sa_snapshot[8][3] , \sa_snapshot[8].f.lower[3] );
tran (\sa_snapshot[8][4] , \sa_snapshot[8].r.part0[4] );
tran (\sa_snapshot[8][4] , \sa_snapshot[8].f.lower[4] );
tran (\sa_snapshot[8][5] , \sa_snapshot[8].r.part0[5] );
tran (\sa_snapshot[8][5] , \sa_snapshot[8].f.lower[5] );
tran (\sa_snapshot[8][6] , \sa_snapshot[8].r.part0[6] );
tran (\sa_snapshot[8][6] , \sa_snapshot[8].f.lower[6] );
tran (\sa_snapshot[8][7] , \sa_snapshot[8].r.part0[7] );
tran (\sa_snapshot[8][7] , \sa_snapshot[8].f.lower[7] );
tran (\sa_snapshot[8][8] , \sa_snapshot[8].r.part0[8] );
tran (\sa_snapshot[8][8] , \sa_snapshot[8].f.lower[8] );
tran (\sa_snapshot[8][9] , \sa_snapshot[8].r.part0[9] );
tran (\sa_snapshot[8][9] , \sa_snapshot[8].f.lower[9] );
tran (\sa_snapshot[8][10] , \sa_snapshot[8].r.part0[10] );
tran (\sa_snapshot[8][10] , \sa_snapshot[8].f.lower[10] );
tran (\sa_snapshot[8][11] , \sa_snapshot[8].r.part0[11] );
tran (\sa_snapshot[8][11] , \sa_snapshot[8].f.lower[11] );
tran (\sa_snapshot[8][12] , \sa_snapshot[8].r.part0[12] );
tran (\sa_snapshot[8][12] , \sa_snapshot[8].f.lower[12] );
tran (\sa_snapshot[8][13] , \sa_snapshot[8].r.part0[13] );
tran (\sa_snapshot[8][13] , \sa_snapshot[8].f.lower[13] );
tran (\sa_snapshot[8][14] , \sa_snapshot[8].r.part0[14] );
tran (\sa_snapshot[8][14] , \sa_snapshot[8].f.lower[14] );
tran (\sa_snapshot[8][15] , \sa_snapshot[8].r.part0[15] );
tran (\sa_snapshot[8][15] , \sa_snapshot[8].f.lower[15] );
tran (\sa_snapshot[8][16] , \sa_snapshot[8].r.part0[16] );
tran (\sa_snapshot[8][16] , \sa_snapshot[8].f.lower[16] );
tran (\sa_snapshot[8][17] , \sa_snapshot[8].r.part0[17] );
tran (\sa_snapshot[8][17] , \sa_snapshot[8].f.lower[17] );
tran (\sa_snapshot[8][18] , \sa_snapshot[8].r.part0[18] );
tran (\sa_snapshot[8][18] , \sa_snapshot[8].f.lower[18] );
tran (\sa_snapshot[8][19] , \sa_snapshot[8].r.part0[19] );
tran (\sa_snapshot[8][19] , \sa_snapshot[8].f.lower[19] );
tran (\sa_snapshot[8][20] , \sa_snapshot[8].r.part0[20] );
tran (\sa_snapshot[8][20] , \sa_snapshot[8].f.lower[20] );
tran (\sa_snapshot[8][21] , \sa_snapshot[8].r.part0[21] );
tran (\sa_snapshot[8][21] , \sa_snapshot[8].f.lower[21] );
tran (\sa_snapshot[8][22] , \sa_snapshot[8].r.part0[22] );
tran (\sa_snapshot[8][22] , \sa_snapshot[8].f.lower[22] );
tran (\sa_snapshot[8][23] , \sa_snapshot[8].r.part0[23] );
tran (\sa_snapshot[8][23] , \sa_snapshot[8].f.lower[23] );
tran (\sa_snapshot[8][24] , \sa_snapshot[8].r.part0[24] );
tran (\sa_snapshot[8][24] , \sa_snapshot[8].f.lower[24] );
tran (\sa_snapshot[8][25] , \sa_snapshot[8].r.part0[25] );
tran (\sa_snapshot[8][25] , \sa_snapshot[8].f.lower[25] );
tran (\sa_snapshot[8][26] , \sa_snapshot[8].r.part0[26] );
tran (\sa_snapshot[8][26] , \sa_snapshot[8].f.lower[26] );
tran (\sa_snapshot[8][27] , \sa_snapshot[8].r.part0[27] );
tran (\sa_snapshot[8][27] , \sa_snapshot[8].f.lower[27] );
tran (\sa_snapshot[8][28] , \sa_snapshot[8].r.part0[28] );
tran (\sa_snapshot[8][28] , \sa_snapshot[8].f.lower[28] );
tran (\sa_snapshot[8][29] , \sa_snapshot[8].r.part0[29] );
tran (\sa_snapshot[8][29] , \sa_snapshot[8].f.lower[29] );
tran (\sa_snapshot[8][30] , \sa_snapshot[8].r.part0[30] );
tran (\sa_snapshot[8][30] , \sa_snapshot[8].f.lower[30] );
tran (\sa_snapshot[8][31] , \sa_snapshot[8].r.part0[31] );
tran (\sa_snapshot[8][31] , \sa_snapshot[8].f.lower[31] );
tran (\sa_snapshot[8][32] , \sa_snapshot[8].r.part1[0] );
tran (\sa_snapshot[8][32] , \sa_snapshot[8].f.upper[0] );
tran (\sa_snapshot[8][33] , \sa_snapshot[8].r.part1[1] );
tran (\sa_snapshot[8][33] , \sa_snapshot[8].f.upper[1] );
tran (\sa_snapshot[8][34] , \sa_snapshot[8].r.part1[2] );
tran (\sa_snapshot[8][34] , \sa_snapshot[8].f.upper[2] );
tran (\sa_snapshot[8][35] , \sa_snapshot[8].r.part1[3] );
tran (\sa_snapshot[8][35] , \sa_snapshot[8].f.upper[3] );
tran (\sa_snapshot[8][36] , \sa_snapshot[8].r.part1[4] );
tran (\sa_snapshot[8][36] , \sa_snapshot[8].f.upper[4] );
tran (\sa_snapshot[8][37] , \sa_snapshot[8].r.part1[5] );
tran (\sa_snapshot[8][37] , \sa_snapshot[8].f.upper[5] );
tran (\sa_snapshot[8][38] , \sa_snapshot[8].r.part1[6] );
tran (\sa_snapshot[8][38] , \sa_snapshot[8].f.upper[6] );
tran (\sa_snapshot[8][39] , \sa_snapshot[8].r.part1[7] );
tran (\sa_snapshot[8][39] , \sa_snapshot[8].f.upper[7] );
tran (\sa_snapshot[8][40] , \sa_snapshot[8].r.part1[8] );
tran (\sa_snapshot[8][40] , \sa_snapshot[8].f.upper[8] );
tran (\sa_snapshot[8][41] , \sa_snapshot[8].r.part1[9] );
tran (\sa_snapshot[8][41] , \sa_snapshot[8].f.upper[9] );
tran (\sa_snapshot[8][42] , \sa_snapshot[8].r.part1[10] );
tran (\sa_snapshot[8][42] , \sa_snapshot[8].f.upper[10] );
tran (\sa_snapshot[8][43] , \sa_snapshot[8].r.part1[11] );
tran (\sa_snapshot[8][43] , \sa_snapshot[8].f.upper[11] );
tran (\sa_snapshot[8][44] , \sa_snapshot[8].r.part1[12] );
tran (\sa_snapshot[8][44] , \sa_snapshot[8].f.upper[12] );
tran (\sa_snapshot[8][45] , \sa_snapshot[8].r.part1[13] );
tran (\sa_snapshot[8][45] , \sa_snapshot[8].f.upper[13] );
tran (\sa_snapshot[8][46] , \sa_snapshot[8].r.part1[14] );
tran (\sa_snapshot[8][46] , \sa_snapshot[8].f.upper[14] );
tran (\sa_snapshot[8][47] , \sa_snapshot[8].r.part1[15] );
tran (\sa_snapshot[8][47] , \sa_snapshot[8].f.upper[15] );
tran (\sa_snapshot[8][48] , \sa_snapshot[8].r.part1[16] );
tran (\sa_snapshot[8][48] , \sa_snapshot[8].f.upper[16] );
tran (\sa_snapshot[8][49] , \sa_snapshot[8].r.part1[17] );
tran (\sa_snapshot[8][49] , \sa_snapshot[8].f.upper[17] );
tran (\sa_snapshot[8][50] , \sa_snapshot[8].r.part1[18] );
tran (\sa_snapshot[8][50] , \sa_snapshot[8].f.unused[0] );
tran (\sa_snapshot[8][51] , \sa_snapshot[8].r.part1[19] );
tran (\sa_snapshot[8][51] , \sa_snapshot[8].f.unused[1] );
tran (\sa_snapshot[8][52] , \sa_snapshot[8].r.part1[20] );
tran (\sa_snapshot[8][52] , \sa_snapshot[8].f.unused[2] );
tran (\sa_snapshot[8][53] , \sa_snapshot[8].r.part1[21] );
tran (\sa_snapshot[8][53] , \sa_snapshot[8].f.unused[3] );
tran (\sa_snapshot[8][54] , \sa_snapshot[8].r.part1[22] );
tran (\sa_snapshot[8][54] , \sa_snapshot[8].f.unused[4] );
tran (\sa_snapshot[8][55] , \sa_snapshot[8].r.part1[23] );
tran (\sa_snapshot[8][55] , \sa_snapshot[8].f.unused[5] );
tran (\sa_snapshot[8][56] , \sa_snapshot[8].r.part1[24] );
tran (\sa_snapshot[8][56] , \sa_snapshot[8].f.unused[6] );
tran (\sa_snapshot[8][57] , \sa_snapshot[8].r.part1[25] );
tran (\sa_snapshot[8][57] , \sa_snapshot[8].f.unused[7] );
tran (\sa_snapshot[8][58] , \sa_snapshot[8].r.part1[26] );
tran (\sa_snapshot[8][58] , \sa_snapshot[8].f.unused[8] );
tran (\sa_snapshot[8][59] , \sa_snapshot[8].r.part1[27] );
tran (\sa_snapshot[8][59] , \sa_snapshot[8].f.unused[9] );
tran (\sa_snapshot[8][60] , \sa_snapshot[8].r.part1[28] );
tran (\sa_snapshot[8][60] , \sa_snapshot[8].f.unused[10] );
tran (\sa_snapshot[8][61] , \sa_snapshot[8].r.part1[29] );
tran (\sa_snapshot[8][61] , \sa_snapshot[8].f.unused[11] );
tran (\sa_snapshot[8][62] , \sa_snapshot[8].r.part1[30] );
tran (\sa_snapshot[8][62] , \sa_snapshot[8].f.unused[12] );
tran (\sa_snapshot[8][63] , \sa_snapshot[8].r.part1[31] );
tran (\sa_snapshot[8][63] , \sa_snapshot[8].f.unused[13] );
tran (\sa_snapshot[9][0] , \sa_snapshot[9].r.part0[0] );
tran (\sa_snapshot[9][0] , \sa_snapshot[9].f.lower[0] );
tran (\sa_snapshot[9][1] , \sa_snapshot[9].r.part0[1] );
tran (\sa_snapshot[9][1] , \sa_snapshot[9].f.lower[1] );
tran (\sa_snapshot[9][2] , \sa_snapshot[9].r.part0[2] );
tran (\sa_snapshot[9][2] , \sa_snapshot[9].f.lower[2] );
tran (\sa_snapshot[9][3] , \sa_snapshot[9].r.part0[3] );
tran (\sa_snapshot[9][3] , \sa_snapshot[9].f.lower[3] );
tran (\sa_snapshot[9][4] , \sa_snapshot[9].r.part0[4] );
tran (\sa_snapshot[9][4] , \sa_snapshot[9].f.lower[4] );
tran (\sa_snapshot[9][5] , \sa_snapshot[9].r.part0[5] );
tran (\sa_snapshot[9][5] , \sa_snapshot[9].f.lower[5] );
tran (\sa_snapshot[9][6] , \sa_snapshot[9].r.part0[6] );
tran (\sa_snapshot[9][6] , \sa_snapshot[9].f.lower[6] );
tran (\sa_snapshot[9][7] , \sa_snapshot[9].r.part0[7] );
tran (\sa_snapshot[9][7] , \sa_snapshot[9].f.lower[7] );
tran (\sa_snapshot[9][8] , \sa_snapshot[9].r.part0[8] );
tran (\sa_snapshot[9][8] , \sa_snapshot[9].f.lower[8] );
tran (\sa_snapshot[9][9] , \sa_snapshot[9].r.part0[9] );
tran (\sa_snapshot[9][9] , \sa_snapshot[9].f.lower[9] );
tran (\sa_snapshot[9][10] , \sa_snapshot[9].r.part0[10] );
tran (\sa_snapshot[9][10] , \sa_snapshot[9].f.lower[10] );
tran (\sa_snapshot[9][11] , \sa_snapshot[9].r.part0[11] );
tran (\sa_snapshot[9][11] , \sa_snapshot[9].f.lower[11] );
tran (\sa_snapshot[9][12] , \sa_snapshot[9].r.part0[12] );
tran (\sa_snapshot[9][12] , \sa_snapshot[9].f.lower[12] );
tran (\sa_snapshot[9][13] , \sa_snapshot[9].r.part0[13] );
tran (\sa_snapshot[9][13] , \sa_snapshot[9].f.lower[13] );
tran (\sa_snapshot[9][14] , \sa_snapshot[9].r.part0[14] );
tran (\sa_snapshot[9][14] , \sa_snapshot[9].f.lower[14] );
tran (\sa_snapshot[9][15] , \sa_snapshot[9].r.part0[15] );
tran (\sa_snapshot[9][15] , \sa_snapshot[9].f.lower[15] );
tran (\sa_snapshot[9][16] , \sa_snapshot[9].r.part0[16] );
tran (\sa_snapshot[9][16] , \sa_snapshot[9].f.lower[16] );
tran (\sa_snapshot[9][17] , \sa_snapshot[9].r.part0[17] );
tran (\sa_snapshot[9][17] , \sa_snapshot[9].f.lower[17] );
tran (\sa_snapshot[9][18] , \sa_snapshot[9].r.part0[18] );
tran (\sa_snapshot[9][18] , \sa_snapshot[9].f.lower[18] );
tran (\sa_snapshot[9][19] , \sa_snapshot[9].r.part0[19] );
tran (\sa_snapshot[9][19] , \sa_snapshot[9].f.lower[19] );
tran (\sa_snapshot[9][20] , \sa_snapshot[9].r.part0[20] );
tran (\sa_snapshot[9][20] , \sa_snapshot[9].f.lower[20] );
tran (\sa_snapshot[9][21] , \sa_snapshot[9].r.part0[21] );
tran (\sa_snapshot[9][21] , \sa_snapshot[9].f.lower[21] );
tran (\sa_snapshot[9][22] , \sa_snapshot[9].r.part0[22] );
tran (\sa_snapshot[9][22] , \sa_snapshot[9].f.lower[22] );
tran (\sa_snapshot[9][23] , \sa_snapshot[9].r.part0[23] );
tran (\sa_snapshot[9][23] , \sa_snapshot[9].f.lower[23] );
tran (\sa_snapshot[9][24] , \sa_snapshot[9].r.part0[24] );
tran (\sa_snapshot[9][24] , \sa_snapshot[9].f.lower[24] );
tran (\sa_snapshot[9][25] , \sa_snapshot[9].r.part0[25] );
tran (\sa_snapshot[9][25] , \sa_snapshot[9].f.lower[25] );
tran (\sa_snapshot[9][26] , \sa_snapshot[9].r.part0[26] );
tran (\sa_snapshot[9][26] , \sa_snapshot[9].f.lower[26] );
tran (\sa_snapshot[9][27] , \sa_snapshot[9].r.part0[27] );
tran (\sa_snapshot[9][27] , \sa_snapshot[9].f.lower[27] );
tran (\sa_snapshot[9][28] , \sa_snapshot[9].r.part0[28] );
tran (\sa_snapshot[9][28] , \sa_snapshot[9].f.lower[28] );
tran (\sa_snapshot[9][29] , \sa_snapshot[9].r.part0[29] );
tran (\sa_snapshot[9][29] , \sa_snapshot[9].f.lower[29] );
tran (\sa_snapshot[9][30] , \sa_snapshot[9].r.part0[30] );
tran (\sa_snapshot[9][30] , \sa_snapshot[9].f.lower[30] );
tran (\sa_snapshot[9][31] , \sa_snapshot[9].r.part0[31] );
tran (\sa_snapshot[9][31] , \sa_snapshot[9].f.lower[31] );
tran (\sa_snapshot[9][32] , \sa_snapshot[9].r.part1[0] );
tran (\sa_snapshot[9][32] , \sa_snapshot[9].f.upper[0] );
tran (\sa_snapshot[9][33] , \sa_snapshot[9].r.part1[1] );
tran (\sa_snapshot[9][33] , \sa_snapshot[9].f.upper[1] );
tran (\sa_snapshot[9][34] , \sa_snapshot[9].r.part1[2] );
tran (\sa_snapshot[9][34] , \sa_snapshot[9].f.upper[2] );
tran (\sa_snapshot[9][35] , \sa_snapshot[9].r.part1[3] );
tran (\sa_snapshot[9][35] , \sa_snapshot[9].f.upper[3] );
tran (\sa_snapshot[9][36] , \sa_snapshot[9].r.part1[4] );
tran (\sa_snapshot[9][36] , \sa_snapshot[9].f.upper[4] );
tran (\sa_snapshot[9][37] , \sa_snapshot[9].r.part1[5] );
tran (\sa_snapshot[9][37] , \sa_snapshot[9].f.upper[5] );
tran (\sa_snapshot[9][38] , \sa_snapshot[9].r.part1[6] );
tran (\sa_snapshot[9][38] , \sa_snapshot[9].f.upper[6] );
tran (\sa_snapshot[9][39] , \sa_snapshot[9].r.part1[7] );
tran (\sa_snapshot[9][39] , \sa_snapshot[9].f.upper[7] );
tran (\sa_snapshot[9][40] , \sa_snapshot[9].r.part1[8] );
tran (\sa_snapshot[9][40] , \sa_snapshot[9].f.upper[8] );
tran (\sa_snapshot[9][41] , \sa_snapshot[9].r.part1[9] );
tran (\sa_snapshot[9][41] , \sa_snapshot[9].f.upper[9] );
tran (\sa_snapshot[9][42] , \sa_snapshot[9].r.part1[10] );
tran (\sa_snapshot[9][42] , \sa_snapshot[9].f.upper[10] );
tran (\sa_snapshot[9][43] , \sa_snapshot[9].r.part1[11] );
tran (\sa_snapshot[9][43] , \sa_snapshot[9].f.upper[11] );
tran (\sa_snapshot[9][44] , \sa_snapshot[9].r.part1[12] );
tran (\sa_snapshot[9][44] , \sa_snapshot[9].f.upper[12] );
tran (\sa_snapshot[9][45] , \sa_snapshot[9].r.part1[13] );
tran (\sa_snapshot[9][45] , \sa_snapshot[9].f.upper[13] );
tran (\sa_snapshot[9][46] , \sa_snapshot[9].r.part1[14] );
tran (\sa_snapshot[9][46] , \sa_snapshot[9].f.upper[14] );
tran (\sa_snapshot[9][47] , \sa_snapshot[9].r.part1[15] );
tran (\sa_snapshot[9][47] , \sa_snapshot[9].f.upper[15] );
tran (\sa_snapshot[9][48] , \sa_snapshot[9].r.part1[16] );
tran (\sa_snapshot[9][48] , \sa_snapshot[9].f.upper[16] );
tran (\sa_snapshot[9][49] , \sa_snapshot[9].r.part1[17] );
tran (\sa_snapshot[9][49] , \sa_snapshot[9].f.upper[17] );
tran (\sa_snapshot[9][50] , \sa_snapshot[9].r.part1[18] );
tran (\sa_snapshot[9][50] , \sa_snapshot[9].f.unused[0] );
tran (\sa_snapshot[9][51] , \sa_snapshot[9].r.part1[19] );
tran (\sa_snapshot[9][51] , \sa_snapshot[9].f.unused[1] );
tran (\sa_snapshot[9][52] , \sa_snapshot[9].r.part1[20] );
tran (\sa_snapshot[9][52] , \sa_snapshot[9].f.unused[2] );
tran (\sa_snapshot[9][53] , \sa_snapshot[9].r.part1[21] );
tran (\sa_snapshot[9][53] , \sa_snapshot[9].f.unused[3] );
tran (\sa_snapshot[9][54] , \sa_snapshot[9].r.part1[22] );
tran (\sa_snapshot[9][54] , \sa_snapshot[9].f.unused[4] );
tran (\sa_snapshot[9][55] , \sa_snapshot[9].r.part1[23] );
tran (\sa_snapshot[9][55] , \sa_snapshot[9].f.unused[5] );
tran (\sa_snapshot[9][56] , \sa_snapshot[9].r.part1[24] );
tran (\sa_snapshot[9][56] , \sa_snapshot[9].f.unused[6] );
tran (\sa_snapshot[9][57] , \sa_snapshot[9].r.part1[25] );
tran (\sa_snapshot[9][57] , \sa_snapshot[9].f.unused[7] );
tran (\sa_snapshot[9][58] , \sa_snapshot[9].r.part1[26] );
tran (\sa_snapshot[9][58] , \sa_snapshot[9].f.unused[8] );
tran (\sa_snapshot[9][59] , \sa_snapshot[9].r.part1[27] );
tran (\sa_snapshot[9][59] , \sa_snapshot[9].f.unused[9] );
tran (\sa_snapshot[9][60] , \sa_snapshot[9].r.part1[28] );
tran (\sa_snapshot[9][60] , \sa_snapshot[9].f.unused[10] );
tran (\sa_snapshot[9][61] , \sa_snapshot[9].r.part1[29] );
tran (\sa_snapshot[9][61] , \sa_snapshot[9].f.unused[11] );
tran (\sa_snapshot[9][62] , \sa_snapshot[9].r.part1[30] );
tran (\sa_snapshot[9][62] , \sa_snapshot[9].f.unused[12] );
tran (\sa_snapshot[9][63] , \sa_snapshot[9].r.part1[31] );
tran (\sa_snapshot[9][63] , \sa_snapshot[9].f.unused[13] );
tran (\sa_snapshot[10][0] , \sa_snapshot[10].r.part0[0] );
tran (\sa_snapshot[10][0] , \sa_snapshot[10].f.lower[0] );
tran (\sa_snapshot[10][1] , \sa_snapshot[10].r.part0[1] );
tran (\sa_snapshot[10][1] , \sa_snapshot[10].f.lower[1] );
tran (\sa_snapshot[10][2] , \sa_snapshot[10].r.part0[2] );
tran (\sa_snapshot[10][2] , \sa_snapshot[10].f.lower[2] );
tran (\sa_snapshot[10][3] , \sa_snapshot[10].r.part0[3] );
tran (\sa_snapshot[10][3] , \sa_snapshot[10].f.lower[3] );
tran (\sa_snapshot[10][4] , \sa_snapshot[10].r.part0[4] );
tran (\sa_snapshot[10][4] , \sa_snapshot[10].f.lower[4] );
tran (\sa_snapshot[10][5] , \sa_snapshot[10].r.part0[5] );
tran (\sa_snapshot[10][5] , \sa_snapshot[10].f.lower[5] );
tran (\sa_snapshot[10][6] , \sa_snapshot[10].r.part0[6] );
tran (\sa_snapshot[10][6] , \sa_snapshot[10].f.lower[6] );
tran (\sa_snapshot[10][7] , \sa_snapshot[10].r.part0[7] );
tran (\sa_snapshot[10][7] , \sa_snapshot[10].f.lower[7] );
tran (\sa_snapshot[10][8] , \sa_snapshot[10].r.part0[8] );
tran (\sa_snapshot[10][8] , \sa_snapshot[10].f.lower[8] );
tran (\sa_snapshot[10][9] , \sa_snapshot[10].r.part0[9] );
tran (\sa_snapshot[10][9] , \sa_snapshot[10].f.lower[9] );
tran (\sa_snapshot[10][10] , \sa_snapshot[10].r.part0[10] );
tran (\sa_snapshot[10][10] , \sa_snapshot[10].f.lower[10] );
tran (\sa_snapshot[10][11] , \sa_snapshot[10].r.part0[11] );
tran (\sa_snapshot[10][11] , \sa_snapshot[10].f.lower[11] );
tran (\sa_snapshot[10][12] , \sa_snapshot[10].r.part0[12] );
tran (\sa_snapshot[10][12] , \sa_snapshot[10].f.lower[12] );
tran (\sa_snapshot[10][13] , \sa_snapshot[10].r.part0[13] );
tran (\sa_snapshot[10][13] , \sa_snapshot[10].f.lower[13] );
tran (\sa_snapshot[10][14] , \sa_snapshot[10].r.part0[14] );
tran (\sa_snapshot[10][14] , \sa_snapshot[10].f.lower[14] );
tran (\sa_snapshot[10][15] , \sa_snapshot[10].r.part0[15] );
tran (\sa_snapshot[10][15] , \sa_snapshot[10].f.lower[15] );
tran (\sa_snapshot[10][16] , \sa_snapshot[10].r.part0[16] );
tran (\sa_snapshot[10][16] , \sa_snapshot[10].f.lower[16] );
tran (\sa_snapshot[10][17] , \sa_snapshot[10].r.part0[17] );
tran (\sa_snapshot[10][17] , \sa_snapshot[10].f.lower[17] );
tran (\sa_snapshot[10][18] , \sa_snapshot[10].r.part0[18] );
tran (\sa_snapshot[10][18] , \sa_snapshot[10].f.lower[18] );
tran (\sa_snapshot[10][19] , \sa_snapshot[10].r.part0[19] );
tran (\sa_snapshot[10][19] , \sa_snapshot[10].f.lower[19] );
tran (\sa_snapshot[10][20] , \sa_snapshot[10].r.part0[20] );
tran (\sa_snapshot[10][20] , \sa_snapshot[10].f.lower[20] );
tran (\sa_snapshot[10][21] , \sa_snapshot[10].r.part0[21] );
tran (\sa_snapshot[10][21] , \sa_snapshot[10].f.lower[21] );
tran (\sa_snapshot[10][22] , \sa_snapshot[10].r.part0[22] );
tran (\sa_snapshot[10][22] , \sa_snapshot[10].f.lower[22] );
tran (\sa_snapshot[10][23] , \sa_snapshot[10].r.part0[23] );
tran (\sa_snapshot[10][23] , \sa_snapshot[10].f.lower[23] );
tran (\sa_snapshot[10][24] , \sa_snapshot[10].r.part0[24] );
tran (\sa_snapshot[10][24] , \sa_snapshot[10].f.lower[24] );
tran (\sa_snapshot[10][25] , \sa_snapshot[10].r.part0[25] );
tran (\sa_snapshot[10][25] , \sa_snapshot[10].f.lower[25] );
tran (\sa_snapshot[10][26] , \sa_snapshot[10].r.part0[26] );
tran (\sa_snapshot[10][26] , \sa_snapshot[10].f.lower[26] );
tran (\sa_snapshot[10][27] , \sa_snapshot[10].r.part0[27] );
tran (\sa_snapshot[10][27] , \sa_snapshot[10].f.lower[27] );
tran (\sa_snapshot[10][28] , \sa_snapshot[10].r.part0[28] );
tran (\sa_snapshot[10][28] , \sa_snapshot[10].f.lower[28] );
tran (\sa_snapshot[10][29] , \sa_snapshot[10].r.part0[29] );
tran (\sa_snapshot[10][29] , \sa_snapshot[10].f.lower[29] );
tran (\sa_snapshot[10][30] , \sa_snapshot[10].r.part0[30] );
tran (\sa_snapshot[10][30] , \sa_snapshot[10].f.lower[30] );
tran (\sa_snapshot[10][31] , \sa_snapshot[10].r.part0[31] );
tran (\sa_snapshot[10][31] , \sa_snapshot[10].f.lower[31] );
tran (\sa_snapshot[10][32] , \sa_snapshot[10].r.part1[0] );
tran (\sa_snapshot[10][32] , \sa_snapshot[10].f.upper[0] );
tran (\sa_snapshot[10][33] , \sa_snapshot[10].r.part1[1] );
tran (\sa_snapshot[10][33] , \sa_snapshot[10].f.upper[1] );
tran (\sa_snapshot[10][34] , \sa_snapshot[10].r.part1[2] );
tran (\sa_snapshot[10][34] , \sa_snapshot[10].f.upper[2] );
tran (\sa_snapshot[10][35] , \sa_snapshot[10].r.part1[3] );
tran (\sa_snapshot[10][35] , \sa_snapshot[10].f.upper[3] );
tran (\sa_snapshot[10][36] , \sa_snapshot[10].r.part1[4] );
tran (\sa_snapshot[10][36] , \sa_snapshot[10].f.upper[4] );
tran (\sa_snapshot[10][37] , \sa_snapshot[10].r.part1[5] );
tran (\sa_snapshot[10][37] , \sa_snapshot[10].f.upper[5] );
tran (\sa_snapshot[10][38] , \sa_snapshot[10].r.part1[6] );
tran (\sa_snapshot[10][38] , \sa_snapshot[10].f.upper[6] );
tran (\sa_snapshot[10][39] , \sa_snapshot[10].r.part1[7] );
tran (\sa_snapshot[10][39] , \sa_snapshot[10].f.upper[7] );
tran (\sa_snapshot[10][40] , \sa_snapshot[10].r.part1[8] );
tran (\sa_snapshot[10][40] , \sa_snapshot[10].f.upper[8] );
tran (\sa_snapshot[10][41] , \sa_snapshot[10].r.part1[9] );
tran (\sa_snapshot[10][41] , \sa_snapshot[10].f.upper[9] );
tran (\sa_snapshot[10][42] , \sa_snapshot[10].r.part1[10] );
tran (\sa_snapshot[10][42] , \sa_snapshot[10].f.upper[10] );
tran (\sa_snapshot[10][43] , \sa_snapshot[10].r.part1[11] );
tran (\sa_snapshot[10][43] , \sa_snapshot[10].f.upper[11] );
tran (\sa_snapshot[10][44] , \sa_snapshot[10].r.part1[12] );
tran (\sa_snapshot[10][44] , \sa_snapshot[10].f.upper[12] );
tran (\sa_snapshot[10][45] , \sa_snapshot[10].r.part1[13] );
tran (\sa_snapshot[10][45] , \sa_snapshot[10].f.upper[13] );
tran (\sa_snapshot[10][46] , \sa_snapshot[10].r.part1[14] );
tran (\sa_snapshot[10][46] , \sa_snapshot[10].f.upper[14] );
tran (\sa_snapshot[10][47] , \sa_snapshot[10].r.part1[15] );
tran (\sa_snapshot[10][47] , \sa_snapshot[10].f.upper[15] );
tran (\sa_snapshot[10][48] , \sa_snapshot[10].r.part1[16] );
tran (\sa_snapshot[10][48] , \sa_snapshot[10].f.upper[16] );
tran (\sa_snapshot[10][49] , \sa_snapshot[10].r.part1[17] );
tran (\sa_snapshot[10][49] , \sa_snapshot[10].f.upper[17] );
tran (\sa_snapshot[10][50] , \sa_snapshot[10].r.part1[18] );
tran (\sa_snapshot[10][50] , \sa_snapshot[10].f.unused[0] );
tran (\sa_snapshot[10][51] , \sa_snapshot[10].r.part1[19] );
tran (\sa_snapshot[10][51] , \sa_snapshot[10].f.unused[1] );
tran (\sa_snapshot[10][52] , \sa_snapshot[10].r.part1[20] );
tran (\sa_snapshot[10][52] , \sa_snapshot[10].f.unused[2] );
tran (\sa_snapshot[10][53] , \sa_snapshot[10].r.part1[21] );
tran (\sa_snapshot[10][53] , \sa_snapshot[10].f.unused[3] );
tran (\sa_snapshot[10][54] , \sa_snapshot[10].r.part1[22] );
tran (\sa_snapshot[10][54] , \sa_snapshot[10].f.unused[4] );
tran (\sa_snapshot[10][55] , \sa_snapshot[10].r.part1[23] );
tran (\sa_snapshot[10][55] , \sa_snapshot[10].f.unused[5] );
tran (\sa_snapshot[10][56] , \sa_snapshot[10].r.part1[24] );
tran (\sa_snapshot[10][56] , \sa_snapshot[10].f.unused[6] );
tran (\sa_snapshot[10][57] , \sa_snapshot[10].r.part1[25] );
tran (\sa_snapshot[10][57] , \sa_snapshot[10].f.unused[7] );
tran (\sa_snapshot[10][58] , \sa_snapshot[10].r.part1[26] );
tran (\sa_snapshot[10][58] , \sa_snapshot[10].f.unused[8] );
tran (\sa_snapshot[10][59] , \sa_snapshot[10].r.part1[27] );
tran (\sa_snapshot[10][59] , \sa_snapshot[10].f.unused[9] );
tran (\sa_snapshot[10][60] , \sa_snapshot[10].r.part1[28] );
tran (\sa_snapshot[10][60] , \sa_snapshot[10].f.unused[10] );
tran (\sa_snapshot[10][61] , \sa_snapshot[10].r.part1[29] );
tran (\sa_snapshot[10][61] , \sa_snapshot[10].f.unused[11] );
tran (\sa_snapshot[10][62] , \sa_snapshot[10].r.part1[30] );
tran (\sa_snapshot[10][62] , \sa_snapshot[10].f.unused[12] );
tran (\sa_snapshot[10][63] , \sa_snapshot[10].r.part1[31] );
tran (\sa_snapshot[10][63] , \sa_snapshot[10].f.unused[13] );
tran (\sa_snapshot[11][0] , \sa_snapshot[11].r.part0[0] );
tran (\sa_snapshot[11][0] , \sa_snapshot[11].f.lower[0] );
tran (\sa_snapshot[11][1] , \sa_snapshot[11].r.part0[1] );
tran (\sa_snapshot[11][1] , \sa_snapshot[11].f.lower[1] );
tran (\sa_snapshot[11][2] , \sa_snapshot[11].r.part0[2] );
tran (\sa_snapshot[11][2] , \sa_snapshot[11].f.lower[2] );
tran (\sa_snapshot[11][3] , \sa_snapshot[11].r.part0[3] );
tran (\sa_snapshot[11][3] , \sa_snapshot[11].f.lower[3] );
tran (\sa_snapshot[11][4] , \sa_snapshot[11].r.part0[4] );
tran (\sa_snapshot[11][4] , \sa_snapshot[11].f.lower[4] );
tran (\sa_snapshot[11][5] , \sa_snapshot[11].r.part0[5] );
tran (\sa_snapshot[11][5] , \sa_snapshot[11].f.lower[5] );
tran (\sa_snapshot[11][6] , \sa_snapshot[11].r.part0[6] );
tran (\sa_snapshot[11][6] , \sa_snapshot[11].f.lower[6] );
tran (\sa_snapshot[11][7] , \sa_snapshot[11].r.part0[7] );
tran (\sa_snapshot[11][7] , \sa_snapshot[11].f.lower[7] );
tran (\sa_snapshot[11][8] , \sa_snapshot[11].r.part0[8] );
tran (\sa_snapshot[11][8] , \sa_snapshot[11].f.lower[8] );
tran (\sa_snapshot[11][9] , \sa_snapshot[11].r.part0[9] );
tran (\sa_snapshot[11][9] , \sa_snapshot[11].f.lower[9] );
tran (\sa_snapshot[11][10] , \sa_snapshot[11].r.part0[10] );
tran (\sa_snapshot[11][10] , \sa_snapshot[11].f.lower[10] );
tran (\sa_snapshot[11][11] , \sa_snapshot[11].r.part0[11] );
tran (\sa_snapshot[11][11] , \sa_snapshot[11].f.lower[11] );
tran (\sa_snapshot[11][12] , \sa_snapshot[11].r.part0[12] );
tran (\sa_snapshot[11][12] , \sa_snapshot[11].f.lower[12] );
tran (\sa_snapshot[11][13] , \sa_snapshot[11].r.part0[13] );
tran (\sa_snapshot[11][13] , \sa_snapshot[11].f.lower[13] );
tran (\sa_snapshot[11][14] , \sa_snapshot[11].r.part0[14] );
tran (\sa_snapshot[11][14] , \sa_snapshot[11].f.lower[14] );
tran (\sa_snapshot[11][15] , \sa_snapshot[11].r.part0[15] );
tran (\sa_snapshot[11][15] , \sa_snapshot[11].f.lower[15] );
tran (\sa_snapshot[11][16] , \sa_snapshot[11].r.part0[16] );
tran (\sa_snapshot[11][16] , \sa_snapshot[11].f.lower[16] );
tran (\sa_snapshot[11][17] , \sa_snapshot[11].r.part0[17] );
tran (\sa_snapshot[11][17] , \sa_snapshot[11].f.lower[17] );
tran (\sa_snapshot[11][18] , \sa_snapshot[11].r.part0[18] );
tran (\sa_snapshot[11][18] , \sa_snapshot[11].f.lower[18] );
tran (\sa_snapshot[11][19] , \sa_snapshot[11].r.part0[19] );
tran (\sa_snapshot[11][19] , \sa_snapshot[11].f.lower[19] );
tran (\sa_snapshot[11][20] , \sa_snapshot[11].r.part0[20] );
tran (\sa_snapshot[11][20] , \sa_snapshot[11].f.lower[20] );
tran (\sa_snapshot[11][21] , \sa_snapshot[11].r.part0[21] );
tran (\sa_snapshot[11][21] , \sa_snapshot[11].f.lower[21] );
tran (\sa_snapshot[11][22] , \sa_snapshot[11].r.part0[22] );
tran (\sa_snapshot[11][22] , \sa_snapshot[11].f.lower[22] );
tran (\sa_snapshot[11][23] , \sa_snapshot[11].r.part0[23] );
tran (\sa_snapshot[11][23] , \sa_snapshot[11].f.lower[23] );
tran (\sa_snapshot[11][24] , \sa_snapshot[11].r.part0[24] );
tran (\sa_snapshot[11][24] , \sa_snapshot[11].f.lower[24] );
tran (\sa_snapshot[11][25] , \sa_snapshot[11].r.part0[25] );
tran (\sa_snapshot[11][25] , \sa_snapshot[11].f.lower[25] );
tran (\sa_snapshot[11][26] , \sa_snapshot[11].r.part0[26] );
tran (\sa_snapshot[11][26] , \sa_snapshot[11].f.lower[26] );
tran (\sa_snapshot[11][27] , \sa_snapshot[11].r.part0[27] );
tran (\sa_snapshot[11][27] , \sa_snapshot[11].f.lower[27] );
tran (\sa_snapshot[11][28] , \sa_snapshot[11].r.part0[28] );
tran (\sa_snapshot[11][28] , \sa_snapshot[11].f.lower[28] );
tran (\sa_snapshot[11][29] , \sa_snapshot[11].r.part0[29] );
tran (\sa_snapshot[11][29] , \sa_snapshot[11].f.lower[29] );
tran (\sa_snapshot[11][30] , \sa_snapshot[11].r.part0[30] );
tran (\sa_snapshot[11][30] , \sa_snapshot[11].f.lower[30] );
tran (\sa_snapshot[11][31] , \sa_snapshot[11].r.part0[31] );
tran (\sa_snapshot[11][31] , \sa_snapshot[11].f.lower[31] );
tran (\sa_snapshot[11][32] , \sa_snapshot[11].r.part1[0] );
tran (\sa_snapshot[11][32] , \sa_snapshot[11].f.upper[0] );
tran (\sa_snapshot[11][33] , \sa_snapshot[11].r.part1[1] );
tran (\sa_snapshot[11][33] , \sa_snapshot[11].f.upper[1] );
tran (\sa_snapshot[11][34] , \sa_snapshot[11].r.part1[2] );
tran (\sa_snapshot[11][34] , \sa_snapshot[11].f.upper[2] );
tran (\sa_snapshot[11][35] , \sa_snapshot[11].r.part1[3] );
tran (\sa_snapshot[11][35] , \sa_snapshot[11].f.upper[3] );
tran (\sa_snapshot[11][36] , \sa_snapshot[11].r.part1[4] );
tran (\sa_snapshot[11][36] , \sa_snapshot[11].f.upper[4] );
tran (\sa_snapshot[11][37] , \sa_snapshot[11].r.part1[5] );
tran (\sa_snapshot[11][37] , \sa_snapshot[11].f.upper[5] );
tran (\sa_snapshot[11][38] , \sa_snapshot[11].r.part1[6] );
tran (\sa_snapshot[11][38] , \sa_snapshot[11].f.upper[6] );
tran (\sa_snapshot[11][39] , \sa_snapshot[11].r.part1[7] );
tran (\sa_snapshot[11][39] , \sa_snapshot[11].f.upper[7] );
tran (\sa_snapshot[11][40] , \sa_snapshot[11].r.part1[8] );
tran (\sa_snapshot[11][40] , \sa_snapshot[11].f.upper[8] );
tran (\sa_snapshot[11][41] , \sa_snapshot[11].r.part1[9] );
tran (\sa_snapshot[11][41] , \sa_snapshot[11].f.upper[9] );
tran (\sa_snapshot[11][42] , \sa_snapshot[11].r.part1[10] );
tran (\sa_snapshot[11][42] , \sa_snapshot[11].f.upper[10] );
tran (\sa_snapshot[11][43] , \sa_snapshot[11].r.part1[11] );
tran (\sa_snapshot[11][43] , \sa_snapshot[11].f.upper[11] );
tran (\sa_snapshot[11][44] , \sa_snapshot[11].r.part1[12] );
tran (\sa_snapshot[11][44] , \sa_snapshot[11].f.upper[12] );
tran (\sa_snapshot[11][45] , \sa_snapshot[11].r.part1[13] );
tran (\sa_snapshot[11][45] , \sa_snapshot[11].f.upper[13] );
tran (\sa_snapshot[11][46] , \sa_snapshot[11].r.part1[14] );
tran (\sa_snapshot[11][46] , \sa_snapshot[11].f.upper[14] );
tran (\sa_snapshot[11][47] , \sa_snapshot[11].r.part1[15] );
tran (\sa_snapshot[11][47] , \sa_snapshot[11].f.upper[15] );
tran (\sa_snapshot[11][48] , \sa_snapshot[11].r.part1[16] );
tran (\sa_snapshot[11][48] , \sa_snapshot[11].f.upper[16] );
tran (\sa_snapshot[11][49] , \sa_snapshot[11].r.part1[17] );
tran (\sa_snapshot[11][49] , \sa_snapshot[11].f.upper[17] );
tran (\sa_snapshot[11][50] , \sa_snapshot[11].r.part1[18] );
tran (\sa_snapshot[11][50] , \sa_snapshot[11].f.unused[0] );
tran (\sa_snapshot[11][51] , \sa_snapshot[11].r.part1[19] );
tran (\sa_snapshot[11][51] , \sa_snapshot[11].f.unused[1] );
tran (\sa_snapshot[11][52] , \sa_snapshot[11].r.part1[20] );
tran (\sa_snapshot[11][52] , \sa_snapshot[11].f.unused[2] );
tran (\sa_snapshot[11][53] , \sa_snapshot[11].r.part1[21] );
tran (\sa_snapshot[11][53] , \sa_snapshot[11].f.unused[3] );
tran (\sa_snapshot[11][54] , \sa_snapshot[11].r.part1[22] );
tran (\sa_snapshot[11][54] , \sa_snapshot[11].f.unused[4] );
tran (\sa_snapshot[11][55] , \sa_snapshot[11].r.part1[23] );
tran (\sa_snapshot[11][55] , \sa_snapshot[11].f.unused[5] );
tran (\sa_snapshot[11][56] , \sa_snapshot[11].r.part1[24] );
tran (\sa_snapshot[11][56] , \sa_snapshot[11].f.unused[6] );
tran (\sa_snapshot[11][57] , \sa_snapshot[11].r.part1[25] );
tran (\sa_snapshot[11][57] , \sa_snapshot[11].f.unused[7] );
tran (\sa_snapshot[11][58] , \sa_snapshot[11].r.part1[26] );
tran (\sa_snapshot[11][58] , \sa_snapshot[11].f.unused[8] );
tran (\sa_snapshot[11][59] , \sa_snapshot[11].r.part1[27] );
tran (\sa_snapshot[11][59] , \sa_snapshot[11].f.unused[9] );
tran (\sa_snapshot[11][60] , \sa_snapshot[11].r.part1[28] );
tran (\sa_snapshot[11][60] , \sa_snapshot[11].f.unused[10] );
tran (\sa_snapshot[11][61] , \sa_snapshot[11].r.part1[29] );
tran (\sa_snapshot[11][61] , \sa_snapshot[11].f.unused[11] );
tran (\sa_snapshot[11][62] , \sa_snapshot[11].r.part1[30] );
tran (\sa_snapshot[11][62] , \sa_snapshot[11].f.unused[12] );
tran (\sa_snapshot[11][63] , \sa_snapshot[11].r.part1[31] );
tran (\sa_snapshot[11][63] , \sa_snapshot[11].f.unused[13] );
tran (\sa_snapshot[12][0] , \sa_snapshot[12].r.part0[0] );
tran (\sa_snapshot[12][0] , \sa_snapshot[12].f.lower[0] );
tran (\sa_snapshot[12][1] , \sa_snapshot[12].r.part0[1] );
tran (\sa_snapshot[12][1] , \sa_snapshot[12].f.lower[1] );
tran (\sa_snapshot[12][2] , \sa_snapshot[12].r.part0[2] );
tran (\sa_snapshot[12][2] , \sa_snapshot[12].f.lower[2] );
tran (\sa_snapshot[12][3] , \sa_snapshot[12].r.part0[3] );
tran (\sa_snapshot[12][3] , \sa_snapshot[12].f.lower[3] );
tran (\sa_snapshot[12][4] , \sa_snapshot[12].r.part0[4] );
tran (\sa_snapshot[12][4] , \sa_snapshot[12].f.lower[4] );
tran (\sa_snapshot[12][5] , \sa_snapshot[12].r.part0[5] );
tran (\sa_snapshot[12][5] , \sa_snapshot[12].f.lower[5] );
tran (\sa_snapshot[12][6] , \sa_snapshot[12].r.part0[6] );
tran (\sa_snapshot[12][6] , \sa_snapshot[12].f.lower[6] );
tran (\sa_snapshot[12][7] , \sa_snapshot[12].r.part0[7] );
tran (\sa_snapshot[12][7] , \sa_snapshot[12].f.lower[7] );
tran (\sa_snapshot[12][8] , \sa_snapshot[12].r.part0[8] );
tran (\sa_snapshot[12][8] , \sa_snapshot[12].f.lower[8] );
tran (\sa_snapshot[12][9] , \sa_snapshot[12].r.part0[9] );
tran (\sa_snapshot[12][9] , \sa_snapshot[12].f.lower[9] );
tran (\sa_snapshot[12][10] , \sa_snapshot[12].r.part0[10] );
tran (\sa_snapshot[12][10] , \sa_snapshot[12].f.lower[10] );
tran (\sa_snapshot[12][11] , \sa_snapshot[12].r.part0[11] );
tran (\sa_snapshot[12][11] , \sa_snapshot[12].f.lower[11] );
tran (\sa_snapshot[12][12] , \sa_snapshot[12].r.part0[12] );
tran (\sa_snapshot[12][12] , \sa_snapshot[12].f.lower[12] );
tran (\sa_snapshot[12][13] , \sa_snapshot[12].r.part0[13] );
tran (\sa_snapshot[12][13] , \sa_snapshot[12].f.lower[13] );
tran (\sa_snapshot[12][14] , \sa_snapshot[12].r.part0[14] );
tran (\sa_snapshot[12][14] , \sa_snapshot[12].f.lower[14] );
tran (\sa_snapshot[12][15] , \sa_snapshot[12].r.part0[15] );
tran (\sa_snapshot[12][15] , \sa_snapshot[12].f.lower[15] );
tran (\sa_snapshot[12][16] , \sa_snapshot[12].r.part0[16] );
tran (\sa_snapshot[12][16] , \sa_snapshot[12].f.lower[16] );
tran (\sa_snapshot[12][17] , \sa_snapshot[12].r.part0[17] );
tran (\sa_snapshot[12][17] , \sa_snapshot[12].f.lower[17] );
tran (\sa_snapshot[12][18] , \sa_snapshot[12].r.part0[18] );
tran (\sa_snapshot[12][18] , \sa_snapshot[12].f.lower[18] );
tran (\sa_snapshot[12][19] , \sa_snapshot[12].r.part0[19] );
tran (\sa_snapshot[12][19] , \sa_snapshot[12].f.lower[19] );
tran (\sa_snapshot[12][20] , \sa_snapshot[12].r.part0[20] );
tran (\sa_snapshot[12][20] , \sa_snapshot[12].f.lower[20] );
tran (\sa_snapshot[12][21] , \sa_snapshot[12].r.part0[21] );
tran (\sa_snapshot[12][21] , \sa_snapshot[12].f.lower[21] );
tran (\sa_snapshot[12][22] , \sa_snapshot[12].r.part0[22] );
tran (\sa_snapshot[12][22] , \sa_snapshot[12].f.lower[22] );
tran (\sa_snapshot[12][23] , \sa_snapshot[12].r.part0[23] );
tran (\sa_snapshot[12][23] , \sa_snapshot[12].f.lower[23] );
tran (\sa_snapshot[12][24] , \sa_snapshot[12].r.part0[24] );
tran (\sa_snapshot[12][24] , \sa_snapshot[12].f.lower[24] );
tran (\sa_snapshot[12][25] , \sa_snapshot[12].r.part0[25] );
tran (\sa_snapshot[12][25] , \sa_snapshot[12].f.lower[25] );
tran (\sa_snapshot[12][26] , \sa_snapshot[12].r.part0[26] );
tran (\sa_snapshot[12][26] , \sa_snapshot[12].f.lower[26] );
tran (\sa_snapshot[12][27] , \sa_snapshot[12].r.part0[27] );
tran (\sa_snapshot[12][27] , \sa_snapshot[12].f.lower[27] );
tran (\sa_snapshot[12][28] , \sa_snapshot[12].r.part0[28] );
tran (\sa_snapshot[12][28] , \sa_snapshot[12].f.lower[28] );
tran (\sa_snapshot[12][29] , \sa_snapshot[12].r.part0[29] );
tran (\sa_snapshot[12][29] , \sa_snapshot[12].f.lower[29] );
tran (\sa_snapshot[12][30] , \sa_snapshot[12].r.part0[30] );
tran (\sa_snapshot[12][30] , \sa_snapshot[12].f.lower[30] );
tran (\sa_snapshot[12][31] , \sa_snapshot[12].r.part0[31] );
tran (\sa_snapshot[12][31] , \sa_snapshot[12].f.lower[31] );
tran (\sa_snapshot[12][32] , \sa_snapshot[12].r.part1[0] );
tran (\sa_snapshot[12][32] , \sa_snapshot[12].f.upper[0] );
tran (\sa_snapshot[12][33] , \sa_snapshot[12].r.part1[1] );
tran (\sa_snapshot[12][33] , \sa_snapshot[12].f.upper[1] );
tran (\sa_snapshot[12][34] , \sa_snapshot[12].r.part1[2] );
tran (\sa_snapshot[12][34] , \sa_snapshot[12].f.upper[2] );
tran (\sa_snapshot[12][35] , \sa_snapshot[12].r.part1[3] );
tran (\sa_snapshot[12][35] , \sa_snapshot[12].f.upper[3] );
tran (\sa_snapshot[12][36] , \sa_snapshot[12].r.part1[4] );
tran (\sa_snapshot[12][36] , \sa_snapshot[12].f.upper[4] );
tran (\sa_snapshot[12][37] , \sa_snapshot[12].r.part1[5] );
tran (\sa_snapshot[12][37] , \sa_snapshot[12].f.upper[5] );
tran (\sa_snapshot[12][38] , \sa_snapshot[12].r.part1[6] );
tran (\sa_snapshot[12][38] , \sa_snapshot[12].f.upper[6] );
tran (\sa_snapshot[12][39] , \sa_snapshot[12].r.part1[7] );
tran (\sa_snapshot[12][39] , \sa_snapshot[12].f.upper[7] );
tran (\sa_snapshot[12][40] , \sa_snapshot[12].r.part1[8] );
tran (\sa_snapshot[12][40] , \sa_snapshot[12].f.upper[8] );
tran (\sa_snapshot[12][41] , \sa_snapshot[12].r.part1[9] );
tran (\sa_snapshot[12][41] , \sa_snapshot[12].f.upper[9] );
tran (\sa_snapshot[12][42] , \sa_snapshot[12].r.part1[10] );
tran (\sa_snapshot[12][42] , \sa_snapshot[12].f.upper[10] );
tran (\sa_snapshot[12][43] , \sa_snapshot[12].r.part1[11] );
tran (\sa_snapshot[12][43] , \sa_snapshot[12].f.upper[11] );
tran (\sa_snapshot[12][44] , \sa_snapshot[12].r.part1[12] );
tran (\sa_snapshot[12][44] , \sa_snapshot[12].f.upper[12] );
tran (\sa_snapshot[12][45] , \sa_snapshot[12].r.part1[13] );
tran (\sa_snapshot[12][45] , \sa_snapshot[12].f.upper[13] );
tran (\sa_snapshot[12][46] , \sa_snapshot[12].r.part1[14] );
tran (\sa_snapshot[12][46] , \sa_snapshot[12].f.upper[14] );
tran (\sa_snapshot[12][47] , \sa_snapshot[12].r.part1[15] );
tran (\sa_snapshot[12][47] , \sa_snapshot[12].f.upper[15] );
tran (\sa_snapshot[12][48] , \sa_snapshot[12].r.part1[16] );
tran (\sa_snapshot[12][48] , \sa_snapshot[12].f.upper[16] );
tran (\sa_snapshot[12][49] , \sa_snapshot[12].r.part1[17] );
tran (\sa_snapshot[12][49] , \sa_snapshot[12].f.upper[17] );
tran (\sa_snapshot[12][50] , \sa_snapshot[12].r.part1[18] );
tran (\sa_snapshot[12][50] , \sa_snapshot[12].f.unused[0] );
tran (\sa_snapshot[12][51] , \sa_snapshot[12].r.part1[19] );
tran (\sa_snapshot[12][51] , \sa_snapshot[12].f.unused[1] );
tran (\sa_snapshot[12][52] , \sa_snapshot[12].r.part1[20] );
tran (\sa_snapshot[12][52] , \sa_snapshot[12].f.unused[2] );
tran (\sa_snapshot[12][53] , \sa_snapshot[12].r.part1[21] );
tran (\sa_snapshot[12][53] , \sa_snapshot[12].f.unused[3] );
tran (\sa_snapshot[12][54] , \sa_snapshot[12].r.part1[22] );
tran (\sa_snapshot[12][54] , \sa_snapshot[12].f.unused[4] );
tran (\sa_snapshot[12][55] , \sa_snapshot[12].r.part1[23] );
tran (\sa_snapshot[12][55] , \sa_snapshot[12].f.unused[5] );
tran (\sa_snapshot[12][56] , \sa_snapshot[12].r.part1[24] );
tran (\sa_snapshot[12][56] , \sa_snapshot[12].f.unused[6] );
tran (\sa_snapshot[12][57] , \sa_snapshot[12].r.part1[25] );
tran (\sa_snapshot[12][57] , \sa_snapshot[12].f.unused[7] );
tran (\sa_snapshot[12][58] , \sa_snapshot[12].r.part1[26] );
tran (\sa_snapshot[12][58] , \sa_snapshot[12].f.unused[8] );
tran (\sa_snapshot[12][59] , \sa_snapshot[12].r.part1[27] );
tran (\sa_snapshot[12][59] , \sa_snapshot[12].f.unused[9] );
tran (\sa_snapshot[12][60] , \sa_snapshot[12].r.part1[28] );
tran (\sa_snapshot[12][60] , \sa_snapshot[12].f.unused[10] );
tran (\sa_snapshot[12][61] , \sa_snapshot[12].r.part1[29] );
tran (\sa_snapshot[12][61] , \sa_snapshot[12].f.unused[11] );
tran (\sa_snapshot[12][62] , \sa_snapshot[12].r.part1[30] );
tran (\sa_snapshot[12][62] , \sa_snapshot[12].f.unused[12] );
tran (\sa_snapshot[12][63] , \sa_snapshot[12].r.part1[31] );
tran (\sa_snapshot[12][63] , \sa_snapshot[12].f.unused[13] );
tran (\sa_snapshot[13][0] , \sa_snapshot[13].r.part0[0] );
tran (\sa_snapshot[13][0] , \sa_snapshot[13].f.lower[0] );
tran (\sa_snapshot[13][1] , \sa_snapshot[13].r.part0[1] );
tran (\sa_snapshot[13][1] , \sa_snapshot[13].f.lower[1] );
tran (\sa_snapshot[13][2] , \sa_snapshot[13].r.part0[2] );
tran (\sa_snapshot[13][2] , \sa_snapshot[13].f.lower[2] );
tran (\sa_snapshot[13][3] , \sa_snapshot[13].r.part0[3] );
tran (\sa_snapshot[13][3] , \sa_snapshot[13].f.lower[3] );
tran (\sa_snapshot[13][4] , \sa_snapshot[13].r.part0[4] );
tran (\sa_snapshot[13][4] , \sa_snapshot[13].f.lower[4] );
tran (\sa_snapshot[13][5] , \sa_snapshot[13].r.part0[5] );
tran (\sa_snapshot[13][5] , \sa_snapshot[13].f.lower[5] );
tran (\sa_snapshot[13][6] , \sa_snapshot[13].r.part0[6] );
tran (\sa_snapshot[13][6] , \sa_snapshot[13].f.lower[6] );
tran (\sa_snapshot[13][7] , \sa_snapshot[13].r.part0[7] );
tran (\sa_snapshot[13][7] , \sa_snapshot[13].f.lower[7] );
tran (\sa_snapshot[13][8] , \sa_snapshot[13].r.part0[8] );
tran (\sa_snapshot[13][8] , \sa_snapshot[13].f.lower[8] );
tran (\sa_snapshot[13][9] , \sa_snapshot[13].r.part0[9] );
tran (\sa_snapshot[13][9] , \sa_snapshot[13].f.lower[9] );
tran (\sa_snapshot[13][10] , \sa_snapshot[13].r.part0[10] );
tran (\sa_snapshot[13][10] , \sa_snapshot[13].f.lower[10] );
tran (\sa_snapshot[13][11] , \sa_snapshot[13].r.part0[11] );
tran (\sa_snapshot[13][11] , \sa_snapshot[13].f.lower[11] );
tran (\sa_snapshot[13][12] , \sa_snapshot[13].r.part0[12] );
tran (\sa_snapshot[13][12] , \sa_snapshot[13].f.lower[12] );
tran (\sa_snapshot[13][13] , \sa_snapshot[13].r.part0[13] );
tran (\sa_snapshot[13][13] , \sa_snapshot[13].f.lower[13] );
tran (\sa_snapshot[13][14] , \sa_snapshot[13].r.part0[14] );
tran (\sa_snapshot[13][14] , \sa_snapshot[13].f.lower[14] );
tran (\sa_snapshot[13][15] , \sa_snapshot[13].r.part0[15] );
tran (\sa_snapshot[13][15] , \sa_snapshot[13].f.lower[15] );
tran (\sa_snapshot[13][16] , \sa_snapshot[13].r.part0[16] );
tran (\sa_snapshot[13][16] , \sa_snapshot[13].f.lower[16] );
tran (\sa_snapshot[13][17] , \sa_snapshot[13].r.part0[17] );
tran (\sa_snapshot[13][17] , \sa_snapshot[13].f.lower[17] );
tran (\sa_snapshot[13][18] , \sa_snapshot[13].r.part0[18] );
tran (\sa_snapshot[13][18] , \sa_snapshot[13].f.lower[18] );
tran (\sa_snapshot[13][19] , \sa_snapshot[13].r.part0[19] );
tran (\sa_snapshot[13][19] , \sa_snapshot[13].f.lower[19] );
tran (\sa_snapshot[13][20] , \sa_snapshot[13].r.part0[20] );
tran (\sa_snapshot[13][20] , \sa_snapshot[13].f.lower[20] );
tran (\sa_snapshot[13][21] , \sa_snapshot[13].r.part0[21] );
tran (\sa_snapshot[13][21] , \sa_snapshot[13].f.lower[21] );
tran (\sa_snapshot[13][22] , \sa_snapshot[13].r.part0[22] );
tran (\sa_snapshot[13][22] , \sa_snapshot[13].f.lower[22] );
tran (\sa_snapshot[13][23] , \sa_snapshot[13].r.part0[23] );
tran (\sa_snapshot[13][23] , \sa_snapshot[13].f.lower[23] );
tran (\sa_snapshot[13][24] , \sa_snapshot[13].r.part0[24] );
tran (\sa_snapshot[13][24] , \sa_snapshot[13].f.lower[24] );
tran (\sa_snapshot[13][25] , \sa_snapshot[13].r.part0[25] );
tran (\sa_snapshot[13][25] , \sa_snapshot[13].f.lower[25] );
tran (\sa_snapshot[13][26] , \sa_snapshot[13].r.part0[26] );
tran (\sa_snapshot[13][26] , \sa_snapshot[13].f.lower[26] );
tran (\sa_snapshot[13][27] , \sa_snapshot[13].r.part0[27] );
tran (\sa_snapshot[13][27] , \sa_snapshot[13].f.lower[27] );
tran (\sa_snapshot[13][28] , \sa_snapshot[13].r.part0[28] );
tran (\sa_snapshot[13][28] , \sa_snapshot[13].f.lower[28] );
tran (\sa_snapshot[13][29] , \sa_snapshot[13].r.part0[29] );
tran (\sa_snapshot[13][29] , \sa_snapshot[13].f.lower[29] );
tran (\sa_snapshot[13][30] , \sa_snapshot[13].r.part0[30] );
tran (\sa_snapshot[13][30] , \sa_snapshot[13].f.lower[30] );
tran (\sa_snapshot[13][31] , \sa_snapshot[13].r.part0[31] );
tran (\sa_snapshot[13][31] , \sa_snapshot[13].f.lower[31] );
tran (\sa_snapshot[13][32] , \sa_snapshot[13].r.part1[0] );
tran (\sa_snapshot[13][32] , \sa_snapshot[13].f.upper[0] );
tran (\sa_snapshot[13][33] , \sa_snapshot[13].r.part1[1] );
tran (\sa_snapshot[13][33] , \sa_snapshot[13].f.upper[1] );
tran (\sa_snapshot[13][34] , \sa_snapshot[13].r.part1[2] );
tran (\sa_snapshot[13][34] , \sa_snapshot[13].f.upper[2] );
tran (\sa_snapshot[13][35] , \sa_snapshot[13].r.part1[3] );
tran (\sa_snapshot[13][35] , \sa_snapshot[13].f.upper[3] );
tran (\sa_snapshot[13][36] , \sa_snapshot[13].r.part1[4] );
tran (\sa_snapshot[13][36] , \sa_snapshot[13].f.upper[4] );
tran (\sa_snapshot[13][37] , \sa_snapshot[13].r.part1[5] );
tran (\sa_snapshot[13][37] , \sa_snapshot[13].f.upper[5] );
tran (\sa_snapshot[13][38] , \sa_snapshot[13].r.part1[6] );
tran (\sa_snapshot[13][38] , \sa_snapshot[13].f.upper[6] );
tran (\sa_snapshot[13][39] , \sa_snapshot[13].r.part1[7] );
tran (\sa_snapshot[13][39] , \sa_snapshot[13].f.upper[7] );
tran (\sa_snapshot[13][40] , \sa_snapshot[13].r.part1[8] );
tran (\sa_snapshot[13][40] , \sa_snapshot[13].f.upper[8] );
tran (\sa_snapshot[13][41] , \sa_snapshot[13].r.part1[9] );
tran (\sa_snapshot[13][41] , \sa_snapshot[13].f.upper[9] );
tran (\sa_snapshot[13][42] , \sa_snapshot[13].r.part1[10] );
tran (\sa_snapshot[13][42] , \sa_snapshot[13].f.upper[10] );
tran (\sa_snapshot[13][43] , \sa_snapshot[13].r.part1[11] );
tran (\sa_snapshot[13][43] , \sa_snapshot[13].f.upper[11] );
tran (\sa_snapshot[13][44] , \sa_snapshot[13].r.part1[12] );
tran (\sa_snapshot[13][44] , \sa_snapshot[13].f.upper[12] );
tran (\sa_snapshot[13][45] , \sa_snapshot[13].r.part1[13] );
tran (\sa_snapshot[13][45] , \sa_snapshot[13].f.upper[13] );
tran (\sa_snapshot[13][46] , \sa_snapshot[13].r.part1[14] );
tran (\sa_snapshot[13][46] , \sa_snapshot[13].f.upper[14] );
tran (\sa_snapshot[13][47] , \sa_snapshot[13].r.part1[15] );
tran (\sa_snapshot[13][47] , \sa_snapshot[13].f.upper[15] );
tran (\sa_snapshot[13][48] , \sa_snapshot[13].r.part1[16] );
tran (\sa_snapshot[13][48] , \sa_snapshot[13].f.upper[16] );
tran (\sa_snapshot[13][49] , \sa_snapshot[13].r.part1[17] );
tran (\sa_snapshot[13][49] , \sa_snapshot[13].f.upper[17] );
tran (\sa_snapshot[13][50] , \sa_snapshot[13].r.part1[18] );
tran (\sa_snapshot[13][50] , \sa_snapshot[13].f.unused[0] );
tran (\sa_snapshot[13][51] , \sa_snapshot[13].r.part1[19] );
tran (\sa_snapshot[13][51] , \sa_snapshot[13].f.unused[1] );
tran (\sa_snapshot[13][52] , \sa_snapshot[13].r.part1[20] );
tran (\sa_snapshot[13][52] , \sa_snapshot[13].f.unused[2] );
tran (\sa_snapshot[13][53] , \sa_snapshot[13].r.part1[21] );
tran (\sa_snapshot[13][53] , \sa_snapshot[13].f.unused[3] );
tran (\sa_snapshot[13][54] , \sa_snapshot[13].r.part1[22] );
tran (\sa_snapshot[13][54] , \sa_snapshot[13].f.unused[4] );
tran (\sa_snapshot[13][55] , \sa_snapshot[13].r.part1[23] );
tran (\sa_snapshot[13][55] , \sa_snapshot[13].f.unused[5] );
tran (\sa_snapshot[13][56] , \sa_snapshot[13].r.part1[24] );
tran (\sa_snapshot[13][56] , \sa_snapshot[13].f.unused[6] );
tran (\sa_snapshot[13][57] , \sa_snapshot[13].r.part1[25] );
tran (\sa_snapshot[13][57] , \sa_snapshot[13].f.unused[7] );
tran (\sa_snapshot[13][58] , \sa_snapshot[13].r.part1[26] );
tran (\sa_snapshot[13][58] , \sa_snapshot[13].f.unused[8] );
tran (\sa_snapshot[13][59] , \sa_snapshot[13].r.part1[27] );
tran (\sa_snapshot[13][59] , \sa_snapshot[13].f.unused[9] );
tran (\sa_snapshot[13][60] , \sa_snapshot[13].r.part1[28] );
tran (\sa_snapshot[13][60] , \sa_snapshot[13].f.unused[10] );
tran (\sa_snapshot[13][61] , \sa_snapshot[13].r.part1[29] );
tran (\sa_snapshot[13][61] , \sa_snapshot[13].f.unused[11] );
tran (\sa_snapshot[13][62] , \sa_snapshot[13].r.part1[30] );
tran (\sa_snapshot[13][62] , \sa_snapshot[13].f.unused[12] );
tran (\sa_snapshot[13][63] , \sa_snapshot[13].r.part1[31] );
tran (\sa_snapshot[13][63] , \sa_snapshot[13].f.unused[13] );
tran (\sa_snapshot[14][0] , \sa_snapshot[14].r.part0[0] );
tran (\sa_snapshot[14][0] , \sa_snapshot[14].f.lower[0] );
tran (\sa_snapshot[14][1] , \sa_snapshot[14].r.part0[1] );
tran (\sa_snapshot[14][1] , \sa_snapshot[14].f.lower[1] );
tran (\sa_snapshot[14][2] , \sa_snapshot[14].r.part0[2] );
tran (\sa_snapshot[14][2] , \sa_snapshot[14].f.lower[2] );
tran (\sa_snapshot[14][3] , \sa_snapshot[14].r.part0[3] );
tran (\sa_snapshot[14][3] , \sa_snapshot[14].f.lower[3] );
tran (\sa_snapshot[14][4] , \sa_snapshot[14].r.part0[4] );
tran (\sa_snapshot[14][4] , \sa_snapshot[14].f.lower[4] );
tran (\sa_snapshot[14][5] , \sa_snapshot[14].r.part0[5] );
tran (\sa_snapshot[14][5] , \sa_snapshot[14].f.lower[5] );
tran (\sa_snapshot[14][6] , \sa_snapshot[14].r.part0[6] );
tran (\sa_snapshot[14][6] , \sa_snapshot[14].f.lower[6] );
tran (\sa_snapshot[14][7] , \sa_snapshot[14].r.part0[7] );
tran (\sa_snapshot[14][7] , \sa_snapshot[14].f.lower[7] );
tran (\sa_snapshot[14][8] , \sa_snapshot[14].r.part0[8] );
tran (\sa_snapshot[14][8] , \sa_snapshot[14].f.lower[8] );
tran (\sa_snapshot[14][9] , \sa_snapshot[14].r.part0[9] );
tran (\sa_snapshot[14][9] , \sa_snapshot[14].f.lower[9] );
tran (\sa_snapshot[14][10] , \sa_snapshot[14].r.part0[10] );
tran (\sa_snapshot[14][10] , \sa_snapshot[14].f.lower[10] );
tran (\sa_snapshot[14][11] , \sa_snapshot[14].r.part0[11] );
tran (\sa_snapshot[14][11] , \sa_snapshot[14].f.lower[11] );
tran (\sa_snapshot[14][12] , \sa_snapshot[14].r.part0[12] );
tran (\sa_snapshot[14][12] , \sa_snapshot[14].f.lower[12] );
tran (\sa_snapshot[14][13] , \sa_snapshot[14].r.part0[13] );
tran (\sa_snapshot[14][13] , \sa_snapshot[14].f.lower[13] );
tran (\sa_snapshot[14][14] , \sa_snapshot[14].r.part0[14] );
tran (\sa_snapshot[14][14] , \sa_snapshot[14].f.lower[14] );
tran (\sa_snapshot[14][15] , \sa_snapshot[14].r.part0[15] );
tran (\sa_snapshot[14][15] , \sa_snapshot[14].f.lower[15] );
tran (\sa_snapshot[14][16] , \sa_snapshot[14].r.part0[16] );
tran (\sa_snapshot[14][16] , \sa_snapshot[14].f.lower[16] );
tran (\sa_snapshot[14][17] , \sa_snapshot[14].r.part0[17] );
tran (\sa_snapshot[14][17] , \sa_snapshot[14].f.lower[17] );
tran (\sa_snapshot[14][18] , \sa_snapshot[14].r.part0[18] );
tran (\sa_snapshot[14][18] , \sa_snapshot[14].f.lower[18] );
tran (\sa_snapshot[14][19] , \sa_snapshot[14].r.part0[19] );
tran (\sa_snapshot[14][19] , \sa_snapshot[14].f.lower[19] );
tran (\sa_snapshot[14][20] , \sa_snapshot[14].r.part0[20] );
tran (\sa_snapshot[14][20] , \sa_snapshot[14].f.lower[20] );
tran (\sa_snapshot[14][21] , \sa_snapshot[14].r.part0[21] );
tran (\sa_snapshot[14][21] , \sa_snapshot[14].f.lower[21] );
tran (\sa_snapshot[14][22] , \sa_snapshot[14].r.part0[22] );
tran (\sa_snapshot[14][22] , \sa_snapshot[14].f.lower[22] );
tran (\sa_snapshot[14][23] , \sa_snapshot[14].r.part0[23] );
tran (\sa_snapshot[14][23] , \sa_snapshot[14].f.lower[23] );
tran (\sa_snapshot[14][24] , \sa_snapshot[14].r.part0[24] );
tran (\sa_snapshot[14][24] , \sa_snapshot[14].f.lower[24] );
tran (\sa_snapshot[14][25] , \sa_snapshot[14].r.part0[25] );
tran (\sa_snapshot[14][25] , \sa_snapshot[14].f.lower[25] );
tran (\sa_snapshot[14][26] , \sa_snapshot[14].r.part0[26] );
tran (\sa_snapshot[14][26] , \sa_snapshot[14].f.lower[26] );
tran (\sa_snapshot[14][27] , \sa_snapshot[14].r.part0[27] );
tran (\sa_snapshot[14][27] , \sa_snapshot[14].f.lower[27] );
tran (\sa_snapshot[14][28] , \sa_snapshot[14].r.part0[28] );
tran (\sa_snapshot[14][28] , \sa_snapshot[14].f.lower[28] );
tran (\sa_snapshot[14][29] , \sa_snapshot[14].r.part0[29] );
tran (\sa_snapshot[14][29] , \sa_snapshot[14].f.lower[29] );
tran (\sa_snapshot[14][30] , \sa_snapshot[14].r.part0[30] );
tran (\sa_snapshot[14][30] , \sa_snapshot[14].f.lower[30] );
tran (\sa_snapshot[14][31] , \sa_snapshot[14].r.part0[31] );
tran (\sa_snapshot[14][31] , \sa_snapshot[14].f.lower[31] );
tran (\sa_snapshot[14][32] , \sa_snapshot[14].r.part1[0] );
tran (\sa_snapshot[14][32] , \sa_snapshot[14].f.upper[0] );
tran (\sa_snapshot[14][33] , \sa_snapshot[14].r.part1[1] );
tran (\sa_snapshot[14][33] , \sa_snapshot[14].f.upper[1] );
tran (\sa_snapshot[14][34] , \sa_snapshot[14].r.part1[2] );
tran (\sa_snapshot[14][34] , \sa_snapshot[14].f.upper[2] );
tran (\sa_snapshot[14][35] , \sa_snapshot[14].r.part1[3] );
tran (\sa_snapshot[14][35] , \sa_snapshot[14].f.upper[3] );
tran (\sa_snapshot[14][36] , \sa_snapshot[14].r.part1[4] );
tran (\sa_snapshot[14][36] , \sa_snapshot[14].f.upper[4] );
tran (\sa_snapshot[14][37] , \sa_snapshot[14].r.part1[5] );
tran (\sa_snapshot[14][37] , \sa_snapshot[14].f.upper[5] );
tran (\sa_snapshot[14][38] , \sa_snapshot[14].r.part1[6] );
tran (\sa_snapshot[14][38] , \sa_snapshot[14].f.upper[6] );
tran (\sa_snapshot[14][39] , \sa_snapshot[14].r.part1[7] );
tran (\sa_snapshot[14][39] , \sa_snapshot[14].f.upper[7] );
tran (\sa_snapshot[14][40] , \sa_snapshot[14].r.part1[8] );
tran (\sa_snapshot[14][40] , \sa_snapshot[14].f.upper[8] );
tran (\sa_snapshot[14][41] , \sa_snapshot[14].r.part1[9] );
tran (\sa_snapshot[14][41] , \sa_snapshot[14].f.upper[9] );
tran (\sa_snapshot[14][42] , \sa_snapshot[14].r.part1[10] );
tran (\sa_snapshot[14][42] , \sa_snapshot[14].f.upper[10] );
tran (\sa_snapshot[14][43] , \sa_snapshot[14].r.part1[11] );
tran (\sa_snapshot[14][43] , \sa_snapshot[14].f.upper[11] );
tran (\sa_snapshot[14][44] , \sa_snapshot[14].r.part1[12] );
tran (\sa_snapshot[14][44] , \sa_snapshot[14].f.upper[12] );
tran (\sa_snapshot[14][45] , \sa_snapshot[14].r.part1[13] );
tran (\sa_snapshot[14][45] , \sa_snapshot[14].f.upper[13] );
tran (\sa_snapshot[14][46] , \sa_snapshot[14].r.part1[14] );
tran (\sa_snapshot[14][46] , \sa_snapshot[14].f.upper[14] );
tran (\sa_snapshot[14][47] , \sa_snapshot[14].r.part1[15] );
tran (\sa_snapshot[14][47] , \sa_snapshot[14].f.upper[15] );
tran (\sa_snapshot[14][48] , \sa_snapshot[14].r.part1[16] );
tran (\sa_snapshot[14][48] , \sa_snapshot[14].f.upper[16] );
tran (\sa_snapshot[14][49] , \sa_snapshot[14].r.part1[17] );
tran (\sa_snapshot[14][49] , \sa_snapshot[14].f.upper[17] );
tran (\sa_snapshot[14][50] , \sa_snapshot[14].r.part1[18] );
tran (\sa_snapshot[14][50] , \sa_snapshot[14].f.unused[0] );
tran (\sa_snapshot[14][51] , \sa_snapshot[14].r.part1[19] );
tran (\sa_snapshot[14][51] , \sa_snapshot[14].f.unused[1] );
tran (\sa_snapshot[14][52] , \sa_snapshot[14].r.part1[20] );
tran (\sa_snapshot[14][52] , \sa_snapshot[14].f.unused[2] );
tran (\sa_snapshot[14][53] , \sa_snapshot[14].r.part1[21] );
tran (\sa_snapshot[14][53] , \sa_snapshot[14].f.unused[3] );
tran (\sa_snapshot[14][54] , \sa_snapshot[14].r.part1[22] );
tran (\sa_snapshot[14][54] , \sa_snapshot[14].f.unused[4] );
tran (\sa_snapshot[14][55] , \sa_snapshot[14].r.part1[23] );
tran (\sa_snapshot[14][55] , \sa_snapshot[14].f.unused[5] );
tran (\sa_snapshot[14][56] , \sa_snapshot[14].r.part1[24] );
tran (\sa_snapshot[14][56] , \sa_snapshot[14].f.unused[6] );
tran (\sa_snapshot[14][57] , \sa_snapshot[14].r.part1[25] );
tran (\sa_snapshot[14][57] , \sa_snapshot[14].f.unused[7] );
tran (\sa_snapshot[14][58] , \sa_snapshot[14].r.part1[26] );
tran (\sa_snapshot[14][58] , \sa_snapshot[14].f.unused[8] );
tran (\sa_snapshot[14][59] , \sa_snapshot[14].r.part1[27] );
tran (\sa_snapshot[14][59] , \sa_snapshot[14].f.unused[9] );
tran (\sa_snapshot[14][60] , \sa_snapshot[14].r.part1[28] );
tran (\sa_snapshot[14][60] , \sa_snapshot[14].f.unused[10] );
tran (\sa_snapshot[14][61] , \sa_snapshot[14].r.part1[29] );
tran (\sa_snapshot[14][61] , \sa_snapshot[14].f.unused[11] );
tran (\sa_snapshot[14][62] , \sa_snapshot[14].r.part1[30] );
tran (\sa_snapshot[14][62] , \sa_snapshot[14].f.unused[12] );
tran (\sa_snapshot[14][63] , \sa_snapshot[14].r.part1[31] );
tran (\sa_snapshot[14][63] , \sa_snapshot[14].f.unused[13] );
tran (\sa_snapshot[15][0] , \sa_snapshot[15].r.part0[0] );
tran (\sa_snapshot[15][0] , \sa_snapshot[15].f.lower[0] );
tran (\sa_snapshot[15][1] , \sa_snapshot[15].r.part0[1] );
tran (\sa_snapshot[15][1] , \sa_snapshot[15].f.lower[1] );
tran (\sa_snapshot[15][2] , \sa_snapshot[15].r.part0[2] );
tran (\sa_snapshot[15][2] , \sa_snapshot[15].f.lower[2] );
tran (\sa_snapshot[15][3] , \sa_snapshot[15].r.part0[3] );
tran (\sa_snapshot[15][3] , \sa_snapshot[15].f.lower[3] );
tran (\sa_snapshot[15][4] , \sa_snapshot[15].r.part0[4] );
tran (\sa_snapshot[15][4] , \sa_snapshot[15].f.lower[4] );
tran (\sa_snapshot[15][5] , \sa_snapshot[15].r.part0[5] );
tran (\sa_snapshot[15][5] , \sa_snapshot[15].f.lower[5] );
tran (\sa_snapshot[15][6] , \sa_snapshot[15].r.part0[6] );
tran (\sa_snapshot[15][6] , \sa_snapshot[15].f.lower[6] );
tran (\sa_snapshot[15][7] , \sa_snapshot[15].r.part0[7] );
tran (\sa_snapshot[15][7] , \sa_snapshot[15].f.lower[7] );
tran (\sa_snapshot[15][8] , \sa_snapshot[15].r.part0[8] );
tran (\sa_snapshot[15][8] , \sa_snapshot[15].f.lower[8] );
tran (\sa_snapshot[15][9] , \sa_snapshot[15].r.part0[9] );
tran (\sa_snapshot[15][9] , \sa_snapshot[15].f.lower[9] );
tran (\sa_snapshot[15][10] , \sa_snapshot[15].r.part0[10] );
tran (\sa_snapshot[15][10] , \sa_snapshot[15].f.lower[10] );
tran (\sa_snapshot[15][11] , \sa_snapshot[15].r.part0[11] );
tran (\sa_snapshot[15][11] , \sa_snapshot[15].f.lower[11] );
tran (\sa_snapshot[15][12] , \sa_snapshot[15].r.part0[12] );
tran (\sa_snapshot[15][12] , \sa_snapshot[15].f.lower[12] );
tran (\sa_snapshot[15][13] , \sa_snapshot[15].r.part0[13] );
tran (\sa_snapshot[15][13] , \sa_snapshot[15].f.lower[13] );
tran (\sa_snapshot[15][14] , \sa_snapshot[15].r.part0[14] );
tran (\sa_snapshot[15][14] , \sa_snapshot[15].f.lower[14] );
tran (\sa_snapshot[15][15] , \sa_snapshot[15].r.part0[15] );
tran (\sa_snapshot[15][15] , \sa_snapshot[15].f.lower[15] );
tran (\sa_snapshot[15][16] , \sa_snapshot[15].r.part0[16] );
tran (\sa_snapshot[15][16] , \sa_snapshot[15].f.lower[16] );
tran (\sa_snapshot[15][17] , \sa_snapshot[15].r.part0[17] );
tran (\sa_snapshot[15][17] , \sa_snapshot[15].f.lower[17] );
tran (\sa_snapshot[15][18] , \sa_snapshot[15].r.part0[18] );
tran (\sa_snapshot[15][18] , \sa_snapshot[15].f.lower[18] );
tran (\sa_snapshot[15][19] , \sa_snapshot[15].r.part0[19] );
tran (\sa_snapshot[15][19] , \sa_snapshot[15].f.lower[19] );
tran (\sa_snapshot[15][20] , \sa_snapshot[15].r.part0[20] );
tran (\sa_snapshot[15][20] , \sa_snapshot[15].f.lower[20] );
tran (\sa_snapshot[15][21] , \sa_snapshot[15].r.part0[21] );
tran (\sa_snapshot[15][21] , \sa_snapshot[15].f.lower[21] );
tran (\sa_snapshot[15][22] , \sa_snapshot[15].r.part0[22] );
tran (\sa_snapshot[15][22] , \sa_snapshot[15].f.lower[22] );
tran (\sa_snapshot[15][23] , \sa_snapshot[15].r.part0[23] );
tran (\sa_snapshot[15][23] , \sa_snapshot[15].f.lower[23] );
tran (\sa_snapshot[15][24] , \sa_snapshot[15].r.part0[24] );
tran (\sa_snapshot[15][24] , \sa_snapshot[15].f.lower[24] );
tran (\sa_snapshot[15][25] , \sa_snapshot[15].r.part0[25] );
tran (\sa_snapshot[15][25] , \sa_snapshot[15].f.lower[25] );
tran (\sa_snapshot[15][26] , \sa_snapshot[15].r.part0[26] );
tran (\sa_snapshot[15][26] , \sa_snapshot[15].f.lower[26] );
tran (\sa_snapshot[15][27] , \sa_snapshot[15].r.part0[27] );
tran (\sa_snapshot[15][27] , \sa_snapshot[15].f.lower[27] );
tran (\sa_snapshot[15][28] , \sa_snapshot[15].r.part0[28] );
tran (\sa_snapshot[15][28] , \sa_snapshot[15].f.lower[28] );
tran (\sa_snapshot[15][29] , \sa_snapshot[15].r.part0[29] );
tran (\sa_snapshot[15][29] , \sa_snapshot[15].f.lower[29] );
tran (\sa_snapshot[15][30] , \sa_snapshot[15].r.part0[30] );
tran (\sa_snapshot[15][30] , \sa_snapshot[15].f.lower[30] );
tran (\sa_snapshot[15][31] , \sa_snapshot[15].r.part0[31] );
tran (\sa_snapshot[15][31] , \sa_snapshot[15].f.lower[31] );
tran (\sa_snapshot[15][32] , \sa_snapshot[15].r.part1[0] );
tran (\sa_snapshot[15][32] , \sa_snapshot[15].f.upper[0] );
tran (\sa_snapshot[15][33] , \sa_snapshot[15].r.part1[1] );
tran (\sa_snapshot[15][33] , \sa_snapshot[15].f.upper[1] );
tran (\sa_snapshot[15][34] , \sa_snapshot[15].r.part1[2] );
tran (\sa_snapshot[15][34] , \sa_snapshot[15].f.upper[2] );
tran (\sa_snapshot[15][35] , \sa_snapshot[15].r.part1[3] );
tran (\sa_snapshot[15][35] , \sa_snapshot[15].f.upper[3] );
tran (\sa_snapshot[15][36] , \sa_snapshot[15].r.part1[4] );
tran (\sa_snapshot[15][36] , \sa_snapshot[15].f.upper[4] );
tran (\sa_snapshot[15][37] , \sa_snapshot[15].r.part1[5] );
tran (\sa_snapshot[15][37] , \sa_snapshot[15].f.upper[5] );
tran (\sa_snapshot[15][38] , \sa_snapshot[15].r.part1[6] );
tran (\sa_snapshot[15][38] , \sa_snapshot[15].f.upper[6] );
tran (\sa_snapshot[15][39] , \sa_snapshot[15].r.part1[7] );
tran (\sa_snapshot[15][39] , \sa_snapshot[15].f.upper[7] );
tran (\sa_snapshot[15][40] , \sa_snapshot[15].r.part1[8] );
tran (\sa_snapshot[15][40] , \sa_snapshot[15].f.upper[8] );
tran (\sa_snapshot[15][41] , \sa_snapshot[15].r.part1[9] );
tran (\sa_snapshot[15][41] , \sa_snapshot[15].f.upper[9] );
tran (\sa_snapshot[15][42] , \sa_snapshot[15].r.part1[10] );
tran (\sa_snapshot[15][42] , \sa_snapshot[15].f.upper[10] );
tran (\sa_snapshot[15][43] , \sa_snapshot[15].r.part1[11] );
tran (\sa_snapshot[15][43] , \sa_snapshot[15].f.upper[11] );
tran (\sa_snapshot[15][44] , \sa_snapshot[15].r.part1[12] );
tran (\sa_snapshot[15][44] , \sa_snapshot[15].f.upper[12] );
tran (\sa_snapshot[15][45] , \sa_snapshot[15].r.part1[13] );
tran (\sa_snapshot[15][45] , \sa_snapshot[15].f.upper[13] );
tran (\sa_snapshot[15][46] , \sa_snapshot[15].r.part1[14] );
tran (\sa_snapshot[15][46] , \sa_snapshot[15].f.upper[14] );
tran (\sa_snapshot[15][47] , \sa_snapshot[15].r.part1[15] );
tran (\sa_snapshot[15][47] , \sa_snapshot[15].f.upper[15] );
tran (\sa_snapshot[15][48] , \sa_snapshot[15].r.part1[16] );
tran (\sa_snapshot[15][48] , \sa_snapshot[15].f.upper[16] );
tran (\sa_snapshot[15][49] , \sa_snapshot[15].r.part1[17] );
tran (\sa_snapshot[15][49] , \sa_snapshot[15].f.upper[17] );
tran (\sa_snapshot[15][50] , \sa_snapshot[15].r.part1[18] );
tran (\sa_snapshot[15][50] , \sa_snapshot[15].f.unused[0] );
tran (\sa_snapshot[15][51] , \sa_snapshot[15].r.part1[19] );
tran (\sa_snapshot[15][51] , \sa_snapshot[15].f.unused[1] );
tran (\sa_snapshot[15][52] , \sa_snapshot[15].r.part1[20] );
tran (\sa_snapshot[15][52] , \sa_snapshot[15].f.unused[2] );
tran (\sa_snapshot[15][53] , \sa_snapshot[15].r.part1[21] );
tran (\sa_snapshot[15][53] , \sa_snapshot[15].f.unused[3] );
tran (\sa_snapshot[15][54] , \sa_snapshot[15].r.part1[22] );
tran (\sa_snapshot[15][54] , \sa_snapshot[15].f.unused[4] );
tran (\sa_snapshot[15][55] , \sa_snapshot[15].r.part1[23] );
tran (\sa_snapshot[15][55] , \sa_snapshot[15].f.unused[5] );
tran (\sa_snapshot[15][56] , \sa_snapshot[15].r.part1[24] );
tran (\sa_snapshot[15][56] , \sa_snapshot[15].f.unused[6] );
tran (\sa_snapshot[15][57] , \sa_snapshot[15].r.part1[25] );
tran (\sa_snapshot[15][57] , \sa_snapshot[15].f.unused[7] );
tran (\sa_snapshot[15][58] , \sa_snapshot[15].r.part1[26] );
tran (\sa_snapshot[15][58] , \sa_snapshot[15].f.unused[8] );
tran (\sa_snapshot[15][59] , \sa_snapshot[15].r.part1[27] );
tran (\sa_snapshot[15][59] , \sa_snapshot[15].f.unused[9] );
tran (\sa_snapshot[15][60] , \sa_snapshot[15].r.part1[28] );
tran (\sa_snapshot[15][60] , \sa_snapshot[15].f.unused[10] );
tran (\sa_snapshot[15][61] , \sa_snapshot[15].r.part1[29] );
tran (\sa_snapshot[15][61] , \sa_snapshot[15].f.unused[11] );
tran (\sa_snapshot[15][62] , \sa_snapshot[15].r.part1[30] );
tran (\sa_snapshot[15][62] , \sa_snapshot[15].f.unused[12] );
tran (\sa_snapshot[15][63] , \sa_snapshot[15].r.part1[31] );
tran (\sa_snapshot[15][63] , \sa_snapshot[15].f.unused[13] );
tran (\sa_snapshot[16][0] , \sa_snapshot[16].r.part0[0] );
tran (\sa_snapshot[16][0] , \sa_snapshot[16].f.lower[0] );
tran (\sa_snapshot[16][1] , \sa_snapshot[16].r.part0[1] );
tran (\sa_snapshot[16][1] , \sa_snapshot[16].f.lower[1] );
tran (\sa_snapshot[16][2] , \sa_snapshot[16].r.part0[2] );
tran (\sa_snapshot[16][2] , \sa_snapshot[16].f.lower[2] );
tran (\sa_snapshot[16][3] , \sa_snapshot[16].r.part0[3] );
tran (\sa_snapshot[16][3] , \sa_snapshot[16].f.lower[3] );
tran (\sa_snapshot[16][4] , \sa_snapshot[16].r.part0[4] );
tran (\sa_snapshot[16][4] , \sa_snapshot[16].f.lower[4] );
tran (\sa_snapshot[16][5] , \sa_snapshot[16].r.part0[5] );
tran (\sa_snapshot[16][5] , \sa_snapshot[16].f.lower[5] );
tran (\sa_snapshot[16][6] , \sa_snapshot[16].r.part0[6] );
tran (\sa_snapshot[16][6] , \sa_snapshot[16].f.lower[6] );
tran (\sa_snapshot[16][7] , \sa_snapshot[16].r.part0[7] );
tran (\sa_snapshot[16][7] , \sa_snapshot[16].f.lower[7] );
tran (\sa_snapshot[16][8] , \sa_snapshot[16].r.part0[8] );
tran (\sa_snapshot[16][8] , \sa_snapshot[16].f.lower[8] );
tran (\sa_snapshot[16][9] , \sa_snapshot[16].r.part0[9] );
tran (\sa_snapshot[16][9] , \sa_snapshot[16].f.lower[9] );
tran (\sa_snapshot[16][10] , \sa_snapshot[16].r.part0[10] );
tran (\sa_snapshot[16][10] , \sa_snapshot[16].f.lower[10] );
tran (\sa_snapshot[16][11] , \sa_snapshot[16].r.part0[11] );
tran (\sa_snapshot[16][11] , \sa_snapshot[16].f.lower[11] );
tran (\sa_snapshot[16][12] , \sa_snapshot[16].r.part0[12] );
tran (\sa_snapshot[16][12] , \sa_snapshot[16].f.lower[12] );
tran (\sa_snapshot[16][13] , \sa_snapshot[16].r.part0[13] );
tran (\sa_snapshot[16][13] , \sa_snapshot[16].f.lower[13] );
tran (\sa_snapshot[16][14] , \sa_snapshot[16].r.part0[14] );
tran (\sa_snapshot[16][14] , \sa_snapshot[16].f.lower[14] );
tran (\sa_snapshot[16][15] , \sa_snapshot[16].r.part0[15] );
tran (\sa_snapshot[16][15] , \sa_snapshot[16].f.lower[15] );
tran (\sa_snapshot[16][16] , \sa_snapshot[16].r.part0[16] );
tran (\sa_snapshot[16][16] , \sa_snapshot[16].f.lower[16] );
tran (\sa_snapshot[16][17] , \sa_snapshot[16].r.part0[17] );
tran (\sa_snapshot[16][17] , \sa_snapshot[16].f.lower[17] );
tran (\sa_snapshot[16][18] , \sa_snapshot[16].r.part0[18] );
tran (\sa_snapshot[16][18] , \sa_snapshot[16].f.lower[18] );
tran (\sa_snapshot[16][19] , \sa_snapshot[16].r.part0[19] );
tran (\sa_snapshot[16][19] , \sa_snapshot[16].f.lower[19] );
tran (\sa_snapshot[16][20] , \sa_snapshot[16].r.part0[20] );
tran (\sa_snapshot[16][20] , \sa_snapshot[16].f.lower[20] );
tran (\sa_snapshot[16][21] , \sa_snapshot[16].r.part0[21] );
tran (\sa_snapshot[16][21] , \sa_snapshot[16].f.lower[21] );
tran (\sa_snapshot[16][22] , \sa_snapshot[16].r.part0[22] );
tran (\sa_snapshot[16][22] , \sa_snapshot[16].f.lower[22] );
tran (\sa_snapshot[16][23] , \sa_snapshot[16].r.part0[23] );
tran (\sa_snapshot[16][23] , \sa_snapshot[16].f.lower[23] );
tran (\sa_snapshot[16][24] , \sa_snapshot[16].r.part0[24] );
tran (\sa_snapshot[16][24] , \sa_snapshot[16].f.lower[24] );
tran (\sa_snapshot[16][25] , \sa_snapshot[16].r.part0[25] );
tran (\sa_snapshot[16][25] , \sa_snapshot[16].f.lower[25] );
tran (\sa_snapshot[16][26] , \sa_snapshot[16].r.part0[26] );
tran (\sa_snapshot[16][26] , \sa_snapshot[16].f.lower[26] );
tran (\sa_snapshot[16][27] , \sa_snapshot[16].r.part0[27] );
tran (\sa_snapshot[16][27] , \sa_snapshot[16].f.lower[27] );
tran (\sa_snapshot[16][28] , \sa_snapshot[16].r.part0[28] );
tran (\sa_snapshot[16][28] , \sa_snapshot[16].f.lower[28] );
tran (\sa_snapshot[16][29] , \sa_snapshot[16].r.part0[29] );
tran (\sa_snapshot[16][29] , \sa_snapshot[16].f.lower[29] );
tran (\sa_snapshot[16][30] , \sa_snapshot[16].r.part0[30] );
tran (\sa_snapshot[16][30] , \sa_snapshot[16].f.lower[30] );
tran (\sa_snapshot[16][31] , \sa_snapshot[16].r.part0[31] );
tran (\sa_snapshot[16][31] , \sa_snapshot[16].f.lower[31] );
tran (\sa_snapshot[16][32] , \sa_snapshot[16].r.part1[0] );
tran (\sa_snapshot[16][32] , \sa_snapshot[16].f.upper[0] );
tran (\sa_snapshot[16][33] , \sa_snapshot[16].r.part1[1] );
tran (\sa_snapshot[16][33] , \sa_snapshot[16].f.upper[1] );
tran (\sa_snapshot[16][34] , \sa_snapshot[16].r.part1[2] );
tran (\sa_snapshot[16][34] , \sa_snapshot[16].f.upper[2] );
tran (\sa_snapshot[16][35] , \sa_snapshot[16].r.part1[3] );
tran (\sa_snapshot[16][35] , \sa_snapshot[16].f.upper[3] );
tran (\sa_snapshot[16][36] , \sa_snapshot[16].r.part1[4] );
tran (\sa_snapshot[16][36] , \sa_snapshot[16].f.upper[4] );
tran (\sa_snapshot[16][37] , \sa_snapshot[16].r.part1[5] );
tran (\sa_snapshot[16][37] , \sa_snapshot[16].f.upper[5] );
tran (\sa_snapshot[16][38] , \sa_snapshot[16].r.part1[6] );
tran (\sa_snapshot[16][38] , \sa_snapshot[16].f.upper[6] );
tran (\sa_snapshot[16][39] , \sa_snapshot[16].r.part1[7] );
tran (\sa_snapshot[16][39] , \sa_snapshot[16].f.upper[7] );
tran (\sa_snapshot[16][40] , \sa_snapshot[16].r.part1[8] );
tran (\sa_snapshot[16][40] , \sa_snapshot[16].f.upper[8] );
tran (\sa_snapshot[16][41] , \sa_snapshot[16].r.part1[9] );
tran (\sa_snapshot[16][41] , \sa_snapshot[16].f.upper[9] );
tran (\sa_snapshot[16][42] , \sa_snapshot[16].r.part1[10] );
tran (\sa_snapshot[16][42] , \sa_snapshot[16].f.upper[10] );
tran (\sa_snapshot[16][43] , \sa_snapshot[16].r.part1[11] );
tran (\sa_snapshot[16][43] , \sa_snapshot[16].f.upper[11] );
tran (\sa_snapshot[16][44] , \sa_snapshot[16].r.part1[12] );
tran (\sa_snapshot[16][44] , \sa_snapshot[16].f.upper[12] );
tran (\sa_snapshot[16][45] , \sa_snapshot[16].r.part1[13] );
tran (\sa_snapshot[16][45] , \sa_snapshot[16].f.upper[13] );
tran (\sa_snapshot[16][46] , \sa_snapshot[16].r.part1[14] );
tran (\sa_snapshot[16][46] , \sa_snapshot[16].f.upper[14] );
tran (\sa_snapshot[16][47] , \sa_snapshot[16].r.part1[15] );
tran (\sa_snapshot[16][47] , \sa_snapshot[16].f.upper[15] );
tran (\sa_snapshot[16][48] , \sa_snapshot[16].r.part1[16] );
tran (\sa_snapshot[16][48] , \sa_snapshot[16].f.upper[16] );
tran (\sa_snapshot[16][49] , \sa_snapshot[16].r.part1[17] );
tran (\sa_snapshot[16][49] , \sa_snapshot[16].f.upper[17] );
tran (\sa_snapshot[16][50] , \sa_snapshot[16].r.part1[18] );
tran (\sa_snapshot[16][50] , \sa_snapshot[16].f.unused[0] );
tran (\sa_snapshot[16][51] , \sa_snapshot[16].r.part1[19] );
tran (\sa_snapshot[16][51] , \sa_snapshot[16].f.unused[1] );
tran (\sa_snapshot[16][52] , \sa_snapshot[16].r.part1[20] );
tran (\sa_snapshot[16][52] , \sa_snapshot[16].f.unused[2] );
tran (\sa_snapshot[16][53] , \sa_snapshot[16].r.part1[21] );
tran (\sa_snapshot[16][53] , \sa_snapshot[16].f.unused[3] );
tran (\sa_snapshot[16][54] , \sa_snapshot[16].r.part1[22] );
tran (\sa_snapshot[16][54] , \sa_snapshot[16].f.unused[4] );
tran (\sa_snapshot[16][55] , \sa_snapshot[16].r.part1[23] );
tran (\sa_snapshot[16][55] , \sa_snapshot[16].f.unused[5] );
tran (\sa_snapshot[16][56] , \sa_snapshot[16].r.part1[24] );
tran (\sa_snapshot[16][56] , \sa_snapshot[16].f.unused[6] );
tran (\sa_snapshot[16][57] , \sa_snapshot[16].r.part1[25] );
tran (\sa_snapshot[16][57] , \sa_snapshot[16].f.unused[7] );
tran (\sa_snapshot[16][58] , \sa_snapshot[16].r.part1[26] );
tran (\sa_snapshot[16][58] , \sa_snapshot[16].f.unused[8] );
tran (\sa_snapshot[16][59] , \sa_snapshot[16].r.part1[27] );
tran (\sa_snapshot[16][59] , \sa_snapshot[16].f.unused[9] );
tran (\sa_snapshot[16][60] , \sa_snapshot[16].r.part1[28] );
tran (\sa_snapshot[16][60] , \sa_snapshot[16].f.unused[10] );
tran (\sa_snapshot[16][61] , \sa_snapshot[16].r.part1[29] );
tran (\sa_snapshot[16][61] , \sa_snapshot[16].f.unused[11] );
tran (\sa_snapshot[16][62] , \sa_snapshot[16].r.part1[30] );
tran (\sa_snapshot[16][62] , \sa_snapshot[16].f.unused[12] );
tran (\sa_snapshot[16][63] , \sa_snapshot[16].r.part1[31] );
tran (\sa_snapshot[16][63] , \sa_snapshot[16].f.unused[13] );
tran (\sa_snapshot[17][0] , \sa_snapshot[17].r.part0[0] );
tran (\sa_snapshot[17][0] , \sa_snapshot[17].f.lower[0] );
tran (\sa_snapshot[17][1] , \sa_snapshot[17].r.part0[1] );
tran (\sa_snapshot[17][1] , \sa_snapshot[17].f.lower[1] );
tran (\sa_snapshot[17][2] , \sa_snapshot[17].r.part0[2] );
tran (\sa_snapshot[17][2] , \sa_snapshot[17].f.lower[2] );
tran (\sa_snapshot[17][3] , \sa_snapshot[17].r.part0[3] );
tran (\sa_snapshot[17][3] , \sa_snapshot[17].f.lower[3] );
tran (\sa_snapshot[17][4] , \sa_snapshot[17].r.part0[4] );
tran (\sa_snapshot[17][4] , \sa_snapshot[17].f.lower[4] );
tran (\sa_snapshot[17][5] , \sa_snapshot[17].r.part0[5] );
tran (\sa_snapshot[17][5] , \sa_snapshot[17].f.lower[5] );
tran (\sa_snapshot[17][6] , \sa_snapshot[17].r.part0[6] );
tran (\sa_snapshot[17][6] , \sa_snapshot[17].f.lower[6] );
tran (\sa_snapshot[17][7] , \sa_snapshot[17].r.part0[7] );
tran (\sa_snapshot[17][7] , \sa_snapshot[17].f.lower[7] );
tran (\sa_snapshot[17][8] , \sa_snapshot[17].r.part0[8] );
tran (\sa_snapshot[17][8] , \sa_snapshot[17].f.lower[8] );
tran (\sa_snapshot[17][9] , \sa_snapshot[17].r.part0[9] );
tran (\sa_snapshot[17][9] , \sa_snapshot[17].f.lower[9] );
tran (\sa_snapshot[17][10] , \sa_snapshot[17].r.part0[10] );
tran (\sa_snapshot[17][10] , \sa_snapshot[17].f.lower[10] );
tran (\sa_snapshot[17][11] , \sa_snapshot[17].r.part0[11] );
tran (\sa_snapshot[17][11] , \sa_snapshot[17].f.lower[11] );
tran (\sa_snapshot[17][12] , \sa_snapshot[17].r.part0[12] );
tran (\sa_snapshot[17][12] , \sa_snapshot[17].f.lower[12] );
tran (\sa_snapshot[17][13] , \sa_snapshot[17].r.part0[13] );
tran (\sa_snapshot[17][13] , \sa_snapshot[17].f.lower[13] );
tran (\sa_snapshot[17][14] , \sa_snapshot[17].r.part0[14] );
tran (\sa_snapshot[17][14] , \sa_snapshot[17].f.lower[14] );
tran (\sa_snapshot[17][15] , \sa_snapshot[17].r.part0[15] );
tran (\sa_snapshot[17][15] , \sa_snapshot[17].f.lower[15] );
tran (\sa_snapshot[17][16] , \sa_snapshot[17].r.part0[16] );
tran (\sa_snapshot[17][16] , \sa_snapshot[17].f.lower[16] );
tran (\sa_snapshot[17][17] , \sa_snapshot[17].r.part0[17] );
tran (\sa_snapshot[17][17] , \sa_snapshot[17].f.lower[17] );
tran (\sa_snapshot[17][18] , \sa_snapshot[17].r.part0[18] );
tran (\sa_snapshot[17][18] , \sa_snapshot[17].f.lower[18] );
tran (\sa_snapshot[17][19] , \sa_snapshot[17].r.part0[19] );
tran (\sa_snapshot[17][19] , \sa_snapshot[17].f.lower[19] );
tran (\sa_snapshot[17][20] , \sa_snapshot[17].r.part0[20] );
tran (\sa_snapshot[17][20] , \sa_snapshot[17].f.lower[20] );
tran (\sa_snapshot[17][21] , \sa_snapshot[17].r.part0[21] );
tran (\sa_snapshot[17][21] , \sa_snapshot[17].f.lower[21] );
tran (\sa_snapshot[17][22] , \sa_snapshot[17].r.part0[22] );
tran (\sa_snapshot[17][22] , \sa_snapshot[17].f.lower[22] );
tran (\sa_snapshot[17][23] , \sa_snapshot[17].r.part0[23] );
tran (\sa_snapshot[17][23] , \sa_snapshot[17].f.lower[23] );
tran (\sa_snapshot[17][24] , \sa_snapshot[17].r.part0[24] );
tran (\sa_snapshot[17][24] , \sa_snapshot[17].f.lower[24] );
tran (\sa_snapshot[17][25] , \sa_snapshot[17].r.part0[25] );
tran (\sa_snapshot[17][25] , \sa_snapshot[17].f.lower[25] );
tran (\sa_snapshot[17][26] , \sa_snapshot[17].r.part0[26] );
tran (\sa_snapshot[17][26] , \sa_snapshot[17].f.lower[26] );
tran (\sa_snapshot[17][27] , \sa_snapshot[17].r.part0[27] );
tran (\sa_snapshot[17][27] , \sa_snapshot[17].f.lower[27] );
tran (\sa_snapshot[17][28] , \sa_snapshot[17].r.part0[28] );
tran (\sa_snapshot[17][28] , \sa_snapshot[17].f.lower[28] );
tran (\sa_snapshot[17][29] , \sa_snapshot[17].r.part0[29] );
tran (\sa_snapshot[17][29] , \sa_snapshot[17].f.lower[29] );
tran (\sa_snapshot[17][30] , \sa_snapshot[17].r.part0[30] );
tran (\sa_snapshot[17][30] , \sa_snapshot[17].f.lower[30] );
tran (\sa_snapshot[17][31] , \sa_snapshot[17].r.part0[31] );
tran (\sa_snapshot[17][31] , \sa_snapshot[17].f.lower[31] );
tran (\sa_snapshot[17][32] , \sa_snapshot[17].r.part1[0] );
tran (\sa_snapshot[17][32] , \sa_snapshot[17].f.upper[0] );
tran (\sa_snapshot[17][33] , \sa_snapshot[17].r.part1[1] );
tran (\sa_snapshot[17][33] , \sa_snapshot[17].f.upper[1] );
tran (\sa_snapshot[17][34] , \sa_snapshot[17].r.part1[2] );
tran (\sa_snapshot[17][34] , \sa_snapshot[17].f.upper[2] );
tran (\sa_snapshot[17][35] , \sa_snapshot[17].r.part1[3] );
tran (\sa_snapshot[17][35] , \sa_snapshot[17].f.upper[3] );
tran (\sa_snapshot[17][36] , \sa_snapshot[17].r.part1[4] );
tran (\sa_snapshot[17][36] , \sa_snapshot[17].f.upper[4] );
tran (\sa_snapshot[17][37] , \sa_snapshot[17].r.part1[5] );
tran (\sa_snapshot[17][37] , \sa_snapshot[17].f.upper[5] );
tran (\sa_snapshot[17][38] , \sa_snapshot[17].r.part1[6] );
tran (\sa_snapshot[17][38] , \sa_snapshot[17].f.upper[6] );
tran (\sa_snapshot[17][39] , \sa_snapshot[17].r.part1[7] );
tran (\sa_snapshot[17][39] , \sa_snapshot[17].f.upper[7] );
tran (\sa_snapshot[17][40] , \sa_snapshot[17].r.part1[8] );
tran (\sa_snapshot[17][40] , \sa_snapshot[17].f.upper[8] );
tran (\sa_snapshot[17][41] , \sa_snapshot[17].r.part1[9] );
tran (\sa_snapshot[17][41] , \sa_snapshot[17].f.upper[9] );
tran (\sa_snapshot[17][42] , \sa_snapshot[17].r.part1[10] );
tran (\sa_snapshot[17][42] , \sa_snapshot[17].f.upper[10] );
tran (\sa_snapshot[17][43] , \sa_snapshot[17].r.part1[11] );
tran (\sa_snapshot[17][43] , \sa_snapshot[17].f.upper[11] );
tran (\sa_snapshot[17][44] , \sa_snapshot[17].r.part1[12] );
tran (\sa_snapshot[17][44] , \sa_snapshot[17].f.upper[12] );
tran (\sa_snapshot[17][45] , \sa_snapshot[17].r.part1[13] );
tran (\sa_snapshot[17][45] , \sa_snapshot[17].f.upper[13] );
tran (\sa_snapshot[17][46] , \sa_snapshot[17].r.part1[14] );
tran (\sa_snapshot[17][46] , \sa_snapshot[17].f.upper[14] );
tran (\sa_snapshot[17][47] , \sa_snapshot[17].r.part1[15] );
tran (\sa_snapshot[17][47] , \sa_snapshot[17].f.upper[15] );
tran (\sa_snapshot[17][48] , \sa_snapshot[17].r.part1[16] );
tran (\sa_snapshot[17][48] , \sa_snapshot[17].f.upper[16] );
tran (\sa_snapshot[17][49] , \sa_snapshot[17].r.part1[17] );
tran (\sa_snapshot[17][49] , \sa_snapshot[17].f.upper[17] );
tran (\sa_snapshot[17][50] , \sa_snapshot[17].r.part1[18] );
tran (\sa_snapshot[17][50] , \sa_snapshot[17].f.unused[0] );
tran (\sa_snapshot[17][51] , \sa_snapshot[17].r.part1[19] );
tran (\sa_snapshot[17][51] , \sa_snapshot[17].f.unused[1] );
tran (\sa_snapshot[17][52] , \sa_snapshot[17].r.part1[20] );
tran (\sa_snapshot[17][52] , \sa_snapshot[17].f.unused[2] );
tran (\sa_snapshot[17][53] , \sa_snapshot[17].r.part1[21] );
tran (\sa_snapshot[17][53] , \sa_snapshot[17].f.unused[3] );
tran (\sa_snapshot[17][54] , \sa_snapshot[17].r.part1[22] );
tran (\sa_snapshot[17][54] , \sa_snapshot[17].f.unused[4] );
tran (\sa_snapshot[17][55] , \sa_snapshot[17].r.part1[23] );
tran (\sa_snapshot[17][55] , \sa_snapshot[17].f.unused[5] );
tran (\sa_snapshot[17][56] , \sa_snapshot[17].r.part1[24] );
tran (\sa_snapshot[17][56] , \sa_snapshot[17].f.unused[6] );
tran (\sa_snapshot[17][57] , \sa_snapshot[17].r.part1[25] );
tran (\sa_snapshot[17][57] , \sa_snapshot[17].f.unused[7] );
tran (\sa_snapshot[17][58] , \sa_snapshot[17].r.part1[26] );
tran (\sa_snapshot[17][58] , \sa_snapshot[17].f.unused[8] );
tran (\sa_snapshot[17][59] , \sa_snapshot[17].r.part1[27] );
tran (\sa_snapshot[17][59] , \sa_snapshot[17].f.unused[9] );
tran (\sa_snapshot[17][60] , \sa_snapshot[17].r.part1[28] );
tran (\sa_snapshot[17][60] , \sa_snapshot[17].f.unused[10] );
tran (\sa_snapshot[17][61] , \sa_snapshot[17].r.part1[29] );
tran (\sa_snapshot[17][61] , \sa_snapshot[17].f.unused[11] );
tran (\sa_snapshot[17][62] , \sa_snapshot[17].r.part1[30] );
tran (\sa_snapshot[17][62] , \sa_snapshot[17].f.unused[12] );
tran (\sa_snapshot[17][63] , \sa_snapshot[17].r.part1[31] );
tran (\sa_snapshot[17][63] , \sa_snapshot[17].f.unused[13] );
tran (\sa_snapshot[18][0] , \sa_snapshot[18].r.part0[0] );
tran (\sa_snapshot[18][0] , \sa_snapshot[18].f.lower[0] );
tran (\sa_snapshot[18][1] , \sa_snapshot[18].r.part0[1] );
tran (\sa_snapshot[18][1] , \sa_snapshot[18].f.lower[1] );
tran (\sa_snapshot[18][2] , \sa_snapshot[18].r.part0[2] );
tran (\sa_snapshot[18][2] , \sa_snapshot[18].f.lower[2] );
tran (\sa_snapshot[18][3] , \sa_snapshot[18].r.part0[3] );
tran (\sa_snapshot[18][3] , \sa_snapshot[18].f.lower[3] );
tran (\sa_snapshot[18][4] , \sa_snapshot[18].r.part0[4] );
tran (\sa_snapshot[18][4] , \sa_snapshot[18].f.lower[4] );
tran (\sa_snapshot[18][5] , \sa_snapshot[18].r.part0[5] );
tran (\sa_snapshot[18][5] , \sa_snapshot[18].f.lower[5] );
tran (\sa_snapshot[18][6] , \sa_snapshot[18].r.part0[6] );
tran (\sa_snapshot[18][6] , \sa_snapshot[18].f.lower[6] );
tran (\sa_snapshot[18][7] , \sa_snapshot[18].r.part0[7] );
tran (\sa_snapshot[18][7] , \sa_snapshot[18].f.lower[7] );
tran (\sa_snapshot[18][8] , \sa_snapshot[18].r.part0[8] );
tran (\sa_snapshot[18][8] , \sa_snapshot[18].f.lower[8] );
tran (\sa_snapshot[18][9] , \sa_snapshot[18].r.part0[9] );
tran (\sa_snapshot[18][9] , \sa_snapshot[18].f.lower[9] );
tran (\sa_snapshot[18][10] , \sa_snapshot[18].r.part0[10] );
tran (\sa_snapshot[18][10] , \sa_snapshot[18].f.lower[10] );
tran (\sa_snapshot[18][11] , \sa_snapshot[18].r.part0[11] );
tran (\sa_snapshot[18][11] , \sa_snapshot[18].f.lower[11] );
tran (\sa_snapshot[18][12] , \sa_snapshot[18].r.part0[12] );
tran (\sa_snapshot[18][12] , \sa_snapshot[18].f.lower[12] );
tran (\sa_snapshot[18][13] , \sa_snapshot[18].r.part0[13] );
tran (\sa_snapshot[18][13] , \sa_snapshot[18].f.lower[13] );
tran (\sa_snapshot[18][14] , \sa_snapshot[18].r.part0[14] );
tran (\sa_snapshot[18][14] , \sa_snapshot[18].f.lower[14] );
tran (\sa_snapshot[18][15] , \sa_snapshot[18].r.part0[15] );
tran (\sa_snapshot[18][15] , \sa_snapshot[18].f.lower[15] );
tran (\sa_snapshot[18][16] , \sa_snapshot[18].r.part0[16] );
tran (\sa_snapshot[18][16] , \sa_snapshot[18].f.lower[16] );
tran (\sa_snapshot[18][17] , \sa_snapshot[18].r.part0[17] );
tran (\sa_snapshot[18][17] , \sa_snapshot[18].f.lower[17] );
tran (\sa_snapshot[18][18] , \sa_snapshot[18].r.part0[18] );
tran (\sa_snapshot[18][18] , \sa_snapshot[18].f.lower[18] );
tran (\sa_snapshot[18][19] , \sa_snapshot[18].r.part0[19] );
tran (\sa_snapshot[18][19] , \sa_snapshot[18].f.lower[19] );
tran (\sa_snapshot[18][20] , \sa_snapshot[18].r.part0[20] );
tran (\sa_snapshot[18][20] , \sa_snapshot[18].f.lower[20] );
tran (\sa_snapshot[18][21] , \sa_snapshot[18].r.part0[21] );
tran (\sa_snapshot[18][21] , \sa_snapshot[18].f.lower[21] );
tran (\sa_snapshot[18][22] , \sa_snapshot[18].r.part0[22] );
tran (\sa_snapshot[18][22] , \sa_snapshot[18].f.lower[22] );
tran (\sa_snapshot[18][23] , \sa_snapshot[18].r.part0[23] );
tran (\sa_snapshot[18][23] , \sa_snapshot[18].f.lower[23] );
tran (\sa_snapshot[18][24] , \sa_snapshot[18].r.part0[24] );
tran (\sa_snapshot[18][24] , \sa_snapshot[18].f.lower[24] );
tran (\sa_snapshot[18][25] , \sa_snapshot[18].r.part0[25] );
tran (\sa_snapshot[18][25] , \sa_snapshot[18].f.lower[25] );
tran (\sa_snapshot[18][26] , \sa_snapshot[18].r.part0[26] );
tran (\sa_snapshot[18][26] , \sa_snapshot[18].f.lower[26] );
tran (\sa_snapshot[18][27] , \sa_snapshot[18].r.part0[27] );
tran (\sa_snapshot[18][27] , \sa_snapshot[18].f.lower[27] );
tran (\sa_snapshot[18][28] , \sa_snapshot[18].r.part0[28] );
tran (\sa_snapshot[18][28] , \sa_snapshot[18].f.lower[28] );
tran (\sa_snapshot[18][29] , \sa_snapshot[18].r.part0[29] );
tran (\sa_snapshot[18][29] , \sa_snapshot[18].f.lower[29] );
tran (\sa_snapshot[18][30] , \sa_snapshot[18].r.part0[30] );
tran (\sa_snapshot[18][30] , \sa_snapshot[18].f.lower[30] );
tran (\sa_snapshot[18][31] , \sa_snapshot[18].r.part0[31] );
tran (\sa_snapshot[18][31] , \sa_snapshot[18].f.lower[31] );
tran (\sa_snapshot[18][32] , \sa_snapshot[18].r.part1[0] );
tran (\sa_snapshot[18][32] , \sa_snapshot[18].f.upper[0] );
tran (\sa_snapshot[18][33] , \sa_snapshot[18].r.part1[1] );
tran (\sa_snapshot[18][33] , \sa_snapshot[18].f.upper[1] );
tran (\sa_snapshot[18][34] , \sa_snapshot[18].r.part1[2] );
tran (\sa_snapshot[18][34] , \sa_snapshot[18].f.upper[2] );
tran (\sa_snapshot[18][35] , \sa_snapshot[18].r.part1[3] );
tran (\sa_snapshot[18][35] , \sa_snapshot[18].f.upper[3] );
tran (\sa_snapshot[18][36] , \sa_snapshot[18].r.part1[4] );
tran (\sa_snapshot[18][36] , \sa_snapshot[18].f.upper[4] );
tran (\sa_snapshot[18][37] , \sa_snapshot[18].r.part1[5] );
tran (\sa_snapshot[18][37] , \sa_snapshot[18].f.upper[5] );
tran (\sa_snapshot[18][38] , \sa_snapshot[18].r.part1[6] );
tran (\sa_snapshot[18][38] , \sa_snapshot[18].f.upper[6] );
tran (\sa_snapshot[18][39] , \sa_snapshot[18].r.part1[7] );
tran (\sa_snapshot[18][39] , \sa_snapshot[18].f.upper[7] );
tran (\sa_snapshot[18][40] , \sa_snapshot[18].r.part1[8] );
tran (\sa_snapshot[18][40] , \sa_snapshot[18].f.upper[8] );
tran (\sa_snapshot[18][41] , \sa_snapshot[18].r.part1[9] );
tran (\sa_snapshot[18][41] , \sa_snapshot[18].f.upper[9] );
tran (\sa_snapshot[18][42] , \sa_snapshot[18].r.part1[10] );
tran (\sa_snapshot[18][42] , \sa_snapshot[18].f.upper[10] );
tran (\sa_snapshot[18][43] , \sa_snapshot[18].r.part1[11] );
tran (\sa_snapshot[18][43] , \sa_snapshot[18].f.upper[11] );
tran (\sa_snapshot[18][44] , \sa_snapshot[18].r.part1[12] );
tran (\sa_snapshot[18][44] , \sa_snapshot[18].f.upper[12] );
tran (\sa_snapshot[18][45] , \sa_snapshot[18].r.part1[13] );
tran (\sa_snapshot[18][45] , \sa_snapshot[18].f.upper[13] );
tran (\sa_snapshot[18][46] , \sa_snapshot[18].r.part1[14] );
tran (\sa_snapshot[18][46] , \sa_snapshot[18].f.upper[14] );
tran (\sa_snapshot[18][47] , \sa_snapshot[18].r.part1[15] );
tran (\sa_snapshot[18][47] , \sa_snapshot[18].f.upper[15] );
tran (\sa_snapshot[18][48] , \sa_snapshot[18].r.part1[16] );
tran (\sa_snapshot[18][48] , \sa_snapshot[18].f.upper[16] );
tran (\sa_snapshot[18][49] , \sa_snapshot[18].r.part1[17] );
tran (\sa_snapshot[18][49] , \sa_snapshot[18].f.upper[17] );
tran (\sa_snapshot[18][50] , \sa_snapshot[18].r.part1[18] );
tran (\sa_snapshot[18][50] , \sa_snapshot[18].f.unused[0] );
tran (\sa_snapshot[18][51] , \sa_snapshot[18].r.part1[19] );
tran (\sa_snapshot[18][51] , \sa_snapshot[18].f.unused[1] );
tran (\sa_snapshot[18][52] , \sa_snapshot[18].r.part1[20] );
tran (\sa_snapshot[18][52] , \sa_snapshot[18].f.unused[2] );
tran (\sa_snapshot[18][53] , \sa_snapshot[18].r.part1[21] );
tran (\sa_snapshot[18][53] , \sa_snapshot[18].f.unused[3] );
tran (\sa_snapshot[18][54] , \sa_snapshot[18].r.part1[22] );
tran (\sa_snapshot[18][54] , \sa_snapshot[18].f.unused[4] );
tran (\sa_snapshot[18][55] , \sa_snapshot[18].r.part1[23] );
tran (\sa_snapshot[18][55] , \sa_snapshot[18].f.unused[5] );
tran (\sa_snapshot[18][56] , \sa_snapshot[18].r.part1[24] );
tran (\sa_snapshot[18][56] , \sa_snapshot[18].f.unused[6] );
tran (\sa_snapshot[18][57] , \sa_snapshot[18].r.part1[25] );
tran (\sa_snapshot[18][57] , \sa_snapshot[18].f.unused[7] );
tran (\sa_snapshot[18][58] , \sa_snapshot[18].r.part1[26] );
tran (\sa_snapshot[18][58] , \sa_snapshot[18].f.unused[8] );
tran (\sa_snapshot[18][59] , \sa_snapshot[18].r.part1[27] );
tran (\sa_snapshot[18][59] , \sa_snapshot[18].f.unused[9] );
tran (\sa_snapshot[18][60] , \sa_snapshot[18].r.part1[28] );
tran (\sa_snapshot[18][60] , \sa_snapshot[18].f.unused[10] );
tran (\sa_snapshot[18][61] , \sa_snapshot[18].r.part1[29] );
tran (\sa_snapshot[18][61] , \sa_snapshot[18].f.unused[11] );
tran (\sa_snapshot[18][62] , \sa_snapshot[18].r.part1[30] );
tran (\sa_snapshot[18][62] , \sa_snapshot[18].f.unused[12] );
tran (\sa_snapshot[18][63] , \sa_snapshot[18].r.part1[31] );
tran (\sa_snapshot[18][63] , \sa_snapshot[18].f.unused[13] );
tran (\sa_snapshot[19][0] , \sa_snapshot[19].r.part0[0] );
tran (\sa_snapshot[19][0] , \sa_snapshot[19].f.lower[0] );
tran (\sa_snapshot[19][1] , \sa_snapshot[19].r.part0[1] );
tran (\sa_snapshot[19][1] , \sa_snapshot[19].f.lower[1] );
tran (\sa_snapshot[19][2] , \sa_snapshot[19].r.part0[2] );
tran (\sa_snapshot[19][2] , \sa_snapshot[19].f.lower[2] );
tran (\sa_snapshot[19][3] , \sa_snapshot[19].r.part0[3] );
tran (\sa_snapshot[19][3] , \sa_snapshot[19].f.lower[3] );
tran (\sa_snapshot[19][4] , \sa_snapshot[19].r.part0[4] );
tran (\sa_snapshot[19][4] , \sa_snapshot[19].f.lower[4] );
tran (\sa_snapshot[19][5] , \sa_snapshot[19].r.part0[5] );
tran (\sa_snapshot[19][5] , \sa_snapshot[19].f.lower[5] );
tran (\sa_snapshot[19][6] , \sa_snapshot[19].r.part0[6] );
tran (\sa_snapshot[19][6] , \sa_snapshot[19].f.lower[6] );
tran (\sa_snapshot[19][7] , \sa_snapshot[19].r.part0[7] );
tran (\sa_snapshot[19][7] , \sa_snapshot[19].f.lower[7] );
tran (\sa_snapshot[19][8] , \sa_snapshot[19].r.part0[8] );
tran (\sa_snapshot[19][8] , \sa_snapshot[19].f.lower[8] );
tran (\sa_snapshot[19][9] , \sa_snapshot[19].r.part0[9] );
tran (\sa_snapshot[19][9] , \sa_snapshot[19].f.lower[9] );
tran (\sa_snapshot[19][10] , \sa_snapshot[19].r.part0[10] );
tran (\sa_snapshot[19][10] , \sa_snapshot[19].f.lower[10] );
tran (\sa_snapshot[19][11] , \sa_snapshot[19].r.part0[11] );
tran (\sa_snapshot[19][11] , \sa_snapshot[19].f.lower[11] );
tran (\sa_snapshot[19][12] , \sa_snapshot[19].r.part0[12] );
tran (\sa_snapshot[19][12] , \sa_snapshot[19].f.lower[12] );
tran (\sa_snapshot[19][13] , \sa_snapshot[19].r.part0[13] );
tran (\sa_snapshot[19][13] , \sa_snapshot[19].f.lower[13] );
tran (\sa_snapshot[19][14] , \sa_snapshot[19].r.part0[14] );
tran (\sa_snapshot[19][14] , \sa_snapshot[19].f.lower[14] );
tran (\sa_snapshot[19][15] , \sa_snapshot[19].r.part0[15] );
tran (\sa_snapshot[19][15] , \sa_snapshot[19].f.lower[15] );
tran (\sa_snapshot[19][16] , \sa_snapshot[19].r.part0[16] );
tran (\sa_snapshot[19][16] , \sa_snapshot[19].f.lower[16] );
tran (\sa_snapshot[19][17] , \sa_snapshot[19].r.part0[17] );
tran (\sa_snapshot[19][17] , \sa_snapshot[19].f.lower[17] );
tran (\sa_snapshot[19][18] , \sa_snapshot[19].r.part0[18] );
tran (\sa_snapshot[19][18] , \sa_snapshot[19].f.lower[18] );
tran (\sa_snapshot[19][19] , \sa_snapshot[19].r.part0[19] );
tran (\sa_snapshot[19][19] , \sa_snapshot[19].f.lower[19] );
tran (\sa_snapshot[19][20] , \sa_snapshot[19].r.part0[20] );
tran (\sa_snapshot[19][20] , \sa_snapshot[19].f.lower[20] );
tran (\sa_snapshot[19][21] , \sa_snapshot[19].r.part0[21] );
tran (\sa_snapshot[19][21] , \sa_snapshot[19].f.lower[21] );
tran (\sa_snapshot[19][22] , \sa_snapshot[19].r.part0[22] );
tran (\sa_snapshot[19][22] , \sa_snapshot[19].f.lower[22] );
tran (\sa_snapshot[19][23] , \sa_snapshot[19].r.part0[23] );
tran (\sa_snapshot[19][23] , \sa_snapshot[19].f.lower[23] );
tran (\sa_snapshot[19][24] , \sa_snapshot[19].r.part0[24] );
tran (\sa_snapshot[19][24] , \sa_snapshot[19].f.lower[24] );
tran (\sa_snapshot[19][25] , \sa_snapshot[19].r.part0[25] );
tran (\sa_snapshot[19][25] , \sa_snapshot[19].f.lower[25] );
tran (\sa_snapshot[19][26] , \sa_snapshot[19].r.part0[26] );
tran (\sa_snapshot[19][26] , \sa_snapshot[19].f.lower[26] );
tran (\sa_snapshot[19][27] , \sa_snapshot[19].r.part0[27] );
tran (\sa_snapshot[19][27] , \sa_snapshot[19].f.lower[27] );
tran (\sa_snapshot[19][28] , \sa_snapshot[19].r.part0[28] );
tran (\sa_snapshot[19][28] , \sa_snapshot[19].f.lower[28] );
tran (\sa_snapshot[19][29] , \sa_snapshot[19].r.part0[29] );
tran (\sa_snapshot[19][29] , \sa_snapshot[19].f.lower[29] );
tran (\sa_snapshot[19][30] , \sa_snapshot[19].r.part0[30] );
tran (\sa_snapshot[19][30] , \sa_snapshot[19].f.lower[30] );
tran (\sa_snapshot[19][31] , \sa_snapshot[19].r.part0[31] );
tran (\sa_snapshot[19][31] , \sa_snapshot[19].f.lower[31] );
tran (\sa_snapshot[19][32] , \sa_snapshot[19].r.part1[0] );
tran (\sa_snapshot[19][32] , \sa_snapshot[19].f.upper[0] );
tran (\sa_snapshot[19][33] , \sa_snapshot[19].r.part1[1] );
tran (\sa_snapshot[19][33] , \sa_snapshot[19].f.upper[1] );
tran (\sa_snapshot[19][34] , \sa_snapshot[19].r.part1[2] );
tran (\sa_snapshot[19][34] , \sa_snapshot[19].f.upper[2] );
tran (\sa_snapshot[19][35] , \sa_snapshot[19].r.part1[3] );
tran (\sa_snapshot[19][35] , \sa_snapshot[19].f.upper[3] );
tran (\sa_snapshot[19][36] , \sa_snapshot[19].r.part1[4] );
tran (\sa_snapshot[19][36] , \sa_snapshot[19].f.upper[4] );
tran (\sa_snapshot[19][37] , \sa_snapshot[19].r.part1[5] );
tran (\sa_snapshot[19][37] , \sa_snapshot[19].f.upper[5] );
tran (\sa_snapshot[19][38] , \sa_snapshot[19].r.part1[6] );
tran (\sa_snapshot[19][38] , \sa_snapshot[19].f.upper[6] );
tran (\sa_snapshot[19][39] , \sa_snapshot[19].r.part1[7] );
tran (\sa_snapshot[19][39] , \sa_snapshot[19].f.upper[7] );
tran (\sa_snapshot[19][40] , \sa_snapshot[19].r.part1[8] );
tran (\sa_snapshot[19][40] , \sa_snapshot[19].f.upper[8] );
tran (\sa_snapshot[19][41] , \sa_snapshot[19].r.part1[9] );
tran (\sa_snapshot[19][41] , \sa_snapshot[19].f.upper[9] );
tran (\sa_snapshot[19][42] , \sa_snapshot[19].r.part1[10] );
tran (\sa_snapshot[19][42] , \sa_snapshot[19].f.upper[10] );
tran (\sa_snapshot[19][43] , \sa_snapshot[19].r.part1[11] );
tran (\sa_snapshot[19][43] , \sa_snapshot[19].f.upper[11] );
tran (\sa_snapshot[19][44] , \sa_snapshot[19].r.part1[12] );
tran (\sa_snapshot[19][44] , \sa_snapshot[19].f.upper[12] );
tran (\sa_snapshot[19][45] , \sa_snapshot[19].r.part1[13] );
tran (\sa_snapshot[19][45] , \sa_snapshot[19].f.upper[13] );
tran (\sa_snapshot[19][46] , \sa_snapshot[19].r.part1[14] );
tran (\sa_snapshot[19][46] , \sa_snapshot[19].f.upper[14] );
tran (\sa_snapshot[19][47] , \sa_snapshot[19].r.part1[15] );
tran (\sa_snapshot[19][47] , \sa_snapshot[19].f.upper[15] );
tran (\sa_snapshot[19][48] , \sa_snapshot[19].r.part1[16] );
tran (\sa_snapshot[19][48] , \sa_snapshot[19].f.upper[16] );
tran (\sa_snapshot[19][49] , \sa_snapshot[19].r.part1[17] );
tran (\sa_snapshot[19][49] , \sa_snapshot[19].f.upper[17] );
tran (\sa_snapshot[19][50] , \sa_snapshot[19].r.part1[18] );
tran (\sa_snapshot[19][50] , \sa_snapshot[19].f.unused[0] );
tran (\sa_snapshot[19][51] , \sa_snapshot[19].r.part1[19] );
tran (\sa_snapshot[19][51] , \sa_snapshot[19].f.unused[1] );
tran (\sa_snapshot[19][52] , \sa_snapshot[19].r.part1[20] );
tran (\sa_snapshot[19][52] , \sa_snapshot[19].f.unused[2] );
tran (\sa_snapshot[19][53] , \sa_snapshot[19].r.part1[21] );
tran (\sa_snapshot[19][53] , \sa_snapshot[19].f.unused[3] );
tran (\sa_snapshot[19][54] , \sa_snapshot[19].r.part1[22] );
tran (\sa_snapshot[19][54] , \sa_snapshot[19].f.unused[4] );
tran (\sa_snapshot[19][55] , \sa_snapshot[19].r.part1[23] );
tran (\sa_snapshot[19][55] , \sa_snapshot[19].f.unused[5] );
tran (\sa_snapshot[19][56] , \sa_snapshot[19].r.part1[24] );
tran (\sa_snapshot[19][56] , \sa_snapshot[19].f.unused[6] );
tran (\sa_snapshot[19][57] , \sa_snapshot[19].r.part1[25] );
tran (\sa_snapshot[19][57] , \sa_snapshot[19].f.unused[7] );
tran (\sa_snapshot[19][58] , \sa_snapshot[19].r.part1[26] );
tran (\sa_snapshot[19][58] , \sa_snapshot[19].f.unused[8] );
tran (\sa_snapshot[19][59] , \sa_snapshot[19].r.part1[27] );
tran (\sa_snapshot[19][59] , \sa_snapshot[19].f.unused[9] );
tran (\sa_snapshot[19][60] , \sa_snapshot[19].r.part1[28] );
tran (\sa_snapshot[19][60] , \sa_snapshot[19].f.unused[10] );
tran (\sa_snapshot[19][61] , \sa_snapshot[19].r.part1[29] );
tran (\sa_snapshot[19][61] , \sa_snapshot[19].f.unused[11] );
tran (\sa_snapshot[19][62] , \sa_snapshot[19].r.part1[30] );
tran (\sa_snapshot[19][62] , \sa_snapshot[19].f.unused[12] );
tran (\sa_snapshot[19][63] , \sa_snapshot[19].r.part1[31] );
tran (\sa_snapshot[19][63] , \sa_snapshot[19].f.unused[13] );
tran (\sa_snapshot[20][0] , \sa_snapshot[20].r.part0[0] );
tran (\sa_snapshot[20][0] , \sa_snapshot[20].f.lower[0] );
tran (\sa_snapshot[20][1] , \sa_snapshot[20].r.part0[1] );
tran (\sa_snapshot[20][1] , \sa_snapshot[20].f.lower[1] );
tran (\sa_snapshot[20][2] , \sa_snapshot[20].r.part0[2] );
tran (\sa_snapshot[20][2] , \sa_snapshot[20].f.lower[2] );
tran (\sa_snapshot[20][3] , \sa_snapshot[20].r.part0[3] );
tran (\sa_snapshot[20][3] , \sa_snapshot[20].f.lower[3] );
tran (\sa_snapshot[20][4] , \sa_snapshot[20].r.part0[4] );
tran (\sa_snapshot[20][4] , \sa_snapshot[20].f.lower[4] );
tran (\sa_snapshot[20][5] , \sa_snapshot[20].r.part0[5] );
tran (\sa_snapshot[20][5] , \sa_snapshot[20].f.lower[5] );
tran (\sa_snapshot[20][6] , \sa_snapshot[20].r.part0[6] );
tran (\sa_snapshot[20][6] , \sa_snapshot[20].f.lower[6] );
tran (\sa_snapshot[20][7] , \sa_snapshot[20].r.part0[7] );
tran (\sa_snapshot[20][7] , \sa_snapshot[20].f.lower[7] );
tran (\sa_snapshot[20][8] , \sa_snapshot[20].r.part0[8] );
tran (\sa_snapshot[20][8] , \sa_snapshot[20].f.lower[8] );
tran (\sa_snapshot[20][9] , \sa_snapshot[20].r.part0[9] );
tran (\sa_snapshot[20][9] , \sa_snapshot[20].f.lower[9] );
tran (\sa_snapshot[20][10] , \sa_snapshot[20].r.part0[10] );
tran (\sa_snapshot[20][10] , \sa_snapshot[20].f.lower[10] );
tran (\sa_snapshot[20][11] , \sa_snapshot[20].r.part0[11] );
tran (\sa_snapshot[20][11] , \sa_snapshot[20].f.lower[11] );
tran (\sa_snapshot[20][12] , \sa_snapshot[20].r.part0[12] );
tran (\sa_snapshot[20][12] , \sa_snapshot[20].f.lower[12] );
tran (\sa_snapshot[20][13] , \sa_snapshot[20].r.part0[13] );
tran (\sa_snapshot[20][13] , \sa_snapshot[20].f.lower[13] );
tran (\sa_snapshot[20][14] , \sa_snapshot[20].r.part0[14] );
tran (\sa_snapshot[20][14] , \sa_snapshot[20].f.lower[14] );
tran (\sa_snapshot[20][15] , \sa_snapshot[20].r.part0[15] );
tran (\sa_snapshot[20][15] , \sa_snapshot[20].f.lower[15] );
tran (\sa_snapshot[20][16] , \sa_snapshot[20].r.part0[16] );
tran (\sa_snapshot[20][16] , \sa_snapshot[20].f.lower[16] );
tran (\sa_snapshot[20][17] , \sa_snapshot[20].r.part0[17] );
tran (\sa_snapshot[20][17] , \sa_snapshot[20].f.lower[17] );
tran (\sa_snapshot[20][18] , \sa_snapshot[20].r.part0[18] );
tran (\sa_snapshot[20][18] , \sa_snapshot[20].f.lower[18] );
tran (\sa_snapshot[20][19] , \sa_snapshot[20].r.part0[19] );
tran (\sa_snapshot[20][19] , \sa_snapshot[20].f.lower[19] );
tran (\sa_snapshot[20][20] , \sa_snapshot[20].r.part0[20] );
tran (\sa_snapshot[20][20] , \sa_snapshot[20].f.lower[20] );
tran (\sa_snapshot[20][21] , \sa_snapshot[20].r.part0[21] );
tran (\sa_snapshot[20][21] , \sa_snapshot[20].f.lower[21] );
tran (\sa_snapshot[20][22] , \sa_snapshot[20].r.part0[22] );
tran (\sa_snapshot[20][22] , \sa_snapshot[20].f.lower[22] );
tran (\sa_snapshot[20][23] , \sa_snapshot[20].r.part0[23] );
tran (\sa_snapshot[20][23] , \sa_snapshot[20].f.lower[23] );
tran (\sa_snapshot[20][24] , \sa_snapshot[20].r.part0[24] );
tran (\sa_snapshot[20][24] , \sa_snapshot[20].f.lower[24] );
tran (\sa_snapshot[20][25] , \sa_snapshot[20].r.part0[25] );
tran (\sa_snapshot[20][25] , \sa_snapshot[20].f.lower[25] );
tran (\sa_snapshot[20][26] , \sa_snapshot[20].r.part0[26] );
tran (\sa_snapshot[20][26] , \sa_snapshot[20].f.lower[26] );
tran (\sa_snapshot[20][27] , \sa_snapshot[20].r.part0[27] );
tran (\sa_snapshot[20][27] , \sa_snapshot[20].f.lower[27] );
tran (\sa_snapshot[20][28] , \sa_snapshot[20].r.part0[28] );
tran (\sa_snapshot[20][28] , \sa_snapshot[20].f.lower[28] );
tran (\sa_snapshot[20][29] , \sa_snapshot[20].r.part0[29] );
tran (\sa_snapshot[20][29] , \sa_snapshot[20].f.lower[29] );
tran (\sa_snapshot[20][30] , \sa_snapshot[20].r.part0[30] );
tran (\sa_snapshot[20][30] , \sa_snapshot[20].f.lower[30] );
tran (\sa_snapshot[20][31] , \sa_snapshot[20].r.part0[31] );
tran (\sa_snapshot[20][31] , \sa_snapshot[20].f.lower[31] );
tran (\sa_snapshot[20][32] , \sa_snapshot[20].r.part1[0] );
tran (\sa_snapshot[20][32] , \sa_snapshot[20].f.upper[0] );
tran (\sa_snapshot[20][33] , \sa_snapshot[20].r.part1[1] );
tran (\sa_snapshot[20][33] , \sa_snapshot[20].f.upper[1] );
tran (\sa_snapshot[20][34] , \sa_snapshot[20].r.part1[2] );
tran (\sa_snapshot[20][34] , \sa_snapshot[20].f.upper[2] );
tran (\sa_snapshot[20][35] , \sa_snapshot[20].r.part1[3] );
tran (\sa_snapshot[20][35] , \sa_snapshot[20].f.upper[3] );
tran (\sa_snapshot[20][36] , \sa_snapshot[20].r.part1[4] );
tran (\sa_snapshot[20][36] , \sa_snapshot[20].f.upper[4] );
tran (\sa_snapshot[20][37] , \sa_snapshot[20].r.part1[5] );
tran (\sa_snapshot[20][37] , \sa_snapshot[20].f.upper[5] );
tran (\sa_snapshot[20][38] , \sa_snapshot[20].r.part1[6] );
tran (\sa_snapshot[20][38] , \sa_snapshot[20].f.upper[6] );
tran (\sa_snapshot[20][39] , \sa_snapshot[20].r.part1[7] );
tran (\sa_snapshot[20][39] , \sa_snapshot[20].f.upper[7] );
tran (\sa_snapshot[20][40] , \sa_snapshot[20].r.part1[8] );
tran (\sa_snapshot[20][40] , \sa_snapshot[20].f.upper[8] );
tran (\sa_snapshot[20][41] , \sa_snapshot[20].r.part1[9] );
tran (\sa_snapshot[20][41] , \sa_snapshot[20].f.upper[9] );
tran (\sa_snapshot[20][42] , \sa_snapshot[20].r.part1[10] );
tran (\sa_snapshot[20][42] , \sa_snapshot[20].f.upper[10] );
tran (\sa_snapshot[20][43] , \sa_snapshot[20].r.part1[11] );
tran (\sa_snapshot[20][43] , \sa_snapshot[20].f.upper[11] );
tran (\sa_snapshot[20][44] , \sa_snapshot[20].r.part1[12] );
tran (\sa_snapshot[20][44] , \sa_snapshot[20].f.upper[12] );
tran (\sa_snapshot[20][45] , \sa_snapshot[20].r.part1[13] );
tran (\sa_snapshot[20][45] , \sa_snapshot[20].f.upper[13] );
tran (\sa_snapshot[20][46] , \sa_snapshot[20].r.part1[14] );
tran (\sa_snapshot[20][46] , \sa_snapshot[20].f.upper[14] );
tran (\sa_snapshot[20][47] , \sa_snapshot[20].r.part1[15] );
tran (\sa_snapshot[20][47] , \sa_snapshot[20].f.upper[15] );
tran (\sa_snapshot[20][48] , \sa_snapshot[20].r.part1[16] );
tran (\sa_snapshot[20][48] , \sa_snapshot[20].f.upper[16] );
tran (\sa_snapshot[20][49] , \sa_snapshot[20].r.part1[17] );
tran (\sa_snapshot[20][49] , \sa_snapshot[20].f.upper[17] );
tran (\sa_snapshot[20][50] , \sa_snapshot[20].r.part1[18] );
tran (\sa_snapshot[20][50] , \sa_snapshot[20].f.unused[0] );
tran (\sa_snapshot[20][51] , \sa_snapshot[20].r.part1[19] );
tran (\sa_snapshot[20][51] , \sa_snapshot[20].f.unused[1] );
tran (\sa_snapshot[20][52] , \sa_snapshot[20].r.part1[20] );
tran (\sa_snapshot[20][52] , \sa_snapshot[20].f.unused[2] );
tran (\sa_snapshot[20][53] , \sa_snapshot[20].r.part1[21] );
tran (\sa_snapshot[20][53] , \sa_snapshot[20].f.unused[3] );
tran (\sa_snapshot[20][54] , \sa_snapshot[20].r.part1[22] );
tran (\sa_snapshot[20][54] , \sa_snapshot[20].f.unused[4] );
tran (\sa_snapshot[20][55] , \sa_snapshot[20].r.part1[23] );
tran (\sa_snapshot[20][55] , \sa_snapshot[20].f.unused[5] );
tran (\sa_snapshot[20][56] , \sa_snapshot[20].r.part1[24] );
tran (\sa_snapshot[20][56] , \sa_snapshot[20].f.unused[6] );
tran (\sa_snapshot[20][57] , \sa_snapshot[20].r.part1[25] );
tran (\sa_snapshot[20][57] , \sa_snapshot[20].f.unused[7] );
tran (\sa_snapshot[20][58] , \sa_snapshot[20].r.part1[26] );
tran (\sa_snapshot[20][58] , \sa_snapshot[20].f.unused[8] );
tran (\sa_snapshot[20][59] , \sa_snapshot[20].r.part1[27] );
tran (\sa_snapshot[20][59] , \sa_snapshot[20].f.unused[9] );
tran (\sa_snapshot[20][60] , \sa_snapshot[20].r.part1[28] );
tran (\sa_snapshot[20][60] , \sa_snapshot[20].f.unused[10] );
tran (\sa_snapshot[20][61] , \sa_snapshot[20].r.part1[29] );
tran (\sa_snapshot[20][61] , \sa_snapshot[20].f.unused[11] );
tran (\sa_snapshot[20][62] , \sa_snapshot[20].r.part1[30] );
tran (\sa_snapshot[20][62] , \sa_snapshot[20].f.unused[12] );
tran (\sa_snapshot[20][63] , \sa_snapshot[20].r.part1[31] );
tran (\sa_snapshot[20][63] , \sa_snapshot[20].f.unused[13] );
tran (\sa_snapshot[21][0] , \sa_snapshot[21].r.part0[0] );
tran (\sa_snapshot[21][0] , \sa_snapshot[21].f.lower[0] );
tran (\sa_snapshot[21][1] , \sa_snapshot[21].r.part0[1] );
tran (\sa_snapshot[21][1] , \sa_snapshot[21].f.lower[1] );
tran (\sa_snapshot[21][2] , \sa_snapshot[21].r.part0[2] );
tran (\sa_snapshot[21][2] , \sa_snapshot[21].f.lower[2] );
tran (\sa_snapshot[21][3] , \sa_snapshot[21].r.part0[3] );
tran (\sa_snapshot[21][3] , \sa_snapshot[21].f.lower[3] );
tran (\sa_snapshot[21][4] , \sa_snapshot[21].r.part0[4] );
tran (\sa_snapshot[21][4] , \sa_snapshot[21].f.lower[4] );
tran (\sa_snapshot[21][5] , \sa_snapshot[21].r.part0[5] );
tran (\sa_snapshot[21][5] , \sa_snapshot[21].f.lower[5] );
tran (\sa_snapshot[21][6] , \sa_snapshot[21].r.part0[6] );
tran (\sa_snapshot[21][6] , \sa_snapshot[21].f.lower[6] );
tran (\sa_snapshot[21][7] , \sa_snapshot[21].r.part0[7] );
tran (\sa_snapshot[21][7] , \sa_snapshot[21].f.lower[7] );
tran (\sa_snapshot[21][8] , \sa_snapshot[21].r.part0[8] );
tran (\sa_snapshot[21][8] , \sa_snapshot[21].f.lower[8] );
tran (\sa_snapshot[21][9] , \sa_snapshot[21].r.part0[9] );
tran (\sa_snapshot[21][9] , \sa_snapshot[21].f.lower[9] );
tran (\sa_snapshot[21][10] , \sa_snapshot[21].r.part0[10] );
tran (\sa_snapshot[21][10] , \sa_snapshot[21].f.lower[10] );
tran (\sa_snapshot[21][11] , \sa_snapshot[21].r.part0[11] );
tran (\sa_snapshot[21][11] , \sa_snapshot[21].f.lower[11] );
tran (\sa_snapshot[21][12] , \sa_snapshot[21].r.part0[12] );
tran (\sa_snapshot[21][12] , \sa_snapshot[21].f.lower[12] );
tran (\sa_snapshot[21][13] , \sa_snapshot[21].r.part0[13] );
tran (\sa_snapshot[21][13] , \sa_snapshot[21].f.lower[13] );
tran (\sa_snapshot[21][14] , \sa_snapshot[21].r.part0[14] );
tran (\sa_snapshot[21][14] , \sa_snapshot[21].f.lower[14] );
tran (\sa_snapshot[21][15] , \sa_snapshot[21].r.part0[15] );
tran (\sa_snapshot[21][15] , \sa_snapshot[21].f.lower[15] );
tran (\sa_snapshot[21][16] , \sa_snapshot[21].r.part0[16] );
tran (\sa_snapshot[21][16] , \sa_snapshot[21].f.lower[16] );
tran (\sa_snapshot[21][17] , \sa_snapshot[21].r.part0[17] );
tran (\sa_snapshot[21][17] , \sa_snapshot[21].f.lower[17] );
tran (\sa_snapshot[21][18] , \sa_snapshot[21].r.part0[18] );
tran (\sa_snapshot[21][18] , \sa_snapshot[21].f.lower[18] );
tran (\sa_snapshot[21][19] , \sa_snapshot[21].r.part0[19] );
tran (\sa_snapshot[21][19] , \sa_snapshot[21].f.lower[19] );
tran (\sa_snapshot[21][20] , \sa_snapshot[21].r.part0[20] );
tran (\sa_snapshot[21][20] , \sa_snapshot[21].f.lower[20] );
tran (\sa_snapshot[21][21] , \sa_snapshot[21].r.part0[21] );
tran (\sa_snapshot[21][21] , \sa_snapshot[21].f.lower[21] );
tran (\sa_snapshot[21][22] , \sa_snapshot[21].r.part0[22] );
tran (\sa_snapshot[21][22] , \sa_snapshot[21].f.lower[22] );
tran (\sa_snapshot[21][23] , \sa_snapshot[21].r.part0[23] );
tran (\sa_snapshot[21][23] , \sa_snapshot[21].f.lower[23] );
tran (\sa_snapshot[21][24] , \sa_snapshot[21].r.part0[24] );
tran (\sa_snapshot[21][24] , \sa_snapshot[21].f.lower[24] );
tran (\sa_snapshot[21][25] , \sa_snapshot[21].r.part0[25] );
tran (\sa_snapshot[21][25] , \sa_snapshot[21].f.lower[25] );
tran (\sa_snapshot[21][26] , \sa_snapshot[21].r.part0[26] );
tran (\sa_snapshot[21][26] , \sa_snapshot[21].f.lower[26] );
tran (\sa_snapshot[21][27] , \sa_snapshot[21].r.part0[27] );
tran (\sa_snapshot[21][27] , \sa_snapshot[21].f.lower[27] );
tran (\sa_snapshot[21][28] , \sa_snapshot[21].r.part0[28] );
tran (\sa_snapshot[21][28] , \sa_snapshot[21].f.lower[28] );
tran (\sa_snapshot[21][29] , \sa_snapshot[21].r.part0[29] );
tran (\sa_snapshot[21][29] , \sa_snapshot[21].f.lower[29] );
tran (\sa_snapshot[21][30] , \sa_snapshot[21].r.part0[30] );
tran (\sa_snapshot[21][30] , \sa_snapshot[21].f.lower[30] );
tran (\sa_snapshot[21][31] , \sa_snapshot[21].r.part0[31] );
tran (\sa_snapshot[21][31] , \sa_snapshot[21].f.lower[31] );
tran (\sa_snapshot[21][32] , \sa_snapshot[21].r.part1[0] );
tran (\sa_snapshot[21][32] , \sa_snapshot[21].f.upper[0] );
tran (\sa_snapshot[21][33] , \sa_snapshot[21].r.part1[1] );
tran (\sa_snapshot[21][33] , \sa_snapshot[21].f.upper[1] );
tran (\sa_snapshot[21][34] , \sa_snapshot[21].r.part1[2] );
tran (\sa_snapshot[21][34] , \sa_snapshot[21].f.upper[2] );
tran (\sa_snapshot[21][35] , \sa_snapshot[21].r.part1[3] );
tran (\sa_snapshot[21][35] , \sa_snapshot[21].f.upper[3] );
tran (\sa_snapshot[21][36] , \sa_snapshot[21].r.part1[4] );
tran (\sa_snapshot[21][36] , \sa_snapshot[21].f.upper[4] );
tran (\sa_snapshot[21][37] , \sa_snapshot[21].r.part1[5] );
tran (\sa_snapshot[21][37] , \sa_snapshot[21].f.upper[5] );
tran (\sa_snapshot[21][38] , \sa_snapshot[21].r.part1[6] );
tran (\sa_snapshot[21][38] , \sa_snapshot[21].f.upper[6] );
tran (\sa_snapshot[21][39] , \sa_snapshot[21].r.part1[7] );
tran (\sa_snapshot[21][39] , \sa_snapshot[21].f.upper[7] );
tran (\sa_snapshot[21][40] , \sa_snapshot[21].r.part1[8] );
tran (\sa_snapshot[21][40] , \sa_snapshot[21].f.upper[8] );
tran (\sa_snapshot[21][41] , \sa_snapshot[21].r.part1[9] );
tran (\sa_snapshot[21][41] , \sa_snapshot[21].f.upper[9] );
tran (\sa_snapshot[21][42] , \sa_snapshot[21].r.part1[10] );
tran (\sa_snapshot[21][42] , \sa_snapshot[21].f.upper[10] );
tran (\sa_snapshot[21][43] , \sa_snapshot[21].r.part1[11] );
tran (\sa_snapshot[21][43] , \sa_snapshot[21].f.upper[11] );
tran (\sa_snapshot[21][44] , \sa_snapshot[21].r.part1[12] );
tran (\sa_snapshot[21][44] , \sa_snapshot[21].f.upper[12] );
tran (\sa_snapshot[21][45] , \sa_snapshot[21].r.part1[13] );
tran (\sa_snapshot[21][45] , \sa_snapshot[21].f.upper[13] );
tran (\sa_snapshot[21][46] , \sa_snapshot[21].r.part1[14] );
tran (\sa_snapshot[21][46] , \sa_snapshot[21].f.upper[14] );
tran (\sa_snapshot[21][47] , \sa_snapshot[21].r.part1[15] );
tran (\sa_snapshot[21][47] , \sa_snapshot[21].f.upper[15] );
tran (\sa_snapshot[21][48] , \sa_snapshot[21].r.part1[16] );
tran (\sa_snapshot[21][48] , \sa_snapshot[21].f.upper[16] );
tran (\sa_snapshot[21][49] , \sa_snapshot[21].r.part1[17] );
tran (\sa_snapshot[21][49] , \sa_snapshot[21].f.upper[17] );
tran (\sa_snapshot[21][50] , \sa_snapshot[21].r.part1[18] );
tran (\sa_snapshot[21][50] , \sa_snapshot[21].f.unused[0] );
tran (\sa_snapshot[21][51] , \sa_snapshot[21].r.part1[19] );
tran (\sa_snapshot[21][51] , \sa_snapshot[21].f.unused[1] );
tran (\sa_snapshot[21][52] , \sa_snapshot[21].r.part1[20] );
tran (\sa_snapshot[21][52] , \sa_snapshot[21].f.unused[2] );
tran (\sa_snapshot[21][53] , \sa_snapshot[21].r.part1[21] );
tran (\sa_snapshot[21][53] , \sa_snapshot[21].f.unused[3] );
tran (\sa_snapshot[21][54] , \sa_snapshot[21].r.part1[22] );
tran (\sa_snapshot[21][54] , \sa_snapshot[21].f.unused[4] );
tran (\sa_snapshot[21][55] , \sa_snapshot[21].r.part1[23] );
tran (\sa_snapshot[21][55] , \sa_snapshot[21].f.unused[5] );
tran (\sa_snapshot[21][56] , \sa_snapshot[21].r.part1[24] );
tran (\sa_snapshot[21][56] , \sa_snapshot[21].f.unused[6] );
tran (\sa_snapshot[21][57] , \sa_snapshot[21].r.part1[25] );
tran (\sa_snapshot[21][57] , \sa_snapshot[21].f.unused[7] );
tran (\sa_snapshot[21][58] , \sa_snapshot[21].r.part1[26] );
tran (\sa_snapshot[21][58] , \sa_snapshot[21].f.unused[8] );
tran (\sa_snapshot[21][59] , \sa_snapshot[21].r.part1[27] );
tran (\sa_snapshot[21][59] , \sa_snapshot[21].f.unused[9] );
tran (\sa_snapshot[21][60] , \sa_snapshot[21].r.part1[28] );
tran (\sa_snapshot[21][60] , \sa_snapshot[21].f.unused[10] );
tran (\sa_snapshot[21][61] , \sa_snapshot[21].r.part1[29] );
tran (\sa_snapshot[21][61] , \sa_snapshot[21].f.unused[11] );
tran (\sa_snapshot[21][62] , \sa_snapshot[21].r.part1[30] );
tran (\sa_snapshot[21][62] , \sa_snapshot[21].f.unused[12] );
tran (\sa_snapshot[21][63] , \sa_snapshot[21].r.part1[31] );
tran (\sa_snapshot[21][63] , \sa_snapshot[21].f.unused[13] );
tran (\sa_snapshot[22][0] , \sa_snapshot[22].r.part0[0] );
tran (\sa_snapshot[22][0] , \sa_snapshot[22].f.lower[0] );
tran (\sa_snapshot[22][1] , \sa_snapshot[22].r.part0[1] );
tran (\sa_snapshot[22][1] , \sa_snapshot[22].f.lower[1] );
tran (\sa_snapshot[22][2] , \sa_snapshot[22].r.part0[2] );
tran (\sa_snapshot[22][2] , \sa_snapshot[22].f.lower[2] );
tran (\sa_snapshot[22][3] , \sa_snapshot[22].r.part0[3] );
tran (\sa_snapshot[22][3] , \sa_snapshot[22].f.lower[3] );
tran (\sa_snapshot[22][4] , \sa_snapshot[22].r.part0[4] );
tran (\sa_snapshot[22][4] , \sa_snapshot[22].f.lower[4] );
tran (\sa_snapshot[22][5] , \sa_snapshot[22].r.part0[5] );
tran (\sa_snapshot[22][5] , \sa_snapshot[22].f.lower[5] );
tran (\sa_snapshot[22][6] , \sa_snapshot[22].r.part0[6] );
tran (\sa_snapshot[22][6] , \sa_snapshot[22].f.lower[6] );
tran (\sa_snapshot[22][7] , \sa_snapshot[22].r.part0[7] );
tran (\sa_snapshot[22][7] , \sa_snapshot[22].f.lower[7] );
tran (\sa_snapshot[22][8] , \sa_snapshot[22].r.part0[8] );
tran (\sa_snapshot[22][8] , \sa_snapshot[22].f.lower[8] );
tran (\sa_snapshot[22][9] , \sa_snapshot[22].r.part0[9] );
tran (\sa_snapshot[22][9] , \sa_snapshot[22].f.lower[9] );
tran (\sa_snapshot[22][10] , \sa_snapshot[22].r.part0[10] );
tran (\sa_snapshot[22][10] , \sa_snapshot[22].f.lower[10] );
tran (\sa_snapshot[22][11] , \sa_snapshot[22].r.part0[11] );
tran (\sa_snapshot[22][11] , \sa_snapshot[22].f.lower[11] );
tran (\sa_snapshot[22][12] , \sa_snapshot[22].r.part0[12] );
tran (\sa_snapshot[22][12] , \sa_snapshot[22].f.lower[12] );
tran (\sa_snapshot[22][13] , \sa_snapshot[22].r.part0[13] );
tran (\sa_snapshot[22][13] , \sa_snapshot[22].f.lower[13] );
tran (\sa_snapshot[22][14] , \sa_snapshot[22].r.part0[14] );
tran (\sa_snapshot[22][14] , \sa_snapshot[22].f.lower[14] );
tran (\sa_snapshot[22][15] , \sa_snapshot[22].r.part0[15] );
tran (\sa_snapshot[22][15] , \sa_snapshot[22].f.lower[15] );
tran (\sa_snapshot[22][16] , \sa_snapshot[22].r.part0[16] );
tran (\sa_snapshot[22][16] , \sa_snapshot[22].f.lower[16] );
tran (\sa_snapshot[22][17] , \sa_snapshot[22].r.part0[17] );
tran (\sa_snapshot[22][17] , \sa_snapshot[22].f.lower[17] );
tran (\sa_snapshot[22][18] , \sa_snapshot[22].r.part0[18] );
tran (\sa_snapshot[22][18] , \sa_snapshot[22].f.lower[18] );
tran (\sa_snapshot[22][19] , \sa_snapshot[22].r.part0[19] );
tran (\sa_snapshot[22][19] , \sa_snapshot[22].f.lower[19] );
tran (\sa_snapshot[22][20] , \sa_snapshot[22].r.part0[20] );
tran (\sa_snapshot[22][20] , \sa_snapshot[22].f.lower[20] );
tran (\sa_snapshot[22][21] , \sa_snapshot[22].r.part0[21] );
tran (\sa_snapshot[22][21] , \sa_snapshot[22].f.lower[21] );
tran (\sa_snapshot[22][22] , \sa_snapshot[22].r.part0[22] );
tran (\sa_snapshot[22][22] , \sa_snapshot[22].f.lower[22] );
tran (\sa_snapshot[22][23] , \sa_snapshot[22].r.part0[23] );
tran (\sa_snapshot[22][23] , \sa_snapshot[22].f.lower[23] );
tran (\sa_snapshot[22][24] , \sa_snapshot[22].r.part0[24] );
tran (\sa_snapshot[22][24] , \sa_snapshot[22].f.lower[24] );
tran (\sa_snapshot[22][25] , \sa_snapshot[22].r.part0[25] );
tran (\sa_snapshot[22][25] , \sa_snapshot[22].f.lower[25] );
tran (\sa_snapshot[22][26] , \sa_snapshot[22].r.part0[26] );
tran (\sa_snapshot[22][26] , \sa_snapshot[22].f.lower[26] );
tran (\sa_snapshot[22][27] , \sa_snapshot[22].r.part0[27] );
tran (\sa_snapshot[22][27] , \sa_snapshot[22].f.lower[27] );
tran (\sa_snapshot[22][28] , \sa_snapshot[22].r.part0[28] );
tran (\sa_snapshot[22][28] , \sa_snapshot[22].f.lower[28] );
tran (\sa_snapshot[22][29] , \sa_snapshot[22].r.part0[29] );
tran (\sa_snapshot[22][29] , \sa_snapshot[22].f.lower[29] );
tran (\sa_snapshot[22][30] , \sa_snapshot[22].r.part0[30] );
tran (\sa_snapshot[22][30] , \sa_snapshot[22].f.lower[30] );
tran (\sa_snapshot[22][31] , \sa_snapshot[22].r.part0[31] );
tran (\sa_snapshot[22][31] , \sa_snapshot[22].f.lower[31] );
tran (\sa_snapshot[22][32] , \sa_snapshot[22].r.part1[0] );
tran (\sa_snapshot[22][32] , \sa_snapshot[22].f.upper[0] );
tran (\sa_snapshot[22][33] , \sa_snapshot[22].r.part1[1] );
tran (\sa_snapshot[22][33] , \sa_snapshot[22].f.upper[1] );
tran (\sa_snapshot[22][34] , \sa_snapshot[22].r.part1[2] );
tran (\sa_snapshot[22][34] , \sa_snapshot[22].f.upper[2] );
tran (\sa_snapshot[22][35] , \sa_snapshot[22].r.part1[3] );
tran (\sa_snapshot[22][35] , \sa_snapshot[22].f.upper[3] );
tran (\sa_snapshot[22][36] , \sa_snapshot[22].r.part1[4] );
tran (\sa_snapshot[22][36] , \sa_snapshot[22].f.upper[4] );
tran (\sa_snapshot[22][37] , \sa_snapshot[22].r.part1[5] );
tran (\sa_snapshot[22][37] , \sa_snapshot[22].f.upper[5] );
tran (\sa_snapshot[22][38] , \sa_snapshot[22].r.part1[6] );
tran (\sa_snapshot[22][38] , \sa_snapshot[22].f.upper[6] );
tran (\sa_snapshot[22][39] , \sa_snapshot[22].r.part1[7] );
tran (\sa_snapshot[22][39] , \sa_snapshot[22].f.upper[7] );
tran (\sa_snapshot[22][40] , \sa_snapshot[22].r.part1[8] );
tran (\sa_snapshot[22][40] , \sa_snapshot[22].f.upper[8] );
tran (\sa_snapshot[22][41] , \sa_snapshot[22].r.part1[9] );
tran (\sa_snapshot[22][41] , \sa_snapshot[22].f.upper[9] );
tran (\sa_snapshot[22][42] , \sa_snapshot[22].r.part1[10] );
tran (\sa_snapshot[22][42] , \sa_snapshot[22].f.upper[10] );
tran (\sa_snapshot[22][43] , \sa_snapshot[22].r.part1[11] );
tran (\sa_snapshot[22][43] , \sa_snapshot[22].f.upper[11] );
tran (\sa_snapshot[22][44] , \sa_snapshot[22].r.part1[12] );
tran (\sa_snapshot[22][44] , \sa_snapshot[22].f.upper[12] );
tran (\sa_snapshot[22][45] , \sa_snapshot[22].r.part1[13] );
tran (\sa_snapshot[22][45] , \sa_snapshot[22].f.upper[13] );
tran (\sa_snapshot[22][46] , \sa_snapshot[22].r.part1[14] );
tran (\sa_snapshot[22][46] , \sa_snapshot[22].f.upper[14] );
tran (\sa_snapshot[22][47] , \sa_snapshot[22].r.part1[15] );
tran (\sa_snapshot[22][47] , \sa_snapshot[22].f.upper[15] );
tran (\sa_snapshot[22][48] , \sa_snapshot[22].r.part1[16] );
tran (\sa_snapshot[22][48] , \sa_snapshot[22].f.upper[16] );
tran (\sa_snapshot[22][49] , \sa_snapshot[22].r.part1[17] );
tran (\sa_snapshot[22][49] , \sa_snapshot[22].f.upper[17] );
tran (\sa_snapshot[22][50] , \sa_snapshot[22].r.part1[18] );
tran (\sa_snapshot[22][50] , \sa_snapshot[22].f.unused[0] );
tran (\sa_snapshot[22][51] , \sa_snapshot[22].r.part1[19] );
tran (\sa_snapshot[22][51] , \sa_snapshot[22].f.unused[1] );
tran (\sa_snapshot[22][52] , \sa_snapshot[22].r.part1[20] );
tran (\sa_snapshot[22][52] , \sa_snapshot[22].f.unused[2] );
tran (\sa_snapshot[22][53] , \sa_snapshot[22].r.part1[21] );
tran (\sa_snapshot[22][53] , \sa_snapshot[22].f.unused[3] );
tran (\sa_snapshot[22][54] , \sa_snapshot[22].r.part1[22] );
tran (\sa_snapshot[22][54] , \sa_snapshot[22].f.unused[4] );
tran (\sa_snapshot[22][55] , \sa_snapshot[22].r.part1[23] );
tran (\sa_snapshot[22][55] , \sa_snapshot[22].f.unused[5] );
tran (\sa_snapshot[22][56] , \sa_snapshot[22].r.part1[24] );
tran (\sa_snapshot[22][56] , \sa_snapshot[22].f.unused[6] );
tran (\sa_snapshot[22][57] , \sa_snapshot[22].r.part1[25] );
tran (\sa_snapshot[22][57] , \sa_snapshot[22].f.unused[7] );
tran (\sa_snapshot[22][58] , \sa_snapshot[22].r.part1[26] );
tran (\sa_snapshot[22][58] , \sa_snapshot[22].f.unused[8] );
tran (\sa_snapshot[22][59] , \sa_snapshot[22].r.part1[27] );
tran (\sa_snapshot[22][59] , \sa_snapshot[22].f.unused[9] );
tran (\sa_snapshot[22][60] , \sa_snapshot[22].r.part1[28] );
tran (\sa_snapshot[22][60] , \sa_snapshot[22].f.unused[10] );
tran (\sa_snapshot[22][61] , \sa_snapshot[22].r.part1[29] );
tran (\sa_snapshot[22][61] , \sa_snapshot[22].f.unused[11] );
tran (\sa_snapshot[22][62] , \sa_snapshot[22].r.part1[30] );
tran (\sa_snapshot[22][62] , \sa_snapshot[22].f.unused[12] );
tran (\sa_snapshot[22][63] , \sa_snapshot[22].r.part1[31] );
tran (\sa_snapshot[22][63] , \sa_snapshot[22].f.unused[13] );
tran (\sa_snapshot[23][0] , \sa_snapshot[23].r.part0[0] );
tran (\sa_snapshot[23][0] , \sa_snapshot[23].f.lower[0] );
tran (\sa_snapshot[23][1] , \sa_snapshot[23].r.part0[1] );
tran (\sa_snapshot[23][1] , \sa_snapshot[23].f.lower[1] );
tran (\sa_snapshot[23][2] , \sa_snapshot[23].r.part0[2] );
tran (\sa_snapshot[23][2] , \sa_snapshot[23].f.lower[2] );
tran (\sa_snapshot[23][3] , \sa_snapshot[23].r.part0[3] );
tran (\sa_snapshot[23][3] , \sa_snapshot[23].f.lower[3] );
tran (\sa_snapshot[23][4] , \sa_snapshot[23].r.part0[4] );
tran (\sa_snapshot[23][4] , \sa_snapshot[23].f.lower[4] );
tran (\sa_snapshot[23][5] , \sa_snapshot[23].r.part0[5] );
tran (\sa_snapshot[23][5] , \sa_snapshot[23].f.lower[5] );
tran (\sa_snapshot[23][6] , \sa_snapshot[23].r.part0[6] );
tran (\sa_snapshot[23][6] , \sa_snapshot[23].f.lower[6] );
tran (\sa_snapshot[23][7] , \sa_snapshot[23].r.part0[7] );
tran (\sa_snapshot[23][7] , \sa_snapshot[23].f.lower[7] );
tran (\sa_snapshot[23][8] , \sa_snapshot[23].r.part0[8] );
tran (\sa_snapshot[23][8] , \sa_snapshot[23].f.lower[8] );
tran (\sa_snapshot[23][9] , \sa_snapshot[23].r.part0[9] );
tran (\sa_snapshot[23][9] , \sa_snapshot[23].f.lower[9] );
tran (\sa_snapshot[23][10] , \sa_snapshot[23].r.part0[10] );
tran (\sa_snapshot[23][10] , \sa_snapshot[23].f.lower[10] );
tran (\sa_snapshot[23][11] , \sa_snapshot[23].r.part0[11] );
tran (\sa_snapshot[23][11] , \sa_snapshot[23].f.lower[11] );
tran (\sa_snapshot[23][12] , \sa_snapshot[23].r.part0[12] );
tran (\sa_snapshot[23][12] , \sa_snapshot[23].f.lower[12] );
tran (\sa_snapshot[23][13] , \sa_snapshot[23].r.part0[13] );
tran (\sa_snapshot[23][13] , \sa_snapshot[23].f.lower[13] );
tran (\sa_snapshot[23][14] , \sa_snapshot[23].r.part0[14] );
tran (\sa_snapshot[23][14] , \sa_snapshot[23].f.lower[14] );
tran (\sa_snapshot[23][15] , \sa_snapshot[23].r.part0[15] );
tran (\sa_snapshot[23][15] , \sa_snapshot[23].f.lower[15] );
tran (\sa_snapshot[23][16] , \sa_snapshot[23].r.part0[16] );
tran (\sa_snapshot[23][16] , \sa_snapshot[23].f.lower[16] );
tran (\sa_snapshot[23][17] , \sa_snapshot[23].r.part0[17] );
tran (\sa_snapshot[23][17] , \sa_snapshot[23].f.lower[17] );
tran (\sa_snapshot[23][18] , \sa_snapshot[23].r.part0[18] );
tran (\sa_snapshot[23][18] , \sa_snapshot[23].f.lower[18] );
tran (\sa_snapshot[23][19] , \sa_snapshot[23].r.part0[19] );
tran (\sa_snapshot[23][19] , \sa_snapshot[23].f.lower[19] );
tran (\sa_snapshot[23][20] , \sa_snapshot[23].r.part0[20] );
tran (\sa_snapshot[23][20] , \sa_snapshot[23].f.lower[20] );
tran (\sa_snapshot[23][21] , \sa_snapshot[23].r.part0[21] );
tran (\sa_snapshot[23][21] , \sa_snapshot[23].f.lower[21] );
tran (\sa_snapshot[23][22] , \sa_snapshot[23].r.part0[22] );
tran (\sa_snapshot[23][22] , \sa_snapshot[23].f.lower[22] );
tran (\sa_snapshot[23][23] , \sa_snapshot[23].r.part0[23] );
tran (\sa_snapshot[23][23] , \sa_snapshot[23].f.lower[23] );
tran (\sa_snapshot[23][24] , \sa_snapshot[23].r.part0[24] );
tran (\sa_snapshot[23][24] , \sa_snapshot[23].f.lower[24] );
tran (\sa_snapshot[23][25] , \sa_snapshot[23].r.part0[25] );
tran (\sa_snapshot[23][25] , \sa_snapshot[23].f.lower[25] );
tran (\sa_snapshot[23][26] , \sa_snapshot[23].r.part0[26] );
tran (\sa_snapshot[23][26] , \sa_snapshot[23].f.lower[26] );
tran (\sa_snapshot[23][27] , \sa_snapshot[23].r.part0[27] );
tran (\sa_snapshot[23][27] , \sa_snapshot[23].f.lower[27] );
tran (\sa_snapshot[23][28] , \sa_snapshot[23].r.part0[28] );
tran (\sa_snapshot[23][28] , \sa_snapshot[23].f.lower[28] );
tran (\sa_snapshot[23][29] , \sa_snapshot[23].r.part0[29] );
tran (\sa_snapshot[23][29] , \sa_snapshot[23].f.lower[29] );
tran (\sa_snapshot[23][30] , \sa_snapshot[23].r.part0[30] );
tran (\sa_snapshot[23][30] , \sa_snapshot[23].f.lower[30] );
tran (\sa_snapshot[23][31] , \sa_snapshot[23].r.part0[31] );
tran (\sa_snapshot[23][31] , \sa_snapshot[23].f.lower[31] );
tran (\sa_snapshot[23][32] , \sa_snapshot[23].r.part1[0] );
tran (\sa_snapshot[23][32] , \sa_snapshot[23].f.upper[0] );
tran (\sa_snapshot[23][33] , \sa_snapshot[23].r.part1[1] );
tran (\sa_snapshot[23][33] , \sa_snapshot[23].f.upper[1] );
tran (\sa_snapshot[23][34] , \sa_snapshot[23].r.part1[2] );
tran (\sa_snapshot[23][34] , \sa_snapshot[23].f.upper[2] );
tran (\sa_snapshot[23][35] , \sa_snapshot[23].r.part1[3] );
tran (\sa_snapshot[23][35] , \sa_snapshot[23].f.upper[3] );
tran (\sa_snapshot[23][36] , \sa_snapshot[23].r.part1[4] );
tran (\sa_snapshot[23][36] , \sa_snapshot[23].f.upper[4] );
tran (\sa_snapshot[23][37] , \sa_snapshot[23].r.part1[5] );
tran (\sa_snapshot[23][37] , \sa_snapshot[23].f.upper[5] );
tran (\sa_snapshot[23][38] , \sa_snapshot[23].r.part1[6] );
tran (\sa_snapshot[23][38] , \sa_snapshot[23].f.upper[6] );
tran (\sa_snapshot[23][39] , \sa_snapshot[23].r.part1[7] );
tran (\sa_snapshot[23][39] , \sa_snapshot[23].f.upper[7] );
tran (\sa_snapshot[23][40] , \sa_snapshot[23].r.part1[8] );
tran (\sa_snapshot[23][40] , \sa_snapshot[23].f.upper[8] );
tran (\sa_snapshot[23][41] , \sa_snapshot[23].r.part1[9] );
tran (\sa_snapshot[23][41] , \sa_snapshot[23].f.upper[9] );
tran (\sa_snapshot[23][42] , \sa_snapshot[23].r.part1[10] );
tran (\sa_snapshot[23][42] , \sa_snapshot[23].f.upper[10] );
tran (\sa_snapshot[23][43] , \sa_snapshot[23].r.part1[11] );
tran (\sa_snapshot[23][43] , \sa_snapshot[23].f.upper[11] );
tran (\sa_snapshot[23][44] , \sa_snapshot[23].r.part1[12] );
tran (\sa_snapshot[23][44] , \sa_snapshot[23].f.upper[12] );
tran (\sa_snapshot[23][45] , \sa_snapshot[23].r.part1[13] );
tran (\sa_snapshot[23][45] , \sa_snapshot[23].f.upper[13] );
tran (\sa_snapshot[23][46] , \sa_snapshot[23].r.part1[14] );
tran (\sa_snapshot[23][46] , \sa_snapshot[23].f.upper[14] );
tran (\sa_snapshot[23][47] , \sa_snapshot[23].r.part1[15] );
tran (\sa_snapshot[23][47] , \sa_snapshot[23].f.upper[15] );
tran (\sa_snapshot[23][48] , \sa_snapshot[23].r.part1[16] );
tran (\sa_snapshot[23][48] , \sa_snapshot[23].f.upper[16] );
tran (\sa_snapshot[23][49] , \sa_snapshot[23].r.part1[17] );
tran (\sa_snapshot[23][49] , \sa_snapshot[23].f.upper[17] );
tran (\sa_snapshot[23][50] , \sa_snapshot[23].r.part1[18] );
tran (\sa_snapshot[23][50] , \sa_snapshot[23].f.unused[0] );
tran (\sa_snapshot[23][51] , \sa_snapshot[23].r.part1[19] );
tran (\sa_snapshot[23][51] , \sa_snapshot[23].f.unused[1] );
tran (\sa_snapshot[23][52] , \sa_snapshot[23].r.part1[20] );
tran (\sa_snapshot[23][52] , \sa_snapshot[23].f.unused[2] );
tran (\sa_snapshot[23][53] , \sa_snapshot[23].r.part1[21] );
tran (\sa_snapshot[23][53] , \sa_snapshot[23].f.unused[3] );
tran (\sa_snapshot[23][54] , \sa_snapshot[23].r.part1[22] );
tran (\sa_snapshot[23][54] , \sa_snapshot[23].f.unused[4] );
tran (\sa_snapshot[23][55] , \sa_snapshot[23].r.part1[23] );
tran (\sa_snapshot[23][55] , \sa_snapshot[23].f.unused[5] );
tran (\sa_snapshot[23][56] , \sa_snapshot[23].r.part1[24] );
tran (\sa_snapshot[23][56] , \sa_snapshot[23].f.unused[6] );
tran (\sa_snapshot[23][57] , \sa_snapshot[23].r.part1[25] );
tran (\sa_snapshot[23][57] , \sa_snapshot[23].f.unused[7] );
tran (\sa_snapshot[23][58] , \sa_snapshot[23].r.part1[26] );
tran (\sa_snapshot[23][58] , \sa_snapshot[23].f.unused[8] );
tran (\sa_snapshot[23][59] , \sa_snapshot[23].r.part1[27] );
tran (\sa_snapshot[23][59] , \sa_snapshot[23].f.unused[9] );
tran (\sa_snapshot[23][60] , \sa_snapshot[23].r.part1[28] );
tran (\sa_snapshot[23][60] , \sa_snapshot[23].f.unused[10] );
tran (\sa_snapshot[23][61] , \sa_snapshot[23].r.part1[29] );
tran (\sa_snapshot[23][61] , \sa_snapshot[23].f.unused[11] );
tran (\sa_snapshot[23][62] , \sa_snapshot[23].r.part1[30] );
tran (\sa_snapshot[23][62] , \sa_snapshot[23].f.unused[12] );
tran (\sa_snapshot[23][63] , \sa_snapshot[23].r.part1[31] );
tran (\sa_snapshot[23][63] , \sa_snapshot[23].f.unused[13] );
tran (\sa_snapshot[24][0] , \sa_snapshot[24].r.part0[0] );
tran (\sa_snapshot[24][0] , \sa_snapshot[24].f.lower[0] );
tran (\sa_snapshot[24][1] , \sa_snapshot[24].r.part0[1] );
tran (\sa_snapshot[24][1] , \sa_snapshot[24].f.lower[1] );
tran (\sa_snapshot[24][2] , \sa_snapshot[24].r.part0[2] );
tran (\sa_snapshot[24][2] , \sa_snapshot[24].f.lower[2] );
tran (\sa_snapshot[24][3] , \sa_snapshot[24].r.part0[3] );
tran (\sa_snapshot[24][3] , \sa_snapshot[24].f.lower[3] );
tran (\sa_snapshot[24][4] , \sa_snapshot[24].r.part0[4] );
tran (\sa_snapshot[24][4] , \sa_snapshot[24].f.lower[4] );
tran (\sa_snapshot[24][5] , \sa_snapshot[24].r.part0[5] );
tran (\sa_snapshot[24][5] , \sa_snapshot[24].f.lower[5] );
tran (\sa_snapshot[24][6] , \sa_snapshot[24].r.part0[6] );
tran (\sa_snapshot[24][6] , \sa_snapshot[24].f.lower[6] );
tran (\sa_snapshot[24][7] , \sa_snapshot[24].r.part0[7] );
tran (\sa_snapshot[24][7] , \sa_snapshot[24].f.lower[7] );
tran (\sa_snapshot[24][8] , \sa_snapshot[24].r.part0[8] );
tran (\sa_snapshot[24][8] , \sa_snapshot[24].f.lower[8] );
tran (\sa_snapshot[24][9] , \sa_snapshot[24].r.part0[9] );
tran (\sa_snapshot[24][9] , \sa_snapshot[24].f.lower[9] );
tran (\sa_snapshot[24][10] , \sa_snapshot[24].r.part0[10] );
tran (\sa_snapshot[24][10] , \sa_snapshot[24].f.lower[10] );
tran (\sa_snapshot[24][11] , \sa_snapshot[24].r.part0[11] );
tran (\sa_snapshot[24][11] , \sa_snapshot[24].f.lower[11] );
tran (\sa_snapshot[24][12] , \sa_snapshot[24].r.part0[12] );
tran (\sa_snapshot[24][12] , \sa_snapshot[24].f.lower[12] );
tran (\sa_snapshot[24][13] , \sa_snapshot[24].r.part0[13] );
tran (\sa_snapshot[24][13] , \sa_snapshot[24].f.lower[13] );
tran (\sa_snapshot[24][14] , \sa_snapshot[24].r.part0[14] );
tran (\sa_snapshot[24][14] , \sa_snapshot[24].f.lower[14] );
tran (\sa_snapshot[24][15] , \sa_snapshot[24].r.part0[15] );
tran (\sa_snapshot[24][15] , \sa_snapshot[24].f.lower[15] );
tran (\sa_snapshot[24][16] , \sa_snapshot[24].r.part0[16] );
tran (\sa_snapshot[24][16] , \sa_snapshot[24].f.lower[16] );
tran (\sa_snapshot[24][17] , \sa_snapshot[24].r.part0[17] );
tran (\sa_snapshot[24][17] , \sa_snapshot[24].f.lower[17] );
tran (\sa_snapshot[24][18] , \sa_snapshot[24].r.part0[18] );
tran (\sa_snapshot[24][18] , \sa_snapshot[24].f.lower[18] );
tran (\sa_snapshot[24][19] , \sa_snapshot[24].r.part0[19] );
tran (\sa_snapshot[24][19] , \sa_snapshot[24].f.lower[19] );
tran (\sa_snapshot[24][20] , \sa_snapshot[24].r.part0[20] );
tran (\sa_snapshot[24][20] , \sa_snapshot[24].f.lower[20] );
tran (\sa_snapshot[24][21] , \sa_snapshot[24].r.part0[21] );
tran (\sa_snapshot[24][21] , \sa_snapshot[24].f.lower[21] );
tran (\sa_snapshot[24][22] , \sa_snapshot[24].r.part0[22] );
tran (\sa_snapshot[24][22] , \sa_snapshot[24].f.lower[22] );
tran (\sa_snapshot[24][23] , \sa_snapshot[24].r.part0[23] );
tran (\sa_snapshot[24][23] , \sa_snapshot[24].f.lower[23] );
tran (\sa_snapshot[24][24] , \sa_snapshot[24].r.part0[24] );
tran (\sa_snapshot[24][24] , \sa_snapshot[24].f.lower[24] );
tran (\sa_snapshot[24][25] , \sa_snapshot[24].r.part0[25] );
tran (\sa_snapshot[24][25] , \sa_snapshot[24].f.lower[25] );
tran (\sa_snapshot[24][26] , \sa_snapshot[24].r.part0[26] );
tran (\sa_snapshot[24][26] , \sa_snapshot[24].f.lower[26] );
tran (\sa_snapshot[24][27] , \sa_snapshot[24].r.part0[27] );
tran (\sa_snapshot[24][27] , \sa_snapshot[24].f.lower[27] );
tran (\sa_snapshot[24][28] , \sa_snapshot[24].r.part0[28] );
tran (\sa_snapshot[24][28] , \sa_snapshot[24].f.lower[28] );
tran (\sa_snapshot[24][29] , \sa_snapshot[24].r.part0[29] );
tran (\sa_snapshot[24][29] , \sa_snapshot[24].f.lower[29] );
tran (\sa_snapshot[24][30] , \sa_snapshot[24].r.part0[30] );
tran (\sa_snapshot[24][30] , \sa_snapshot[24].f.lower[30] );
tran (\sa_snapshot[24][31] , \sa_snapshot[24].r.part0[31] );
tran (\sa_snapshot[24][31] , \sa_snapshot[24].f.lower[31] );
tran (\sa_snapshot[24][32] , \sa_snapshot[24].r.part1[0] );
tran (\sa_snapshot[24][32] , \sa_snapshot[24].f.upper[0] );
tran (\sa_snapshot[24][33] , \sa_snapshot[24].r.part1[1] );
tran (\sa_snapshot[24][33] , \sa_snapshot[24].f.upper[1] );
tran (\sa_snapshot[24][34] , \sa_snapshot[24].r.part1[2] );
tran (\sa_snapshot[24][34] , \sa_snapshot[24].f.upper[2] );
tran (\sa_snapshot[24][35] , \sa_snapshot[24].r.part1[3] );
tran (\sa_snapshot[24][35] , \sa_snapshot[24].f.upper[3] );
tran (\sa_snapshot[24][36] , \sa_snapshot[24].r.part1[4] );
tran (\sa_snapshot[24][36] , \sa_snapshot[24].f.upper[4] );
tran (\sa_snapshot[24][37] , \sa_snapshot[24].r.part1[5] );
tran (\sa_snapshot[24][37] , \sa_snapshot[24].f.upper[5] );
tran (\sa_snapshot[24][38] , \sa_snapshot[24].r.part1[6] );
tran (\sa_snapshot[24][38] , \sa_snapshot[24].f.upper[6] );
tran (\sa_snapshot[24][39] , \sa_snapshot[24].r.part1[7] );
tran (\sa_snapshot[24][39] , \sa_snapshot[24].f.upper[7] );
tran (\sa_snapshot[24][40] , \sa_snapshot[24].r.part1[8] );
tran (\sa_snapshot[24][40] , \sa_snapshot[24].f.upper[8] );
tran (\sa_snapshot[24][41] , \sa_snapshot[24].r.part1[9] );
tran (\sa_snapshot[24][41] , \sa_snapshot[24].f.upper[9] );
tran (\sa_snapshot[24][42] , \sa_snapshot[24].r.part1[10] );
tran (\sa_snapshot[24][42] , \sa_snapshot[24].f.upper[10] );
tran (\sa_snapshot[24][43] , \sa_snapshot[24].r.part1[11] );
tran (\sa_snapshot[24][43] , \sa_snapshot[24].f.upper[11] );
tran (\sa_snapshot[24][44] , \sa_snapshot[24].r.part1[12] );
tran (\sa_snapshot[24][44] , \sa_snapshot[24].f.upper[12] );
tran (\sa_snapshot[24][45] , \sa_snapshot[24].r.part1[13] );
tran (\sa_snapshot[24][45] , \sa_snapshot[24].f.upper[13] );
tran (\sa_snapshot[24][46] , \sa_snapshot[24].r.part1[14] );
tran (\sa_snapshot[24][46] , \sa_snapshot[24].f.upper[14] );
tran (\sa_snapshot[24][47] , \sa_snapshot[24].r.part1[15] );
tran (\sa_snapshot[24][47] , \sa_snapshot[24].f.upper[15] );
tran (\sa_snapshot[24][48] , \sa_snapshot[24].r.part1[16] );
tran (\sa_snapshot[24][48] , \sa_snapshot[24].f.upper[16] );
tran (\sa_snapshot[24][49] , \sa_snapshot[24].r.part1[17] );
tran (\sa_snapshot[24][49] , \sa_snapshot[24].f.upper[17] );
tran (\sa_snapshot[24][50] , \sa_snapshot[24].r.part1[18] );
tran (\sa_snapshot[24][50] , \sa_snapshot[24].f.unused[0] );
tran (\sa_snapshot[24][51] , \sa_snapshot[24].r.part1[19] );
tran (\sa_snapshot[24][51] , \sa_snapshot[24].f.unused[1] );
tran (\sa_snapshot[24][52] , \sa_snapshot[24].r.part1[20] );
tran (\sa_snapshot[24][52] , \sa_snapshot[24].f.unused[2] );
tran (\sa_snapshot[24][53] , \sa_snapshot[24].r.part1[21] );
tran (\sa_snapshot[24][53] , \sa_snapshot[24].f.unused[3] );
tran (\sa_snapshot[24][54] , \sa_snapshot[24].r.part1[22] );
tran (\sa_snapshot[24][54] , \sa_snapshot[24].f.unused[4] );
tran (\sa_snapshot[24][55] , \sa_snapshot[24].r.part1[23] );
tran (\sa_snapshot[24][55] , \sa_snapshot[24].f.unused[5] );
tran (\sa_snapshot[24][56] , \sa_snapshot[24].r.part1[24] );
tran (\sa_snapshot[24][56] , \sa_snapshot[24].f.unused[6] );
tran (\sa_snapshot[24][57] , \sa_snapshot[24].r.part1[25] );
tran (\sa_snapshot[24][57] , \sa_snapshot[24].f.unused[7] );
tran (\sa_snapshot[24][58] , \sa_snapshot[24].r.part1[26] );
tran (\sa_snapshot[24][58] , \sa_snapshot[24].f.unused[8] );
tran (\sa_snapshot[24][59] , \sa_snapshot[24].r.part1[27] );
tran (\sa_snapshot[24][59] , \sa_snapshot[24].f.unused[9] );
tran (\sa_snapshot[24][60] , \sa_snapshot[24].r.part1[28] );
tran (\sa_snapshot[24][60] , \sa_snapshot[24].f.unused[10] );
tran (\sa_snapshot[24][61] , \sa_snapshot[24].r.part1[29] );
tran (\sa_snapshot[24][61] , \sa_snapshot[24].f.unused[11] );
tran (\sa_snapshot[24][62] , \sa_snapshot[24].r.part1[30] );
tran (\sa_snapshot[24][62] , \sa_snapshot[24].f.unused[12] );
tran (\sa_snapshot[24][63] , \sa_snapshot[24].r.part1[31] );
tran (\sa_snapshot[24][63] , \sa_snapshot[24].f.unused[13] );
tran (\sa_snapshot[25][0] , \sa_snapshot[25].r.part0[0] );
tran (\sa_snapshot[25][0] , \sa_snapshot[25].f.lower[0] );
tran (\sa_snapshot[25][1] , \sa_snapshot[25].r.part0[1] );
tran (\sa_snapshot[25][1] , \sa_snapshot[25].f.lower[1] );
tran (\sa_snapshot[25][2] , \sa_snapshot[25].r.part0[2] );
tran (\sa_snapshot[25][2] , \sa_snapshot[25].f.lower[2] );
tran (\sa_snapshot[25][3] , \sa_snapshot[25].r.part0[3] );
tran (\sa_snapshot[25][3] , \sa_snapshot[25].f.lower[3] );
tran (\sa_snapshot[25][4] , \sa_snapshot[25].r.part0[4] );
tran (\sa_snapshot[25][4] , \sa_snapshot[25].f.lower[4] );
tran (\sa_snapshot[25][5] , \sa_snapshot[25].r.part0[5] );
tran (\sa_snapshot[25][5] , \sa_snapshot[25].f.lower[5] );
tran (\sa_snapshot[25][6] , \sa_snapshot[25].r.part0[6] );
tran (\sa_snapshot[25][6] , \sa_snapshot[25].f.lower[6] );
tran (\sa_snapshot[25][7] , \sa_snapshot[25].r.part0[7] );
tran (\sa_snapshot[25][7] , \sa_snapshot[25].f.lower[7] );
tran (\sa_snapshot[25][8] , \sa_snapshot[25].r.part0[8] );
tran (\sa_snapshot[25][8] , \sa_snapshot[25].f.lower[8] );
tran (\sa_snapshot[25][9] , \sa_snapshot[25].r.part0[9] );
tran (\sa_snapshot[25][9] , \sa_snapshot[25].f.lower[9] );
tran (\sa_snapshot[25][10] , \sa_snapshot[25].r.part0[10] );
tran (\sa_snapshot[25][10] , \sa_snapshot[25].f.lower[10] );
tran (\sa_snapshot[25][11] , \sa_snapshot[25].r.part0[11] );
tran (\sa_snapshot[25][11] , \sa_snapshot[25].f.lower[11] );
tran (\sa_snapshot[25][12] , \sa_snapshot[25].r.part0[12] );
tran (\sa_snapshot[25][12] , \sa_snapshot[25].f.lower[12] );
tran (\sa_snapshot[25][13] , \sa_snapshot[25].r.part0[13] );
tran (\sa_snapshot[25][13] , \sa_snapshot[25].f.lower[13] );
tran (\sa_snapshot[25][14] , \sa_snapshot[25].r.part0[14] );
tran (\sa_snapshot[25][14] , \sa_snapshot[25].f.lower[14] );
tran (\sa_snapshot[25][15] , \sa_snapshot[25].r.part0[15] );
tran (\sa_snapshot[25][15] , \sa_snapshot[25].f.lower[15] );
tran (\sa_snapshot[25][16] , \sa_snapshot[25].r.part0[16] );
tran (\sa_snapshot[25][16] , \sa_snapshot[25].f.lower[16] );
tran (\sa_snapshot[25][17] , \sa_snapshot[25].r.part0[17] );
tran (\sa_snapshot[25][17] , \sa_snapshot[25].f.lower[17] );
tran (\sa_snapshot[25][18] , \sa_snapshot[25].r.part0[18] );
tran (\sa_snapshot[25][18] , \sa_snapshot[25].f.lower[18] );
tran (\sa_snapshot[25][19] , \sa_snapshot[25].r.part0[19] );
tran (\sa_snapshot[25][19] , \sa_snapshot[25].f.lower[19] );
tran (\sa_snapshot[25][20] , \sa_snapshot[25].r.part0[20] );
tran (\sa_snapshot[25][20] , \sa_snapshot[25].f.lower[20] );
tran (\sa_snapshot[25][21] , \sa_snapshot[25].r.part0[21] );
tran (\sa_snapshot[25][21] , \sa_snapshot[25].f.lower[21] );
tran (\sa_snapshot[25][22] , \sa_snapshot[25].r.part0[22] );
tran (\sa_snapshot[25][22] , \sa_snapshot[25].f.lower[22] );
tran (\sa_snapshot[25][23] , \sa_snapshot[25].r.part0[23] );
tran (\sa_snapshot[25][23] , \sa_snapshot[25].f.lower[23] );
tran (\sa_snapshot[25][24] , \sa_snapshot[25].r.part0[24] );
tran (\sa_snapshot[25][24] , \sa_snapshot[25].f.lower[24] );
tran (\sa_snapshot[25][25] , \sa_snapshot[25].r.part0[25] );
tran (\sa_snapshot[25][25] , \sa_snapshot[25].f.lower[25] );
tran (\sa_snapshot[25][26] , \sa_snapshot[25].r.part0[26] );
tran (\sa_snapshot[25][26] , \sa_snapshot[25].f.lower[26] );
tran (\sa_snapshot[25][27] , \sa_snapshot[25].r.part0[27] );
tran (\sa_snapshot[25][27] , \sa_snapshot[25].f.lower[27] );
tran (\sa_snapshot[25][28] , \sa_snapshot[25].r.part0[28] );
tran (\sa_snapshot[25][28] , \sa_snapshot[25].f.lower[28] );
tran (\sa_snapshot[25][29] , \sa_snapshot[25].r.part0[29] );
tran (\sa_snapshot[25][29] , \sa_snapshot[25].f.lower[29] );
tran (\sa_snapshot[25][30] , \sa_snapshot[25].r.part0[30] );
tran (\sa_snapshot[25][30] , \sa_snapshot[25].f.lower[30] );
tran (\sa_snapshot[25][31] , \sa_snapshot[25].r.part0[31] );
tran (\sa_snapshot[25][31] , \sa_snapshot[25].f.lower[31] );
tran (\sa_snapshot[25][32] , \sa_snapshot[25].r.part1[0] );
tran (\sa_snapshot[25][32] , \sa_snapshot[25].f.upper[0] );
tran (\sa_snapshot[25][33] , \sa_snapshot[25].r.part1[1] );
tran (\sa_snapshot[25][33] , \sa_snapshot[25].f.upper[1] );
tran (\sa_snapshot[25][34] , \sa_snapshot[25].r.part1[2] );
tran (\sa_snapshot[25][34] , \sa_snapshot[25].f.upper[2] );
tran (\sa_snapshot[25][35] , \sa_snapshot[25].r.part1[3] );
tran (\sa_snapshot[25][35] , \sa_snapshot[25].f.upper[3] );
tran (\sa_snapshot[25][36] , \sa_snapshot[25].r.part1[4] );
tran (\sa_snapshot[25][36] , \sa_snapshot[25].f.upper[4] );
tran (\sa_snapshot[25][37] , \sa_snapshot[25].r.part1[5] );
tran (\sa_snapshot[25][37] , \sa_snapshot[25].f.upper[5] );
tran (\sa_snapshot[25][38] , \sa_snapshot[25].r.part1[6] );
tran (\sa_snapshot[25][38] , \sa_snapshot[25].f.upper[6] );
tran (\sa_snapshot[25][39] , \sa_snapshot[25].r.part1[7] );
tran (\sa_snapshot[25][39] , \sa_snapshot[25].f.upper[7] );
tran (\sa_snapshot[25][40] , \sa_snapshot[25].r.part1[8] );
tran (\sa_snapshot[25][40] , \sa_snapshot[25].f.upper[8] );
tran (\sa_snapshot[25][41] , \sa_snapshot[25].r.part1[9] );
tran (\sa_snapshot[25][41] , \sa_snapshot[25].f.upper[9] );
tran (\sa_snapshot[25][42] , \sa_snapshot[25].r.part1[10] );
tran (\sa_snapshot[25][42] , \sa_snapshot[25].f.upper[10] );
tran (\sa_snapshot[25][43] , \sa_snapshot[25].r.part1[11] );
tran (\sa_snapshot[25][43] , \sa_snapshot[25].f.upper[11] );
tran (\sa_snapshot[25][44] , \sa_snapshot[25].r.part1[12] );
tran (\sa_snapshot[25][44] , \sa_snapshot[25].f.upper[12] );
tran (\sa_snapshot[25][45] , \sa_snapshot[25].r.part1[13] );
tran (\sa_snapshot[25][45] , \sa_snapshot[25].f.upper[13] );
tran (\sa_snapshot[25][46] , \sa_snapshot[25].r.part1[14] );
tran (\sa_snapshot[25][46] , \sa_snapshot[25].f.upper[14] );
tran (\sa_snapshot[25][47] , \sa_snapshot[25].r.part1[15] );
tran (\sa_snapshot[25][47] , \sa_snapshot[25].f.upper[15] );
tran (\sa_snapshot[25][48] , \sa_snapshot[25].r.part1[16] );
tran (\sa_snapshot[25][48] , \sa_snapshot[25].f.upper[16] );
tran (\sa_snapshot[25][49] , \sa_snapshot[25].r.part1[17] );
tran (\sa_snapshot[25][49] , \sa_snapshot[25].f.upper[17] );
tran (\sa_snapshot[25][50] , \sa_snapshot[25].r.part1[18] );
tran (\sa_snapshot[25][50] , \sa_snapshot[25].f.unused[0] );
tran (\sa_snapshot[25][51] , \sa_snapshot[25].r.part1[19] );
tran (\sa_snapshot[25][51] , \sa_snapshot[25].f.unused[1] );
tran (\sa_snapshot[25][52] , \sa_snapshot[25].r.part1[20] );
tran (\sa_snapshot[25][52] , \sa_snapshot[25].f.unused[2] );
tran (\sa_snapshot[25][53] , \sa_snapshot[25].r.part1[21] );
tran (\sa_snapshot[25][53] , \sa_snapshot[25].f.unused[3] );
tran (\sa_snapshot[25][54] , \sa_snapshot[25].r.part1[22] );
tran (\sa_snapshot[25][54] , \sa_snapshot[25].f.unused[4] );
tran (\sa_snapshot[25][55] , \sa_snapshot[25].r.part1[23] );
tran (\sa_snapshot[25][55] , \sa_snapshot[25].f.unused[5] );
tran (\sa_snapshot[25][56] , \sa_snapshot[25].r.part1[24] );
tran (\sa_snapshot[25][56] , \sa_snapshot[25].f.unused[6] );
tran (\sa_snapshot[25][57] , \sa_snapshot[25].r.part1[25] );
tran (\sa_snapshot[25][57] , \sa_snapshot[25].f.unused[7] );
tran (\sa_snapshot[25][58] , \sa_snapshot[25].r.part1[26] );
tran (\sa_snapshot[25][58] , \sa_snapshot[25].f.unused[8] );
tran (\sa_snapshot[25][59] , \sa_snapshot[25].r.part1[27] );
tran (\sa_snapshot[25][59] , \sa_snapshot[25].f.unused[9] );
tran (\sa_snapshot[25][60] , \sa_snapshot[25].r.part1[28] );
tran (\sa_snapshot[25][60] , \sa_snapshot[25].f.unused[10] );
tran (\sa_snapshot[25][61] , \sa_snapshot[25].r.part1[29] );
tran (\sa_snapshot[25][61] , \sa_snapshot[25].f.unused[11] );
tran (\sa_snapshot[25][62] , \sa_snapshot[25].r.part1[30] );
tran (\sa_snapshot[25][62] , \sa_snapshot[25].f.unused[12] );
tran (\sa_snapshot[25][63] , \sa_snapshot[25].r.part1[31] );
tran (\sa_snapshot[25][63] , \sa_snapshot[25].f.unused[13] );
tran (\sa_snapshot[26][0] , \sa_snapshot[26].r.part0[0] );
tran (\sa_snapshot[26][0] , \sa_snapshot[26].f.lower[0] );
tran (\sa_snapshot[26][1] , \sa_snapshot[26].r.part0[1] );
tran (\sa_snapshot[26][1] , \sa_snapshot[26].f.lower[1] );
tran (\sa_snapshot[26][2] , \sa_snapshot[26].r.part0[2] );
tran (\sa_snapshot[26][2] , \sa_snapshot[26].f.lower[2] );
tran (\sa_snapshot[26][3] , \sa_snapshot[26].r.part0[3] );
tran (\sa_snapshot[26][3] , \sa_snapshot[26].f.lower[3] );
tran (\sa_snapshot[26][4] , \sa_snapshot[26].r.part0[4] );
tran (\sa_snapshot[26][4] , \sa_snapshot[26].f.lower[4] );
tran (\sa_snapshot[26][5] , \sa_snapshot[26].r.part0[5] );
tran (\sa_snapshot[26][5] , \sa_snapshot[26].f.lower[5] );
tran (\sa_snapshot[26][6] , \sa_snapshot[26].r.part0[6] );
tran (\sa_snapshot[26][6] , \sa_snapshot[26].f.lower[6] );
tran (\sa_snapshot[26][7] , \sa_snapshot[26].r.part0[7] );
tran (\sa_snapshot[26][7] , \sa_snapshot[26].f.lower[7] );
tran (\sa_snapshot[26][8] , \sa_snapshot[26].r.part0[8] );
tran (\sa_snapshot[26][8] , \sa_snapshot[26].f.lower[8] );
tran (\sa_snapshot[26][9] , \sa_snapshot[26].r.part0[9] );
tran (\sa_snapshot[26][9] , \sa_snapshot[26].f.lower[9] );
tran (\sa_snapshot[26][10] , \sa_snapshot[26].r.part0[10] );
tran (\sa_snapshot[26][10] , \sa_snapshot[26].f.lower[10] );
tran (\sa_snapshot[26][11] , \sa_snapshot[26].r.part0[11] );
tran (\sa_snapshot[26][11] , \sa_snapshot[26].f.lower[11] );
tran (\sa_snapshot[26][12] , \sa_snapshot[26].r.part0[12] );
tran (\sa_snapshot[26][12] , \sa_snapshot[26].f.lower[12] );
tran (\sa_snapshot[26][13] , \sa_snapshot[26].r.part0[13] );
tran (\sa_snapshot[26][13] , \sa_snapshot[26].f.lower[13] );
tran (\sa_snapshot[26][14] , \sa_snapshot[26].r.part0[14] );
tran (\sa_snapshot[26][14] , \sa_snapshot[26].f.lower[14] );
tran (\sa_snapshot[26][15] , \sa_snapshot[26].r.part0[15] );
tran (\sa_snapshot[26][15] , \sa_snapshot[26].f.lower[15] );
tran (\sa_snapshot[26][16] , \sa_snapshot[26].r.part0[16] );
tran (\sa_snapshot[26][16] , \sa_snapshot[26].f.lower[16] );
tran (\sa_snapshot[26][17] , \sa_snapshot[26].r.part0[17] );
tran (\sa_snapshot[26][17] , \sa_snapshot[26].f.lower[17] );
tran (\sa_snapshot[26][18] , \sa_snapshot[26].r.part0[18] );
tran (\sa_snapshot[26][18] , \sa_snapshot[26].f.lower[18] );
tran (\sa_snapshot[26][19] , \sa_snapshot[26].r.part0[19] );
tran (\sa_snapshot[26][19] , \sa_snapshot[26].f.lower[19] );
tran (\sa_snapshot[26][20] , \sa_snapshot[26].r.part0[20] );
tran (\sa_snapshot[26][20] , \sa_snapshot[26].f.lower[20] );
tran (\sa_snapshot[26][21] , \sa_snapshot[26].r.part0[21] );
tran (\sa_snapshot[26][21] , \sa_snapshot[26].f.lower[21] );
tran (\sa_snapshot[26][22] , \sa_snapshot[26].r.part0[22] );
tran (\sa_snapshot[26][22] , \sa_snapshot[26].f.lower[22] );
tran (\sa_snapshot[26][23] , \sa_snapshot[26].r.part0[23] );
tran (\sa_snapshot[26][23] , \sa_snapshot[26].f.lower[23] );
tran (\sa_snapshot[26][24] , \sa_snapshot[26].r.part0[24] );
tran (\sa_snapshot[26][24] , \sa_snapshot[26].f.lower[24] );
tran (\sa_snapshot[26][25] , \sa_snapshot[26].r.part0[25] );
tran (\sa_snapshot[26][25] , \sa_snapshot[26].f.lower[25] );
tran (\sa_snapshot[26][26] , \sa_snapshot[26].r.part0[26] );
tran (\sa_snapshot[26][26] , \sa_snapshot[26].f.lower[26] );
tran (\sa_snapshot[26][27] , \sa_snapshot[26].r.part0[27] );
tran (\sa_snapshot[26][27] , \sa_snapshot[26].f.lower[27] );
tran (\sa_snapshot[26][28] , \sa_snapshot[26].r.part0[28] );
tran (\sa_snapshot[26][28] , \sa_snapshot[26].f.lower[28] );
tran (\sa_snapshot[26][29] , \sa_snapshot[26].r.part0[29] );
tran (\sa_snapshot[26][29] , \sa_snapshot[26].f.lower[29] );
tran (\sa_snapshot[26][30] , \sa_snapshot[26].r.part0[30] );
tran (\sa_snapshot[26][30] , \sa_snapshot[26].f.lower[30] );
tran (\sa_snapshot[26][31] , \sa_snapshot[26].r.part0[31] );
tran (\sa_snapshot[26][31] , \sa_snapshot[26].f.lower[31] );
tran (\sa_snapshot[26][32] , \sa_snapshot[26].r.part1[0] );
tran (\sa_snapshot[26][32] , \sa_snapshot[26].f.upper[0] );
tran (\sa_snapshot[26][33] , \sa_snapshot[26].r.part1[1] );
tran (\sa_snapshot[26][33] , \sa_snapshot[26].f.upper[1] );
tran (\sa_snapshot[26][34] , \sa_snapshot[26].r.part1[2] );
tran (\sa_snapshot[26][34] , \sa_snapshot[26].f.upper[2] );
tran (\sa_snapshot[26][35] , \sa_snapshot[26].r.part1[3] );
tran (\sa_snapshot[26][35] , \sa_snapshot[26].f.upper[3] );
tran (\sa_snapshot[26][36] , \sa_snapshot[26].r.part1[4] );
tran (\sa_snapshot[26][36] , \sa_snapshot[26].f.upper[4] );
tran (\sa_snapshot[26][37] , \sa_snapshot[26].r.part1[5] );
tran (\sa_snapshot[26][37] , \sa_snapshot[26].f.upper[5] );
tran (\sa_snapshot[26][38] , \sa_snapshot[26].r.part1[6] );
tran (\sa_snapshot[26][38] , \sa_snapshot[26].f.upper[6] );
tran (\sa_snapshot[26][39] , \sa_snapshot[26].r.part1[7] );
tran (\sa_snapshot[26][39] , \sa_snapshot[26].f.upper[7] );
tran (\sa_snapshot[26][40] , \sa_snapshot[26].r.part1[8] );
tran (\sa_snapshot[26][40] , \sa_snapshot[26].f.upper[8] );
tran (\sa_snapshot[26][41] , \sa_snapshot[26].r.part1[9] );
tran (\sa_snapshot[26][41] , \sa_snapshot[26].f.upper[9] );
tran (\sa_snapshot[26][42] , \sa_snapshot[26].r.part1[10] );
tran (\sa_snapshot[26][42] , \sa_snapshot[26].f.upper[10] );
tran (\sa_snapshot[26][43] , \sa_snapshot[26].r.part1[11] );
tran (\sa_snapshot[26][43] , \sa_snapshot[26].f.upper[11] );
tran (\sa_snapshot[26][44] , \sa_snapshot[26].r.part1[12] );
tran (\sa_snapshot[26][44] , \sa_snapshot[26].f.upper[12] );
tran (\sa_snapshot[26][45] , \sa_snapshot[26].r.part1[13] );
tran (\sa_snapshot[26][45] , \sa_snapshot[26].f.upper[13] );
tran (\sa_snapshot[26][46] , \sa_snapshot[26].r.part1[14] );
tran (\sa_snapshot[26][46] , \sa_snapshot[26].f.upper[14] );
tran (\sa_snapshot[26][47] , \sa_snapshot[26].r.part1[15] );
tran (\sa_snapshot[26][47] , \sa_snapshot[26].f.upper[15] );
tran (\sa_snapshot[26][48] , \sa_snapshot[26].r.part1[16] );
tran (\sa_snapshot[26][48] , \sa_snapshot[26].f.upper[16] );
tran (\sa_snapshot[26][49] , \sa_snapshot[26].r.part1[17] );
tran (\sa_snapshot[26][49] , \sa_snapshot[26].f.upper[17] );
tran (\sa_snapshot[26][50] , \sa_snapshot[26].r.part1[18] );
tran (\sa_snapshot[26][50] , \sa_snapshot[26].f.unused[0] );
tran (\sa_snapshot[26][51] , \sa_snapshot[26].r.part1[19] );
tran (\sa_snapshot[26][51] , \sa_snapshot[26].f.unused[1] );
tran (\sa_snapshot[26][52] , \sa_snapshot[26].r.part1[20] );
tran (\sa_snapshot[26][52] , \sa_snapshot[26].f.unused[2] );
tran (\sa_snapshot[26][53] , \sa_snapshot[26].r.part1[21] );
tran (\sa_snapshot[26][53] , \sa_snapshot[26].f.unused[3] );
tran (\sa_snapshot[26][54] , \sa_snapshot[26].r.part1[22] );
tran (\sa_snapshot[26][54] , \sa_snapshot[26].f.unused[4] );
tran (\sa_snapshot[26][55] , \sa_snapshot[26].r.part1[23] );
tran (\sa_snapshot[26][55] , \sa_snapshot[26].f.unused[5] );
tran (\sa_snapshot[26][56] , \sa_snapshot[26].r.part1[24] );
tran (\sa_snapshot[26][56] , \sa_snapshot[26].f.unused[6] );
tran (\sa_snapshot[26][57] , \sa_snapshot[26].r.part1[25] );
tran (\sa_snapshot[26][57] , \sa_snapshot[26].f.unused[7] );
tran (\sa_snapshot[26][58] , \sa_snapshot[26].r.part1[26] );
tran (\sa_snapshot[26][58] , \sa_snapshot[26].f.unused[8] );
tran (\sa_snapshot[26][59] , \sa_snapshot[26].r.part1[27] );
tran (\sa_snapshot[26][59] , \sa_snapshot[26].f.unused[9] );
tran (\sa_snapshot[26][60] , \sa_snapshot[26].r.part1[28] );
tran (\sa_snapshot[26][60] , \sa_snapshot[26].f.unused[10] );
tran (\sa_snapshot[26][61] , \sa_snapshot[26].r.part1[29] );
tran (\sa_snapshot[26][61] , \sa_snapshot[26].f.unused[11] );
tran (\sa_snapshot[26][62] , \sa_snapshot[26].r.part1[30] );
tran (\sa_snapshot[26][62] , \sa_snapshot[26].f.unused[12] );
tran (\sa_snapshot[26][63] , \sa_snapshot[26].r.part1[31] );
tran (\sa_snapshot[26][63] , \sa_snapshot[26].f.unused[13] );
tran (\sa_snapshot[27][0] , \sa_snapshot[27].r.part0[0] );
tran (\sa_snapshot[27][0] , \sa_snapshot[27].f.lower[0] );
tran (\sa_snapshot[27][1] , \sa_snapshot[27].r.part0[1] );
tran (\sa_snapshot[27][1] , \sa_snapshot[27].f.lower[1] );
tran (\sa_snapshot[27][2] , \sa_snapshot[27].r.part0[2] );
tran (\sa_snapshot[27][2] , \sa_snapshot[27].f.lower[2] );
tran (\sa_snapshot[27][3] , \sa_snapshot[27].r.part0[3] );
tran (\sa_snapshot[27][3] , \sa_snapshot[27].f.lower[3] );
tran (\sa_snapshot[27][4] , \sa_snapshot[27].r.part0[4] );
tran (\sa_snapshot[27][4] , \sa_snapshot[27].f.lower[4] );
tran (\sa_snapshot[27][5] , \sa_snapshot[27].r.part0[5] );
tran (\sa_snapshot[27][5] , \sa_snapshot[27].f.lower[5] );
tran (\sa_snapshot[27][6] , \sa_snapshot[27].r.part0[6] );
tran (\sa_snapshot[27][6] , \sa_snapshot[27].f.lower[6] );
tran (\sa_snapshot[27][7] , \sa_snapshot[27].r.part0[7] );
tran (\sa_snapshot[27][7] , \sa_snapshot[27].f.lower[7] );
tran (\sa_snapshot[27][8] , \sa_snapshot[27].r.part0[8] );
tran (\sa_snapshot[27][8] , \sa_snapshot[27].f.lower[8] );
tran (\sa_snapshot[27][9] , \sa_snapshot[27].r.part0[9] );
tran (\sa_snapshot[27][9] , \sa_snapshot[27].f.lower[9] );
tran (\sa_snapshot[27][10] , \sa_snapshot[27].r.part0[10] );
tran (\sa_snapshot[27][10] , \sa_snapshot[27].f.lower[10] );
tran (\sa_snapshot[27][11] , \sa_snapshot[27].r.part0[11] );
tran (\sa_snapshot[27][11] , \sa_snapshot[27].f.lower[11] );
tran (\sa_snapshot[27][12] , \sa_snapshot[27].r.part0[12] );
tran (\sa_snapshot[27][12] , \sa_snapshot[27].f.lower[12] );
tran (\sa_snapshot[27][13] , \sa_snapshot[27].r.part0[13] );
tran (\sa_snapshot[27][13] , \sa_snapshot[27].f.lower[13] );
tran (\sa_snapshot[27][14] , \sa_snapshot[27].r.part0[14] );
tran (\sa_snapshot[27][14] , \sa_snapshot[27].f.lower[14] );
tran (\sa_snapshot[27][15] , \sa_snapshot[27].r.part0[15] );
tran (\sa_snapshot[27][15] , \sa_snapshot[27].f.lower[15] );
tran (\sa_snapshot[27][16] , \sa_snapshot[27].r.part0[16] );
tran (\sa_snapshot[27][16] , \sa_snapshot[27].f.lower[16] );
tran (\sa_snapshot[27][17] , \sa_snapshot[27].r.part0[17] );
tran (\sa_snapshot[27][17] , \sa_snapshot[27].f.lower[17] );
tran (\sa_snapshot[27][18] , \sa_snapshot[27].r.part0[18] );
tran (\sa_snapshot[27][18] , \sa_snapshot[27].f.lower[18] );
tran (\sa_snapshot[27][19] , \sa_snapshot[27].r.part0[19] );
tran (\sa_snapshot[27][19] , \sa_snapshot[27].f.lower[19] );
tran (\sa_snapshot[27][20] , \sa_snapshot[27].r.part0[20] );
tran (\sa_snapshot[27][20] , \sa_snapshot[27].f.lower[20] );
tran (\sa_snapshot[27][21] , \sa_snapshot[27].r.part0[21] );
tran (\sa_snapshot[27][21] , \sa_snapshot[27].f.lower[21] );
tran (\sa_snapshot[27][22] , \sa_snapshot[27].r.part0[22] );
tran (\sa_snapshot[27][22] , \sa_snapshot[27].f.lower[22] );
tran (\sa_snapshot[27][23] , \sa_snapshot[27].r.part0[23] );
tran (\sa_snapshot[27][23] , \sa_snapshot[27].f.lower[23] );
tran (\sa_snapshot[27][24] , \sa_snapshot[27].r.part0[24] );
tran (\sa_snapshot[27][24] , \sa_snapshot[27].f.lower[24] );
tran (\sa_snapshot[27][25] , \sa_snapshot[27].r.part0[25] );
tran (\sa_snapshot[27][25] , \sa_snapshot[27].f.lower[25] );
tran (\sa_snapshot[27][26] , \sa_snapshot[27].r.part0[26] );
tran (\sa_snapshot[27][26] , \sa_snapshot[27].f.lower[26] );
tran (\sa_snapshot[27][27] , \sa_snapshot[27].r.part0[27] );
tran (\sa_snapshot[27][27] , \sa_snapshot[27].f.lower[27] );
tran (\sa_snapshot[27][28] , \sa_snapshot[27].r.part0[28] );
tran (\sa_snapshot[27][28] , \sa_snapshot[27].f.lower[28] );
tran (\sa_snapshot[27][29] , \sa_snapshot[27].r.part0[29] );
tran (\sa_snapshot[27][29] , \sa_snapshot[27].f.lower[29] );
tran (\sa_snapshot[27][30] , \sa_snapshot[27].r.part0[30] );
tran (\sa_snapshot[27][30] , \sa_snapshot[27].f.lower[30] );
tran (\sa_snapshot[27][31] , \sa_snapshot[27].r.part0[31] );
tran (\sa_snapshot[27][31] , \sa_snapshot[27].f.lower[31] );
tran (\sa_snapshot[27][32] , \sa_snapshot[27].r.part1[0] );
tran (\sa_snapshot[27][32] , \sa_snapshot[27].f.upper[0] );
tran (\sa_snapshot[27][33] , \sa_snapshot[27].r.part1[1] );
tran (\sa_snapshot[27][33] , \sa_snapshot[27].f.upper[1] );
tran (\sa_snapshot[27][34] , \sa_snapshot[27].r.part1[2] );
tran (\sa_snapshot[27][34] , \sa_snapshot[27].f.upper[2] );
tran (\sa_snapshot[27][35] , \sa_snapshot[27].r.part1[3] );
tran (\sa_snapshot[27][35] , \sa_snapshot[27].f.upper[3] );
tran (\sa_snapshot[27][36] , \sa_snapshot[27].r.part1[4] );
tran (\sa_snapshot[27][36] , \sa_snapshot[27].f.upper[4] );
tran (\sa_snapshot[27][37] , \sa_snapshot[27].r.part1[5] );
tran (\sa_snapshot[27][37] , \sa_snapshot[27].f.upper[5] );
tran (\sa_snapshot[27][38] , \sa_snapshot[27].r.part1[6] );
tran (\sa_snapshot[27][38] , \sa_snapshot[27].f.upper[6] );
tran (\sa_snapshot[27][39] , \sa_snapshot[27].r.part1[7] );
tran (\sa_snapshot[27][39] , \sa_snapshot[27].f.upper[7] );
tran (\sa_snapshot[27][40] , \sa_snapshot[27].r.part1[8] );
tran (\sa_snapshot[27][40] , \sa_snapshot[27].f.upper[8] );
tran (\sa_snapshot[27][41] , \sa_snapshot[27].r.part1[9] );
tran (\sa_snapshot[27][41] , \sa_snapshot[27].f.upper[9] );
tran (\sa_snapshot[27][42] , \sa_snapshot[27].r.part1[10] );
tran (\sa_snapshot[27][42] , \sa_snapshot[27].f.upper[10] );
tran (\sa_snapshot[27][43] , \sa_snapshot[27].r.part1[11] );
tran (\sa_snapshot[27][43] , \sa_snapshot[27].f.upper[11] );
tran (\sa_snapshot[27][44] , \sa_snapshot[27].r.part1[12] );
tran (\sa_snapshot[27][44] , \sa_snapshot[27].f.upper[12] );
tran (\sa_snapshot[27][45] , \sa_snapshot[27].r.part1[13] );
tran (\sa_snapshot[27][45] , \sa_snapshot[27].f.upper[13] );
tran (\sa_snapshot[27][46] , \sa_snapshot[27].r.part1[14] );
tran (\sa_snapshot[27][46] , \sa_snapshot[27].f.upper[14] );
tran (\sa_snapshot[27][47] , \sa_snapshot[27].r.part1[15] );
tran (\sa_snapshot[27][47] , \sa_snapshot[27].f.upper[15] );
tran (\sa_snapshot[27][48] , \sa_snapshot[27].r.part1[16] );
tran (\sa_snapshot[27][48] , \sa_snapshot[27].f.upper[16] );
tran (\sa_snapshot[27][49] , \sa_snapshot[27].r.part1[17] );
tran (\sa_snapshot[27][49] , \sa_snapshot[27].f.upper[17] );
tran (\sa_snapshot[27][50] , \sa_snapshot[27].r.part1[18] );
tran (\sa_snapshot[27][50] , \sa_snapshot[27].f.unused[0] );
tran (\sa_snapshot[27][51] , \sa_snapshot[27].r.part1[19] );
tran (\sa_snapshot[27][51] , \sa_snapshot[27].f.unused[1] );
tran (\sa_snapshot[27][52] , \sa_snapshot[27].r.part1[20] );
tran (\sa_snapshot[27][52] , \sa_snapshot[27].f.unused[2] );
tran (\sa_snapshot[27][53] , \sa_snapshot[27].r.part1[21] );
tran (\sa_snapshot[27][53] , \sa_snapshot[27].f.unused[3] );
tran (\sa_snapshot[27][54] , \sa_snapshot[27].r.part1[22] );
tran (\sa_snapshot[27][54] , \sa_snapshot[27].f.unused[4] );
tran (\sa_snapshot[27][55] , \sa_snapshot[27].r.part1[23] );
tran (\sa_snapshot[27][55] , \sa_snapshot[27].f.unused[5] );
tran (\sa_snapshot[27][56] , \sa_snapshot[27].r.part1[24] );
tran (\sa_snapshot[27][56] , \sa_snapshot[27].f.unused[6] );
tran (\sa_snapshot[27][57] , \sa_snapshot[27].r.part1[25] );
tran (\sa_snapshot[27][57] , \sa_snapshot[27].f.unused[7] );
tran (\sa_snapshot[27][58] , \sa_snapshot[27].r.part1[26] );
tran (\sa_snapshot[27][58] , \sa_snapshot[27].f.unused[8] );
tran (\sa_snapshot[27][59] , \sa_snapshot[27].r.part1[27] );
tran (\sa_snapshot[27][59] , \sa_snapshot[27].f.unused[9] );
tran (\sa_snapshot[27][60] , \sa_snapshot[27].r.part1[28] );
tran (\sa_snapshot[27][60] , \sa_snapshot[27].f.unused[10] );
tran (\sa_snapshot[27][61] , \sa_snapshot[27].r.part1[29] );
tran (\sa_snapshot[27][61] , \sa_snapshot[27].f.unused[11] );
tran (\sa_snapshot[27][62] , \sa_snapshot[27].r.part1[30] );
tran (\sa_snapshot[27][62] , \sa_snapshot[27].f.unused[12] );
tran (\sa_snapshot[27][63] , \sa_snapshot[27].r.part1[31] );
tran (\sa_snapshot[27][63] , \sa_snapshot[27].f.unused[13] );
tran (\sa_snapshot[28][0] , \sa_snapshot[28].r.part0[0] );
tran (\sa_snapshot[28][0] , \sa_snapshot[28].f.lower[0] );
tran (\sa_snapshot[28][1] , \sa_snapshot[28].r.part0[1] );
tran (\sa_snapshot[28][1] , \sa_snapshot[28].f.lower[1] );
tran (\sa_snapshot[28][2] , \sa_snapshot[28].r.part0[2] );
tran (\sa_snapshot[28][2] , \sa_snapshot[28].f.lower[2] );
tran (\sa_snapshot[28][3] , \sa_snapshot[28].r.part0[3] );
tran (\sa_snapshot[28][3] , \sa_snapshot[28].f.lower[3] );
tran (\sa_snapshot[28][4] , \sa_snapshot[28].r.part0[4] );
tran (\sa_snapshot[28][4] , \sa_snapshot[28].f.lower[4] );
tran (\sa_snapshot[28][5] , \sa_snapshot[28].r.part0[5] );
tran (\sa_snapshot[28][5] , \sa_snapshot[28].f.lower[5] );
tran (\sa_snapshot[28][6] , \sa_snapshot[28].r.part0[6] );
tran (\sa_snapshot[28][6] , \sa_snapshot[28].f.lower[6] );
tran (\sa_snapshot[28][7] , \sa_snapshot[28].r.part0[7] );
tran (\sa_snapshot[28][7] , \sa_snapshot[28].f.lower[7] );
tran (\sa_snapshot[28][8] , \sa_snapshot[28].r.part0[8] );
tran (\sa_snapshot[28][8] , \sa_snapshot[28].f.lower[8] );
tran (\sa_snapshot[28][9] , \sa_snapshot[28].r.part0[9] );
tran (\sa_snapshot[28][9] , \sa_snapshot[28].f.lower[9] );
tran (\sa_snapshot[28][10] , \sa_snapshot[28].r.part0[10] );
tran (\sa_snapshot[28][10] , \sa_snapshot[28].f.lower[10] );
tran (\sa_snapshot[28][11] , \sa_snapshot[28].r.part0[11] );
tran (\sa_snapshot[28][11] , \sa_snapshot[28].f.lower[11] );
tran (\sa_snapshot[28][12] , \sa_snapshot[28].r.part0[12] );
tran (\sa_snapshot[28][12] , \sa_snapshot[28].f.lower[12] );
tran (\sa_snapshot[28][13] , \sa_snapshot[28].r.part0[13] );
tran (\sa_snapshot[28][13] , \sa_snapshot[28].f.lower[13] );
tran (\sa_snapshot[28][14] , \sa_snapshot[28].r.part0[14] );
tran (\sa_snapshot[28][14] , \sa_snapshot[28].f.lower[14] );
tran (\sa_snapshot[28][15] , \sa_snapshot[28].r.part0[15] );
tran (\sa_snapshot[28][15] , \sa_snapshot[28].f.lower[15] );
tran (\sa_snapshot[28][16] , \sa_snapshot[28].r.part0[16] );
tran (\sa_snapshot[28][16] , \sa_snapshot[28].f.lower[16] );
tran (\sa_snapshot[28][17] , \sa_snapshot[28].r.part0[17] );
tran (\sa_snapshot[28][17] , \sa_snapshot[28].f.lower[17] );
tran (\sa_snapshot[28][18] , \sa_snapshot[28].r.part0[18] );
tran (\sa_snapshot[28][18] , \sa_snapshot[28].f.lower[18] );
tran (\sa_snapshot[28][19] , \sa_snapshot[28].r.part0[19] );
tran (\sa_snapshot[28][19] , \sa_snapshot[28].f.lower[19] );
tran (\sa_snapshot[28][20] , \sa_snapshot[28].r.part0[20] );
tran (\sa_snapshot[28][20] , \sa_snapshot[28].f.lower[20] );
tran (\sa_snapshot[28][21] , \sa_snapshot[28].r.part0[21] );
tran (\sa_snapshot[28][21] , \sa_snapshot[28].f.lower[21] );
tran (\sa_snapshot[28][22] , \sa_snapshot[28].r.part0[22] );
tran (\sa_snapshot[28][22] , \sa_snapshot[28].f.lower[22] );
tran (\sa_snapshot[28][23] , \sa_snapshot[28].r.part0[23] );
tran (\sa_snapshot[28][23] , \sa_snapshot[28].f.lower[23] );
tran (\sa_snapshot[28][24] , \sa_snapshot[28].r.part0[24] );
tran (\sa_snapshot[28][24] , \sa_snapshot[28].f.lower[24] );
tran (\sa_snapshot[28][25] , \sa_snapshot[28].r.part0[25] );
tran (\sa_snapshot[28][25] , \sa_snapshot[28].f.lower[25] );
tran (\sa_snapshot[28][26] , \sa_snapshot[28].r.part0[26] );
tran (\sa_snapshot[28][26] , \sa_snapshot[28].f.lower[26] );
tran (\sa_snapshot[28][27] , \sa_snapshot[28].r.part0[27] );
tran (\sa_snapshot[28][27] , \sa_snapshot[28].f.lower[27] );
tran (\sa_snapshot[28][28] , \sa_snapshot[28].r.part0[28] );
tran (\sa_snapshot[28][28] , \sa_snapshot[28].f.lower[28] );
tran (\sa_snapshot[28][29] , \sa_snapshot[28].r.part0[29] );
tran (\sa_snapshot[28][29] , \sa_snapshot[28].f.lower[29] );
tran (\sa_snapshot[28][30] , \sa_snapshot[28].r.part0[30] );
tran (\sa_snapshot[28][30] , \sa_snapshot[28].f.lower[30] );
tran (\sa_snapshot[28][31] , \sa_snapshot[28].r.part0[31] );
tran (\sa_snapshot[28][31] , \sa_snapshot[28].f.lower[31] );
tran (\sa_snapshot[28][32] , \sa_snapshot[28].r.part1[0] );
tran (\sa_snapshot[28][32] , \sa_snapshot[28].f.upper[0] );
tran (\sa_snapshot[28][33] , \sa_snapshot[28].r.part1[1] );
tran (\sa_snapshot[28][33] , \sa_snapshot[28].f.upper[1] );
tran (\sa_snapshot[28][34] , \sa_snapshot[28].r.part1[2] );
tran (\sa_snapshot[28][34] , \sa_snapshot[28].f.upper[2] );
tran (\sa_snapshot[28][35] , \sa_snapshot[28].r.part1[3] );
tran (\sa_snapshot[28][35] , \sa_snapshot[28].f.upper[3] );
tran (\sa_snapshot[28][36] , \sa_snapshot[28].r.part1[4] );
tran (\sa_snapshot[28][36] , \sa_snapshot[28].f.upper[4] );
tran (\sa_snapshot[28][37] , \sa_snapshot[28].r.part1[5] );
tran (\sa_snapshot[28][37] , \sa_snapshot[28].f.upper[5] );
tran (\sa_snapshot[28][38] , \sa_snapshot[28].r.part1[6] );
tran (\sa_snapshot[28][38] , \sa_snapshot[28].f.upper[6] );
tran (\sa_snapshot[28][39] , \sa_snapshot[28].r.part1[7] );
tran (\sa_snapshot[28][39] , \sa_snapshot[28].f.upper[7] );
tran (\sa_snapshot[28][40] , \sa_snapshot[28].r.part1[8] );
tran (\sa_snapshot[28][40] , \sa_snapshot[28].f.upper[8] );
tran (\sa_snapshot[28][41] , \sa_snapshot[28].r.part1[9] );
tran (\sa_snapshot[28][41] , \sa_snapshot[28].f.upper[9] );
tran (\sa_snapshot[28][42] , \sa_snapshot[28].r.part1[10] );
tran (\sa_snapshot[28][42] , \sa_snapshot[28].f.upper[10] );
tran (\sa_snapshot[28][43] , \sa_snapshot[28].r.part1[11] );
tran (\sa_snapshot[28][43] , \sa_snapshot[28].f.upper[11] );
tran (\sa_snapshot[28][44] , \sa_snapshot[28].r.part1[12] );
tran (\sa_snapshot[28][44] , \sa_snapshot[28].f.upper[12] );
tran (\sa_snapshot[28][45] , \sa_snapshot[28].r.part1[13] );
tran (\sa_snapshot[28][45] , \sa_snapshot[28].f.upper[13] );
tran (\sa_snapshot[28][46] , \sa_snapshot[28].r.part1[14] );
tran (\sa_snapshot[28][46] , \sa_snapshot[28].f.upper[14] );
tran (\sa_snapshot[28][47] , \sa_snapshot[28].r.part1[15] );
tran (\sa_snapshot[28][47] , \sa_snapshot[28].f.upper[15] );
tran (\sa_snapshot[28][48] , \sa_snapshot[28].r.part1[16] );
tran (\sa_snapshot[28][48] , \sa_snapshot[28].f.upper[16] );
tran (\sa_snapshot[28][49] , \sa_snapshot[28].r.part1[17] );
tran (\sa_snapshot[28][49] , \sa_snapshot[28].f.upper[17] );
tran (\sa_snapshot[28][50] , \sa_snapshot[28].r.part1[18] );
tran (\sa_snapshot[28][50] , \sa_snapshot[28].f.unused[0] );
tran (\sa_snapshot[28][51] , \sa_snapshot[28].r.part1[19] );
tran (\sa_snapshot[28][51] , \sa_snapshot[28].f.unused[1] );
tran (\sa_snapshot[28][52] , \sa_snapshot[28].r.part1[20] );
tran (\sa_snapshot[28][52] , \sa_snapshot[28].f.unused[2] );
tran (\sa_snapshot[28][53] , \sa_snapshot[28].r.part1[21] );
tran (\sa_snapshot[28][53] , \sa_snapshot[28].f.unused[3] );
tran (\sa_snapshot[28][54] , \sa_snapshot[28].r.part1[22] );
tran (\sa_snapshot[28][54] , \sa_snapshot[28].f.unused[4] );
tran (\sa_snapshot[28][55] , \sa_snapshot[28].r.part1[23] );
tran (\sa_snapshot[28][55] , \sa_snapshot[28].f.unused[5] );
tran (\sa_snapshot[28][56] , \sa_snapshot[28].r.part1[24] );
tran (\sa_snapshot[28][56] , \sa_snapshot[28].f.unused[6] );
tran (\sa_snapshot[28][57] , \sa_snapshot[28].r.part1[25] );
tran (\sa_snapshot[28][57] , \sa_snapshot[28].f.unused[7] );
tran (\sa_snapshot[28][58] , \sa_snapshot[28].r.part1[26] );
tran (\sa_snapshot[28][58] , \sa_snapshot[28].f.unused[8] );
tran (\sa_snapshot[28][59] , \sa_snapshot[28].r.part1[27] );
tran (\sa_snapshot[28][59] , \sa_snapshot[28].f.unused[9] );
tran (\sa_snapshot[28][60] , \sa_snapshot[28].r.part1[28] );
tran (\sa_snapshot[28][60] , \sa_snapshot[28].f.unused[10] );
tran (\sa_snapshot[28][61] , \sa_snapshot[28].r.part1[29] );
tran (\sa_snapshot[28][61] , \sa_snapshot[28].f.unused[11] );
tran (\sa_snapshot[28][62] , \sa_snapshot[28].r.part1[30] );
tran (\sa_snapshot[28][62] , \sa_snapshot[28].f.unused[12] );
tran (\sa_snapshot[28][63] , \sa_snapshot[28].r.part1[31] );
tran (\sa_snapshot[28][63] , \sa_snapshot[28].f.unused[13] );
tran (\sa_snapshot[29][0] , \sa_snapshot[29].r.part0[0] );
tran (\sa_snapshot[29][0] , \sa_snapshot[29].f.lower[0] );
tran (\sa_snapshot[29][1] , \sa_snapshot[29].r.part0[1] );
tran (\sa_snapshot[29][1] , \sa_snapshot[29].f.lower[1] );
tran (\sa_snapshot[29][2] , \sa_snapshot[29].r.part0[2] );
tran (\sa_snapshot[29][2] , \sa_snapshot[29].f.lower[2] );
tran (\sa_snapshot[29][3] , \sa_snapshot[29].r.part0[3] );
tran (\sa_snapshot[29][3] , \sa_snapshot[29].f.lower[3] );
tran (\sa_snapshot[29][4] , \sa_snapshot[29].r.part0[4] );
tran (\sa_snapshot[29][4] , \sa_snapshot[29].f.lower[4] );
tran (\sa_snapshot[29][5] , \sa_snapshot[29].r.part0[5] );
tran (\sa_snapshot[29][5] , \sa_snapshot[29].f.lower[5] );
tran (\sa_snapshot[29][6] , \sa_snapshot[29].r.part0[6] );
tran (\sa_snapshot[29][6] , \sa_snapshot[29].f.lower[6] );
tran (\sa_snapshot[29][7] , \sa_snapshot[29].r.part0[7] );
tran (\sa_snapshot[29][7] , \sa_snapshot[29].f.lower[7] );
tran (\sa_snapshot[29][8] , \sa_snapshot[29].r.part0[8] );
tran (\sa_snapshot[29][8] , \sa_snapshot[29].f.lower[8] );
tran (\sa_snapshot[29][9] , \sa_snapshot[29].r.part0[9] );
tran (\sa_snapshot[29][9] , \sa_snapshot[29].f.lower[9] );
tran (\sa_snapshot[29][10] , \sa_snapshot[29].r.part0[10] );
tran (\sa_snapshot[29][10] , \sa_snapshot[29].f.lower[10] );
tran (\sa_snapshot[29][11] , \sa_snapshot[29].r.part0[11] );
tran (\sa_snapshot[29][11] , \sa_snapshot[29].f.lower[11] );
tran (\sa_snapshot[29][12] , \sa_snapshot[29].r.part0[12] );
tran (\sa_snapshot[29][12] , \sa_snapshot[29].f.lower[12] );
tran (\sa_snapshot[29][13] , \sa_snapshot[29].r.part0[13] );
tran (\sa_snapshot[29][13] , \sa_snapshot[29].f.lower[13] );
tran (\sa_snapshot[29][14] , \sa_snapshot[29].r.part0[14] );
tran (\sa_snapshot[29][14] , \sa_snapshot[29].f.lower[14] );
tran (\sa_snapshot[29][15] , \sa_snapshot[29].r.part0[15] );
tran (\sa_snapshot[29][15] , \sa_snapshot[29].f.lower[15] );
tran (\sa_snapshot[29][16] , \sa_snapshot[29].r.part0[16] );
tran (\sa_snapshot[29][16] , \sa_snapshot[29].f.lower[16] );
tran (\sa_snapshot[29][17] , \sa_snapshot[29].r.part0[17] );
tran (\sa_snapshot[29][17] , \sa_snapshot[29].f.lower[17] );
tran (\sa_snapshot[29][18] , \sa_snapshot[29].r.part0[18] );
tran (\sa_snapshot[29][18] , \sa_snapshot[29].f.lower[18] );
tran (\sa_snapshot[29][19] , \sa_snapshot[29].r.part0[19] );
tran (\sa_snapshot[29][19] , \sa_snapshot[29].f.lower[19] );
tran (\sa_snapshot[29][20] , \sa_snapshot[29].r.part0[20] );
tran (\sa_snapshot[29][20] , \sa_snapshot[29].f.lower[20] );
tran (\sa_snapshot[29][21] , \sa_snapshot[29].r.part0[21] );
tran (\sa_snapshot[29][21] , \sa_snapshot[29].f.lower[21] );
tran (\sa_snapshot[29][22] , \sa_snapshot[29].r.part0[22] );
tran (\sa_snapshot[29][22] , \sa_snapshot[29].f.lower[22] );
tran (\sa_snapshot[29][23] , \sa_snapshot[29].r.part0[23] );
tran (\sa_snapshot[29][23] , \sa_snapshot[29].f.lower[23] );
tran (\sa_snapshot[29][24] , \sa_snapshot[29].r.part0[24] );
tran (\sa_snapshot[29][24] , \sa_snapshot[29].f.lower[24] );
tran (\sa_snapshot[29][25] , \sa_snapshot[29].r.part0[25] );
tran (\sa_snapshot[29][25] , \sa_snapshot[29].f.lower[25] );
tran (\sa_snapshot[29][26] , \sa_snapshot[29].r.part0[26] );
tran (\sa_snapshot[29][26] , \sa_snapshot[29].f.lower[26] );
tran (\sa_snapshot[29][27] , \sa_snapshot[29].r.part0[27] );
tran (\sa_snapshot[29][27] , \sa_snapshot[29].f.lower[27] );
tran (\sa_snapshot[29][28] , \sa_snapshot[29].r.part0[28] );
tran (\sa_snapshot[29][28] , \sa_snapshot[29].f.lower[28] );
tran (\sa_snapshot[29][29] , \sa_snapshot[29].r.part0[29] );
tran (\sa_snapshot[29][29] , \sa_snapshot[29].f.lower[29] );
tran (\sa_snapshot[29][30] , \sa_snapshot[29].r.part0[30] );
tran (\sa_snapshot[29][30] , \sa_snapshot[29].f.lower[30] );
tran (\sa_snapshot[29][31] , \sa_snapshot[29].r.part0[31] );
tran (\sa_snapshot[29][31] , \sa_snapshot[29].f.lower[31] );
tran (\sa_snapshot[29][32] , \sa_snapshot[29].r.part1[0] );
tran (\sa_snapshot[29][32] , \sa_snapshot[29].f.upper[0] );
tran (\sa_snapshot[29][33] , \sa_snapshot[29].r.part1[1] );
tran (\sa_snapshot[29][33] , \sa_snapshot[29].f.upper[1] );
tran (\sa_snapshot[29][34] , \sa_snapshot[29].r.part1[2] );
tran (\sa_snapshot[29][34] , \sa_snapshot[29].f.upper[2] );
tran (\sa_snapshot[29][35] , \sa_snapshot[29].r.part1[3] );
tran (\sa_snapshot[29][35] , \sa_snapshot[29].f.upper[3] );
tran (\sa_snapshot[29][36] , \sa_snapshot[29].r.part1[4] );
tran (\sa_snapshot[29][36] , \sa_snapshot[29].f.upper[4] );
tran (\sa_snapshot[29][37] , \sa_snapshot[29].r.part1[5] );
tran (\sa_snapshot[29][37] , \sa_snapshot[29].f.upper[5] );
tran (\sa_snapshot[29][38] , \sa_snapshot[29].r.part1[6] );
tran (\sa_snapshot[29][38] , \sa_snapshot[29].f.upper[6] );
tran (\sa_snapshot[29][39] , \sa_snapshot[29].r.part1[7] );
tran (\sa_snapshot[29][39] , \sa_snapshot[29].f.upper[7] );
tran (\sa_snapshot[29][40] , \sa_snapshot[29].r.part1[8] );
tran (\sa_snapshot[29][40] , \sa_snapshot[29].f.upper[8] );
tran (\sa_snapshot[29][41] , \sa_snapshot[29].r.part1[9] );
tran (\sa_snapshot[29][41] , \sa_snapshot[29].f.upper[9] );
tran (\sa_snapshot[29][42] , \sa_snapshot[29].r.part1[10] );
tran (\sa_snapshot[29][42] , \sa_snapshot[29].f.upper[10] );
tran (\sa_snapshot[29][43] , \sa_snapshot[29].r.part1[11] );
tran (\sa_snapshot[29][43] , \sa_snapshot[29].f.upper[11] );
tran (\sa_snapshot[29][44] , \sa_snapshot[29].r.part1[12] );
tran (\sa_snapshot[29][44] , \sa_snapshot[29].f.upper[12] );
tran (\sa_snapshot[29][45] , \sa_snapshot[29].r.part1[13] );
tran (\sa_snapshot[29][45] , \sa_snapshot[29].f.upper[13] );
tran (\sa_snapshot[29][46] , \sa_snapshot[29].r.part1[14] );
tran (\sa_snapshot[29][46] , \sa_snapshot[29].f.upper[14] );
tran (\sa_snapshot[29][47] , \sa_snapshot[29].r.part1[15] );
tran (\sa_snapshot[29][47] , \sa_snapshot[29].f.upper[15] );
tran (\sa_snapshot[29][48] , \sa_snapshot[29].r.part1[16] );
tran (\sa_snapshot[29][48] , \sa_snapshot[29].f.upper[16] );
tran (\sa_snapshot[29][49] , \sa_snapshot[29].r.part1[17] );
tran (\sa_snapshot[29][49] , \sa_snapshot[29].f.upper[17] );
tran (\sa_snapshot[29][50] , \sa_snapshot[29].r.part1[18] );
tran (\sa_snapshot[29][50] , \sa_snapshot[29].f.unused[0] );
tran (\sa_snapshot[29][51] , \sa_snapshot[29].r.part1[19] );
tran (\sa_snapshot[29][51] , \sa_snapshot[29].f.unused[1] );
tran (\sa_snapshot[29][52] , \sa_snapshot[29].r.part1[20] );
tran (\sa_snapshot[29][52] , \sa_snapshot[29].f.unused[2] );
tran (\sa_snapshot[29][53] , \sa_snapshot[29].r.part1[21] );
tran (\sa_snapshot[29][53] , \sa_snapshot[29].f.unused[3] );
tran (\sa_snapshot[29][54] , \sa_snapshot[29].r.part1[22] );
tran (\sa_snapshot[29][54] , \sa_snapshot[29].f.unused[4] );
tran (\sa_snapshot[29][55] , \sa_snapshot[29].r.part1[23] );
tran (\sa_snapshot[29][55] , \sa_snapshot[29].f.unused[5] );
tran (\sa_snapshot[29][56] , \sa_snapshot[29].r.part1[24] );
tran (\sa_snapshot[29][56] , \sa_snapshot[29].f.unused[6] );
tran (\sa_snapshot[29][57] , \sa_snapshot[29].r.part1[25] );
tran (\sa_snapshot[29][57] , \sa_snapshot[29].f.unused[7] );
tran (\sa_snapshot[29][58] , \sa_snapshot[29].r.part1[26] );
tran (\sa_snapshot[29][58] , \sa_snapshot[29].f.unused[8] );
tran (\sa_snapshot[29][59] , \sa_snapshot[29].r.part1[27] );
tran (\sa_snapshot[29][59] , \sa_snapshot[29].f.unused[9] );
tran (\sa_snapshot[29][60] , \sa_snapshot[29].r.part1[28] );
tran (\sa_snapshot[29][60] , \sa_snapshot[29].f.unused[10] );
tran (\sa_snapshot[29][61] , \sa_snapshot[29].r.part1[29] );
tran (\sa_snapshot[29][61] , \sa_snapshot[29].f.unused[11] );
tran (\sa_snapshot[29][62] , \sa_snapshot[29].r.part1[30] );
tran (\sa_snapshot[29][62] , \sa_snapshot[29].f.unused[12] );
tran (\sa_snapshot[29][63] , \sa_snapshot[29].r.part1[31] );
tran (\sa_snapshot[29][63] , \sa_snapshot[29].f.unused[13] );
tran (\sa_snapshot[30][0] , \sa_snapshot[30].r.part0[0] );
tran (\sa_snapshot[30][0] , \sa_snapshot[30].f.lower[0] );
tran (\sa_snapshot[30][1] , \sa_snapshot[30].r.part0[1] );
tran (\sa_snapshot[30][1] , \sa_snapshot[30].f.lower[1] );
tran (\sa_snapshot[30][2] , \sa_snapshot[30].r.part0[2] );
tran (\sa_snapshot[30][2] , \sa_snapshot[30].f.lower[2] );
tran (\sa_snapshot[30][3] , \sa_snapshot[30].r.part0[3] );
tran (\sa_snapshot[30][3] , \sa_snapshot[30].f.lower[3] );
tran (\sa_snapshot[30][4] , \sa_snapshot[30].r.part0[4] );
tran (\sa_snapshot[30][4] , \sa_snapshot[30].f.lower[4] );
tran (\sa_snapshot[30][5] , \sa_snapshot[30].r.part0[5] );
tran (\sa_snapshot[30][5] , \sa_snapshot[30].f.lower[5] );
tran (\sa_snapshot[30][6] , \sa_snapshot[30].r.part0[6] );
tran (\sa_snapshot[30][6] , \sa_snapshot[30].f.lower[6] );
tran (\sa_snapshot[30][7] , \sa_snapshot[30].r.part0[7] );
tran (\sa_snapshot[30][7] , \sa_snapshot[30].f.lower[7] );
tran (\sa_snapshot[30][8] , \sa_snapshot[30].r.part0[8] );
tran (\sa_snapshot[30][8] , \sa_snapshot[30].f.lower[8] );
tran (\sa_snapshot[30][9] , \sa_snapshot[30].r.part0[9] );
tran (\sa_snapshot[30][9] , \sa_snapshot[30].f.lower[9] );
tran (\sa_snapshot[30][10] , \sa_snapshot[30].r.part0[10] );
tran (\sa_snapshot[30][10] , \sa_snapshot[30].f.lower[10] );
tran (\sa_snapshot[30][11] , \sa_snapshot[30].r.part0[11] );
tran (\sa_snapshot[30][11] , \sa_snapshot[30].f.lower[11] );
tran (\sa_snapshot[30][12] , \sa_snapshot[30].r.part0[12] );
tran (\sa_snapshot[30][12] , \sa_snapshot[30].f.lower[12] );
tran (\sa_snapshot[30][13] , \sa_snapshot[30].r.part0[13] );
tran (\sa_snapshot[30][13] , \sa_snapshot[30].f.lower[13] );
tran (\sa_snapshot[30][14] , \sa_snapshot[30].r.part0[14] );
tran (\sa_snapshot[30][14] , \sa_snapshot[30].f.lower[14] );
tran (\sa_snapshot[30][15] , \sa_snapshot[30].r.part0[15] );
tran (\sa_snapshot[30][15] , \sa_snapshot[30].f.lower[15] );
tran (\sa_snapshot[30][16] , \sa_snapshot[30].r.part0[16] );
tran (\sa_snapshot[30][16] , \sa_snapshot[30].f.lower[16] );
tran (\sa_snapshot[30][17] , \sa_snapshot[30].r.part0[17] );
tran (\sa_snapshot[30][17] , \sa_snapshot[30].f.lower[17] );
tran (\sa_snapshot[30][18] , \sa_snapshot[30].r.part0[18] );
tran (\sa_snapshot[30][18] , \sa_snapshot[30].f.lower[18] );
tran (\sa_snapshot[30][19] , \sa_snapshot[30].r.part0[19] );
tran (\sa_snapshot[30][19] , \sa_snapshot[30].f.lower[19] );
tran (\sa_snapshot[30][20] , \sa_snapshot[30].r.part0[20] );
tran (\sa_snapshot[30][20] , \sa_snapshot[30].f.lower[20] );
tran (\sa_snapshot[30][21] , \sa_snapshot[30].r.part0[21] );
tran (\sa_snapshot[30][21] , \sa_snapshot[30].f.lower[21] );
tran (\sa_snapshot[30][22] , \sa_snapshot[30].r.part0[22] );
tran (\sa_snapshot[30][22] , \sa_snapshot[30].f.lower[22] );
tran (\sa_snapshot[30][23] , \sa_snapshot[30].r.part0[23] );
tran (\sa_snapshot[30][23] , \sa_snapshot[30].f.lower[23] );
tran (\sa_snapshot[30][24] , \sa_snapshot[30].r.part0[24] );
tran (\sa_snapshot[30][24] , \sa_snapshot[30].f.lower[24] );
tran (\sa_snapshot[30][25] , \sa_snapshot[30].r.part0[25] );
tran (\sa_snapshot[30][25] , \sa_snapshot[30].f.lower[25] );
tran (\sa_snapshot[30][26] , \sa_snapshot[30].r.part0[26] );
tran (\sa_snapshot[30][26] , \sa_snapshot[30].f.lower[26] );
tran (\sa_snapshot[30][27] , \sa_snapshot[30].r.part0[27] );
tran (\sa_snapshot[30][27] , \sa_snapshot[30].f.lower[27] );
tran (\sa_snapshot[30][28] , \sa_snapshot[30].r.part0[28] );
tran (\sa_snapshot[30][28] , \sa_snapshot[30].f.lower[28] );
tran (\sa_snapshot[30][29] , \sa_snapshot[30].r.part0[29] );
tran (\sa_snapshot[30][29] , \sa_snapshot[30].f.lower[29] );
tran (\sa_snapshot[30][30] , \sa_snapshot[30].r.part0[30] );
tran (\sa_snapshot[30][30] , \sa_snapshot[30].f.lower[30] );
tran (\sa_snapshot[30][31] , \sa_snapshot[30].r.part0[31] );
tran (\sa_snapshot[30][31] , \sa_snapshot[30].f.lower[31] );
tran (\sa_snapshot[30][32] , \sa_snapshot[30].r.part1[0] );
tran (\sa_snapshot[30][32] , \sa_snapshot[30].f.upper[0] );
tran (\sa_snapshot[30][33] , \sa_snapshot[30].r.part1[1] );
tran (\sa_snapshot[30][33] , \sa_snapshot[30].f.upper[1] );
tran (\sa_snapshot[30][34] , \sa_snapshot[30].r.part1[2] );
tran (\sa_snapshot[30][34] , \sa_snapshot[30].f.upper[2] );
tran (\sa_snapshot[30][35] , \sa_snapshot[30].r.part1[3] );
tran (\sa_snapshot[30][35] , \sa_snapshot[30].f.upper[3] );
tran (\sa_snapshot[30][36] , \sa_snapshot[30].r.part1[4] );
tran (\sa_snapshot[30][36] , \sa_snapshot[30].f.upper[4] );
tran (\sa_snapshot[30][37] , \sa_snapshot[30].r.part1[5] );
tran (\sa_snapshot[30][37] , \sa_snapshot[30].f.upper[5] );
tran (\sa_snapshot[30][38] , \sa_snapshot[30].r.part1[6] );
tran (\sa_snapshot[30][38] , \sa_snapshot[30].f.upper[6] );
tran (\sa_snapshot[30][39] , \sa_snapshot[30].r.part1[7] );
tran (\sa_snapshot[30][39] , \sa_snapshot[30].f.upper[7] );
tran (\sa_snapshot[30][40] , \sa_snapshot[30].r.part1[8] );
tran (\sa_snapshot[30][40] , \sa_snapshot[30].f.upper[8] );
tran (\sa_snapshot[30][41] , \sa_snapshot[30].r.part1[9] );
tran (\sa_snapshot[30][41] , \sa_snapshot[30].f.upper[9] );
tran (\sa_snapshot[30][42] , \sa_snapshot[30].r.part1[10] );
tran (\sa_snapshot[30][42] , \sa_snapshot[30].f.upper[10] );
tran (\sa_snapshot[30][43] , \sa_snapshot[30].r.part1[11] );
tran (\sa_snapshot[30][43] , \sa_snapshot[30].f.upper[11] );
tran (\sa_snapshot[30][44] , \sa_snapshot[30].r.part1[12] );
tran (\sa_snapshot[30][44] , \sa_snapshot[30].f.upper[12] );
tran (\sa_snapshot[30][45] , \sa_snapshot[30].r.part1[13] );
tran (\sa_snapshot[30][45] , \sa_snapshot[30].f.upper[13] );
tran (\sa_snapshot[30][46] , \sa_snapshot[30].r.part1[14] );
tran (\sa_snapshot[30][46] , \sa_snapshot[30].f.upper[14] );
tran (\sa_snapshot[30][47] , \sa_snapshot[30].r.part1[15] );
tran (\sa_snapshot[30][47] , \sa_snapshot[30].f.upper[15] );
tran (\sa_snapshot[30][48] , \sa_snapshot[30].r.part1[16] );
tran (\sa_snapshot[30][48] , \sa_snapshot[30].f.upper[16] );
tran (\sa_snapshot[30][49] , \sa_snapshot[30].r.part1[17] );
tran (\sa_snapshot[30][49] , \sa_snapshot[30].f.upper[17] );
tran (\sa_snapshot[30][50] , \sa_snapshot[30].r.part1[18] );
tran (\sa_snapshot[30][50] , \sa_snapshot[30].f.unused[0] );
tran (\sa_snapshot[30][51] , \sa_snapshot[30].r.part1[19] );
tran (\sa_snapshot[30][51] , \sa_snapshot[30].f.unused[1] );
tran (\sa_snapshot[30][52] , \sa_snapshot[30].r.part1[20] );
tran (\sa_snapshot[30][52] , \sa_snapshot[30].f.unused[2] );
tran (\sa_snapshot[30][53] , \sa_snapshot[30].r.part1[21] );
tran (\sa_snapshot[30][53] , \sa_snapshot[30].f.unused[3] );
tran (\sa_snapshot[30][54] , \sa_snapshot[30].r.part1[22] );
tran (\sa_snapshot[30][54] , \sa_snapshot[30].f.unused[4] );
tran (\sa_snapshot[30][55] , \sa_snapshot[30].r.part1[23] );
tran (\sa_snapshot[30][55] , \sa_snapshot[30].f.unused[5] );
tran (\sa_snapshot[30][56] , \sa_snapshot[30].r.part1[24] );
tran (\sa_snapshot[30][56] , \sa_snapshot[30].f.unused[6] );
tran (\sa_snapshot[30][57] , \sa_snapshot[30].r.part1[25] );
tran (\sa_snapshot[30][57] , \sa_snapshot[30].f.unused[7] );
tran (\sa_snapshot[30][58] , \sa_snapshot[30].r.part1[26] );
tran (\sa_snapshot[30][58] , \sa_snapshot[30].f.unused[8] );
tran (\sa_snapshot[30][59] , \sa_snapshot[30].r.part1[27] );
tran (\sa_snapshot[30][59] , \sa_snapshot[30].f.unused[9] );
tran (\sa_snapshot[30][60] , \sa_snapshot[30].r.part1[28] );
tran (\sa_snapshot[30][60] , \sa_snapshot[30].f.unused[10] );
tran (\sa_snapshot[30][61] , \sa_snapshot[30].r.part1[29] );
tran (\sa_snapshot[30][61] , \sa_snapshot[30].f.unused[11] );
tran (\sa_snapshot[30][62] , \sa_snapshot[30].r.part1[30] );
tran (\sa_snapshot[30][62] , \sa_snapshot[30].f.unused[12] );
tran (\sa_snapshot[30][63] , \sa_snapshot[30].r.part1[31] );
tran (\sa_snapshot[30][63] , \sa_snapshot[30].f.unused[13] );
tran (\sa_snapshot[31][0] , \sa_snapshot[31].r.part0[0] );
tran (\sa_snapshot[31][0] , \sa_snapshot[31].f.lower[0] );
tran (\sa_snapshot[31][1] , \sa_snapshot[31].r.part0[1] );
tran (\sa_snapshot[31][1] , \sa_snapshot[31].f.lower[1] );
tran (\sa_snapshot[31][2] , \sa_snapshot[31].r.part0[2] );
tran (\sa_snapshot[31][2] , \sa_snapshot[31].f.lower[2] );
tran (\sa_snapshot[31][3] , \sa_snapshot[31].r.part0[3] );
tran (\sa_snapshot[31][3] , \sa_snapshot[31].f.lower[3] );
tran (\sa_snapshot[31][4] , \sa_snapshot[31].r.part0[4] );
tran (\sa_snapshot[31][4] , \sa_snapshot[31].f.lower[4] );
tran (\sa_snapshot[31][5] , \sa_snapshot[31].r.part0[5] );
tran (\sa_snapshot[31][5] , \sa_snapshot[31].f.lower[5] );
tran (\sa_snapshot[31][6] , \sa_snapshot[31].r.part0[6] );
tran (\sa_snapshot[31][6] , \sa_snapshot[31].f.lower[6] );
tran (\sa_snapshot[31][7] , \sa_snapshot[31].r.part0[7] );
tran (\sa_snapshot[31][7] , \sa_snapshot[31].f.lower[7] );
tran (\sa_snapshot[31][8] , \sa_snapshot[31].r.part0[8] );
tran (\sa_snapshot[31][8] , \sa_snapshot[31].f.lower[8] );
tran (\sa_snapshot[31][9] , \sa_snapshot[31].r.part0[9] );
tran (\sa_snapshot[31][9] , \sa_snapshot[31].f.lower[9] );
tran (\sa_snapshot[31][10] , \sa_snapshot[31].r.part0[10] );
tran (\sa_snapshot[31][10] , \sa_snapshot[31].f.lower[10] );
tran (\sa_snapshot[31][11] , \sa_snapshot[31].r.part0[11] );
tran (\sa_snapshot[31][11] , \sa_snapshot[31].f.lower[11] );
tran (\sa_snapshot[31][12] , \sa_snapshot[31].r.part0[12] );
tran (\sa_snapshot[31][12] , \sa_snapshot[31].f.lower[12] );
tran (\sa_snapshot[31][13] , \sa_snapshot[31].r.part0[13] );
tran (\sa_snapshot[31][13] , \sa_snapshot[31].f.lower[13] );
tran (\sa_snapshot[31][14] , \sa_snapshot[31].r.part0[14] );
tran (\sa_snapshot[31][14] , \sa_snapshot[31].f.lower[14] );
tran (\sa_snapshot[31][15] , \sa_snapshot[31].r.part0[15] );
tran (\sa_snapshot[31][15] , \sa_snapshot[31].f.lower[15] );
tran (\sa_snapshot[31][16] , \sa_snapshot[31].r.part0[16] );
tran (\sa_snapshot[31][16] , \sa_snapshot[31].f.lower[16] );
tran (\sa_snapshot[31][17] , \sa_snapshot[31].r.part0[17] );
tran (\sa_snapshot[31][17] , \sa_snapshot[31].f.lower[17] );
tran (\sa_snapshot[31][18] , \sa_snapshot[31].r.part0[18] );
tran (\sa_snapshot[31][18] , \sa_snapshot[31].f.lower[18] );
tran (\sa_snapshot[31][19] , \sa_snapshot[31].r.part0[19] );
tran (\sa_snapshot[31][19] , \sa_snapshot[31].f.lower[19] );
tran (\sa_snapshot[31][20] , \sa_snapshot[31].r.part0[20] );
tran (\sa_snapshot[31][20] , \sa_snapshot[31].f.lower[20] );
tran (\sa_snapshot[31][21] , \sa_snapshot[31].r.part0[21] );
tran (\sa_snapshot[31][21] , \sa_snapshot[31].f.lower[21] );
tran (\sa_snapshot[31][22] , \sa_snapshot[31].r.part0[22] );
tran (\sa_snapshot[31][22] , \sa_snapshot[31].f.lower[22] );
tran (\sa_snapshot[31][23] , \sa_snapshot[31].r.part0[23] );
tran (\sa_snapshot[31][23] , \sa_snapshot[31].f.lower[23] );
tran (\sa_snapshot[31][24] , \sa_snapshot[31].r.part0[24] );
tran (\sa_snapshot[31][24] , \sa_snapshot[31].f.lower[24] );
tran (\sa_snapshot[31][25] , \sa_snapshot[31].r.part0[25] );
tran (\sa_snapshot[31][25] , \sa_snapshot[31].f.lower[25] );
tran (\sa_snapshot[31][26] , \sa_snapshot[31].r.part0[26] );
tran (\sa_snapshot[31][26] , \sa_snapshot[31].f.lower[26] );
tran (\sa_snapshot[31][27] , \sa_snapshot[31].r.part0[27] );
tran (\sa_snapshot[31][27] , \sa_snapshot[31].f.lower[27] );
tran (\sa_snapshot[31][28] , \sa_snapshot[31].r.part0[28] );
tran (\sa_snapshot[31][28] , \sa_snapshot[31].f.lower[28] );
tran (\sa_snapshot[31][29] , \sa_snapshot[31].r.part0[29] );
tran (\sa_snapshot[31][29] , \sa_snapshot[31].f.lower[29] );
tran (\sa_snapshot[31][30] , \sa_snapshot[31].r.part0[30] );
tran (\sa_snapshot[31][30] , \sa_snapshot[31].f.lower[30] );
tran (\sa_snapshot[31][31] , \sa_snapshot[31].r.part0[31] );
tran (\sa_snapshot[31][31] , \sa_snapshot[31].f.lower[31] );
tran (\sa_snapshot[31][32] , \sa_snapshot[31].r.part1[0] );
tran (\sa_snapshot[31][32] , \sa_snapshot[31].f.upper[0] );
tran (\sa_snapshot[31][33] , \sa_snapshot[31].r.part1[1] );
tran (\sa_snapshot[31][33] , \sa_snapshot[31].f.upper[1] );
tran (\sa_snapshot[31][34] , \sa_snapshot[31].r.part1[2] );
tran (\sa_snapshot[31][34] , \sa_snapshot[31].f.upper[2] );
tran (\sa_snapshot[31][35] , \sa_snapshot[31].r.part1[3] );
tran (\sa_snapshot[31][35] , \sa_snapshot[31].f.upper[3] );
tran (\sa_snapshot[31][36] , \sa_snapshot[31].r.part1[4] );
tran (\sa_snapshot[31][36] , \sa_snapshot[31].f.upper[4] );
tran (\sa_snapshot[31][37] , \sa_snapshot[31].r.part1[5] );
tran (\sa_snapshot[31][37] , \sa_snapshot[31].f.upper[5] );
tran (\sa_snapshot[31][38] , \sa_snapshot[31].r.part1[6] );
tran (\sa_snapshot[31][38] , \sa_snapshot[31].f.upper[6] );
tran (\sa_snapshot[31][39] , \sa_snapshot[31].r.part1[7] );
tran (\sa_snapshot[31][39] , \sa_snapshot[31].f.upper[7] );
tran (\sa_snapshot[31][40] , \sa_snapshot[31].r.part1[8] );
tran (\sa_snapshot[31][40] , \sa_snapshot[31].f.upper[8] );
tran (\sa_snapshot[31][41] , \sa_snapshot[31].r.part1[9] );
tran (\sa_snapshot[31][41] , \sa_snapshot[31].f.upper[9] );
tran (\sa_snapshot[31][42] , \sa_snapshot[31].r.part1[10] );
tran (\sa_snapshot[31][42] , \sa_snapshot[31].f.upper[10] );
tran (\sa_snapshot[31][43] , \sa_snapshot[31].r.part1[11] );
tran (\sa_snapshot[31][43] , \sa_snapshot[31].f.upper[11] );
tran (\sa_snapshot[31][44] , \sa_snapshot[31].r.part1[12] );
tran (\sa_snapshot[31][44] , \sa_snapshot[31].f.upper[12] );
tran (\sa_snapshot[31][45] , \sa_snapshot[31].r.part1[13] );
tran (\sa_snapshot[31][45] , \sa_snapshot[31].f.upper[13] );
tran (\sa_snapshot[31][46] , \sa_snapshot[31].r.part1[14] );
tran (\sa_snapshot[31][46] , \sa_snapshot[31].f.upper[14] );
tran (\sa_snapshot[31][47] , \sa_snapshot[31].r.part1[15] );
tran (\sa_snapshot[31][47] , \sa_snapshot[31].f.upper[15] );
tran (\sa_snapshot[31][48] , \sa_snapshot[31].r.part1[16] );
tran (\sa_snapshot[31][48] , \sa_snapshot[31].f.upper[16] );
tran (\sa_snapshot[31][49] , \sa_snapshot[31].r.part1[17] );
tran (\sa_snapshot[31][49] , \sa_snapshot[31].f.upper[17] );
tran (\sa_snapshot[31][50] , \sa_snapshot[31].r.part1[18] );
tran (\sa_snapshot[31][50] , \sa_snapshot[31].f.unused[0] );
tran (\sa_snapshot[31][51] , \sa_snapshot[31].r.part1[19] );
tran (\sa_snapshot[31][51] , \sa_snapshot[31].f.unused[1] );
tran (\sa_snapshot[31][52] , \sa_snapshot[31].r.part1[20] );
tran (\sa_snapshot[31][52] , \sa_snapshot[31].f.unused[2] );
tran (\sa_snapshot[31][53] , \sa_snapshot[31].r.part1[21] );
tran (\sa_snapshot[31][53] , \sa_snapshot[31].f.unused[3] );
tran (\sa_snapshot[31][54] , \sa_snapshot[31].r.part1[22] );
tran (\sa_snapshot[31][54] , \sa_snapshot[31].f.unused[4] );
tran (\sa_snapshot[31][55] , \sa_snapshot[31].r.part1[23] );
tran (\sa_snapshot[31][55] , \sa_snapshot[31].f.unused[5] );
tran (\sa_snapshot[31][56] , \sa_snapshot[31].r.part1[24] );
tran (\sa_snapshot[31][56] , \sa_snapshot[31].f.unused[6] );
tran (\sa_snapshot[31][57] , \sa_snapshot[31].r.part1[25] );
tran (\sa_snapshot[31][57] , \sa_snapshot[31].f.unused[7] );
tran (\sa_snapshot[31][58] , \sa_snapshot[31].r.part1[26] );
tran (\sa_snapshot[31][58] , \sa_snapshot[31].f.unused[8] );
tran (\sa_snapshot[31][59] , \sa_snapshot[31].r.part1[27] );
tran (\sa_snapshot[31][59] , \sa_snapshot[31].f.unused[9] );
tran (\sa_snapshot[31][60] , \sa_snapshot[31].r.part1[28] );
tran (\sa_snapshot[31][60] , \sa_snapshot[31].f.unused[10] );
tran (\sa_snapshot[31][61] , \sa_snapshot[31].r.part1[29] );
tran (\sa_snapshot[31][61] , \sa_snapshot[31].f.unused[11] );
tran (\sa_snapshot[31][62] , \sa_snapshot[31].r.part1[30] );
tran (\sa_snapshot[31][62] , \sa_snapshot[31].f.unused[12] );
tran (\sa_snapshot[31][63] , \sa_snapshot[31].r.part1[31] );
tran (\sa_snapshot[31][63] , \sa_snapshot[31].f.unused[13] );
tran (\sa_count[0][0] , \sa_count[0].r.part0[0] );
tran (\sa_count[0][0] , \sa_count[0].f.lower[0] );
tran (\sa_count[0][1] , \sa_count[0].r.part0[1] );
tran (\sa_count[0][1] , \sa_count[0].f.lower[1] );
tran (\sa_count[0][2] , \sa_count[0].r.part0[2] );
tran (\sa_count[0][2] , \sa_count[0].f.lower[2] );
tran (\sa_count[0][3] , \sa_count[0].r.part0[3] );
tran (\sa_count[0][3] , \sa_count[0].f.lower[3] );
tran (\sa_count[0][4] , \sa_count[0].r.part0[4] );
tran (\sa_count[0][4] , \sa_count[0].f.lower[4] );
tran (\sa_count[0][5] , \sa_count[0].r.part0[5] );
tran (\sa_count[0][5] , \sa_count[0].f.lower[5] );
tran (\sa_count[0][6] , \sa_count[0].r.part0[6] );
tran (\sa_count[0][6] , \sa_count[0].f.lower[6] );
tran (\sa_count[0][7] , \sa_count[0].r.part0[7] );
tran (\sa_count[0][7] , \sa_count[0].f.lower[7] );
tran (\sa_count[0][8] , \sa_count[0].r.part0[8] );
tran (\sa_count[0][8] , \sa_count[0].f.lower[8] );
tran (\sa_count[0][9] , \sa_count[0].r.part0[9] );
tran (\sa_count[0][9] , \sa_count[0].f.lower[9] );
tran (\sa_count[0][10] , \sa_count[0].r.part0[10] );
tran (\sa_count[0][10] , \sa_count[0].f.lower[10] );
tran (\sa_count[0][11] , \sa_count[0].r.part0[11] );
tran (\sa_count[0][11] , \sa_count[0].f.lower[11] );
tran (\sa_count[0][12] , \sa_count[0].r.part0[12] );
tran (\sa_count[0][12] , \sa_count[0].f.lower[12] );
tran (\sa_count[0][13] , \sa_count[0].r.part0[13] );
tran (\sa_count[0][13] , \sa_count[0].f.lower[13] );
tran (\sa_count[0][14] , \sa_count[0].r.part0[14] );
tran (\sa_count[0][14] , \sa_count[0].f.lower[14] );
tran (\sa_count[0][15] , \sa_count[0].r.part0[15] );
tran (\sa_count[0][15] , \sa_count[0].f.lower[15] );
tran (\sa_count[0][16] , \sa_count[0].r.part0[16] );
tran (\sa_count[0][16] , \sa_count[0].f.lower[16] );
tran (\sa_count[0][17] , \sa_count[0].r.part0[17] );
tran (\sa_count[0][17] , \sa_count[0].f.lower[17] );
tran (\sa_count[0][18] , \sa_count[0].r.part0[18] );
tran (\sa_count[0][18] , \sa_count[0].f.lower[18] );
tran (\sa_count[0][19] , \sa_count[0].r.part0[19] );
tran (\sa_count[0][19] , \sa_count[0].f.lower[19] );
tran (\sa_count[0][20] , \sa_count[0].r.part0[20] );
tran (\sa_count[0][20] , \sa_count[0].f.lower[20] );
tran (\sa_count[0][21] , \sa_count[0].r.part0[21] );
tran (\sa_count[0][21] , \sa_count[0].f.lower[21] );
tran (\sa_count[0][22] , \sa_count[0].r.part0[22] );
tran (\sa_count[0][22] , \sa_count[0].f.lower[22] );
tran (\sa_count[0][23] , \sa_count[0].r.part0[23] );
tran (\sa_count[0][23] , \sa_count[0].f.lower[23] );
tran (\sa_count[0][24] , \sa_count[0].r.part0[24] );
tran (\sa_count[0][24] , \sa_count[0].f.lower[24] );
tran (\sa_count[0][25] , \sa_count[0].r.part0[25] );
tran (\sa_count[0][25] , \sa_count[0].f.lower[25] );
tran (\sa_count[0][26] , \sa_count[0].r.part0[26] );
tran (\sa_count[0][26] , \sa_count[0].f.lower[26] );
tran (\sa_count[0][27] , \sa_count[0].r.part0[27] );
tran (\sa_count[0][27] , \sa_count[0].f.lower[27] );
tran (\sa_count[0][28] , \sa_count[0].r.part0[28] );
tran (\sa_count[0][28] , \sa_count[0].f.lower[28] );
tran (\sa_count[0][29] , \sa_count[0].r.part0[29] );
tran (\sa_count[0][29] , \sa_count[0].f.lower[29] );
tran (\sa_count[0][30] , \sa_count[0].r.part0[30] );
tran (\sa_count[0][30] , \sa_count[0].f.lower[30] );
tran (\sa_count[0][31] , \sa_count[0].r.part0[31] );
tran (\sa_count[0][31] , \sa_count[0].f.lower[31] );
tran (\sa_count[0][32] , \sa_count[0].r.part1[0] );
tran (\sa_count[0][32] , \sa_count[0].f.upper[0] );
tran (\sa_count[0][33] , \sa_count[0].r.part1[1] );
tran (\sa_count[0][33] , \sa_count[0].f.upper[1] );
tran (\sa_count[0][34] , \sa_count[0].r.part1[2] );
tran (\sa_count[0][34] , \sa_count[0].f.upper[2] );
tran (\sa_count[0][35] , \sa_count[0].r.part1[3] );
tran (\sa_count[0][35] , \sa_count[0].f.upper[3] );
tran (\sa_count[0][36] , \sa_count[0].r.part1[4] );
tran (\sa_count[0][36] , \sa_count[0].f.upper[4] );
tran (\sa_count[0][37] , \sa_count[0].r.part1[5] );
tran (\sa_count[0][37] , \sa_count[0].f.upper[5] );
tran (\sa_count[0][38] , \sa_count[0].r.part1[6] );
tran (\sa_count[0][38] , \sa_count[0].f.upper[6] );
tran (\sa_count[0][39] , \sa_count[0].r.part1[7] );
tran (\sa_count[0][39] , \sa_count[0].f.upper[7] );
tran (\sa_count[0][40] , \sa_count[0].r.part1[8] );
tran (\sa_count[0][40] , \sa_count[0].f.upper[8] );
tran (\sa_count[0][41] , \sa_count[0].r.part1[9] );
tran (\sa_count[0][41] , \sa_count[0].f.upper[9] );
tran (\sa_count[0][42] , \sa_count[0].r.part1[10] );
tran (\sa_count[0][42] , \sa_count[0].f.upper[10] );
tran (\sa_count[0][43] , \sa_count[0].r.part1[11] );
tran (\sa_count[0][43] , \sa_count[0].f.upper[11] );
tran (\sa_count[0][44] , \sa_count[0].r.part1[12] );
tran (\sa_count[0][44] , \sa_count[0].f.upper[12] );
tran (\sa_count[0][45] , \sa_count[0].r.part1[13] );
tran (\sa_count[0][45] , \sa_count[0].f.upper[13] );
tran (\sa_count[0][46] , \sa_count[0].r.part1[14] );
tran (\sa_count[0][46] , \sa_count[0].f.upper[14] );
tran (\sa_count[0][47] , \sa_count[0].r.part1[15] );
tran (\sa_count[0][47] , \sa_count[0].f.upper[15] );
tran (\sa_count[0][48] , \sa_count[0].r.part1[16] );
tran (\sa_count[0][48] , \sa_count[0].f.upper[16] );
tran (\sa_count[0][49] , \sa_count[0].r.part1[17] );
tran (\sa_count[0][49] , \sa_count[0].f.upper[17] );
tran (\sa_count[0][50] , \sa_count[0].r.part1[18] );
tran (\sa_count[0][50] , \sa_count[0].f.unused[0] );
tran (\sa_count[0][51] , \sa_count[0].r.part1[19] );
tran (\sa_count[0][51] , \sa_count[0].f.unused[1] );
tran (\sa_count[0][52] , \sa_count[0].r.part1[20] );
tran (\sa_count[0][52] , \sa_count[0].f.unused[2] );
tran (\sa_count[0][53] , \sa_count[0].r.part1[21] );
tran (\sa_count[0][53] , \sa_count[0].f.unused[3] );
tran (\sa_count[0][54] , \sa_count[0].r.part1[22] );
tran (\sa_count[0][54] , \sa_count[0].f.unused[4] );
tran (\sa_count[0][55] , \sa_count[0].r.part1[23] );
tran (\sa_count[0][55] , \sa_count[0].f.unused[5] );
tran (\sa_count[0][56] , \sa_count[0].r.part1[24] );
tran (\sa_count[0][56] , \sa_count[0].f.unused[6] );
tran (\sa_count[0][57] , \sa_count[0].r.part1[25] );
tran (\sa_count[0][57] , \sa_count[0].f.unused[7] );
tran (\sa_count[0][58] , \sa_count[0].r.part1[26] );
tran (\sa_count[0][58] , \sa_count[0].f.unused[8] );
tran (\sa_count[0][59] , \sa_count[0].r.part1[27] );
tran (\sa_count[0][59] , \sa_count[0].f.unused[9] );
tran (\sa_count[0][60] , \sa_count[0].r.part1[28] );
tran (\sa_count[0][60] , \sa_count[0].f.unused[10] );
tran (\sa_count[0][61] , \sa_count[0].r.part1[29] );
tran (\sa_count[0][61] , \sa_count[0].f.unused[11] );
tran (\sa_count[0][62] , \sa_count[0].r.part1[30] );
tran (\sa_count[0][62] , \sa_count[0].f.unused[12] );
tran (\sa_count[0][63] , \sa_count[0].r.part1[31] );
tran (\sa_count[0][63] , \sa_count[0].f.unused[13] );
tran (\sa_count[1][0] , \sa_count[1].r.part0[0] );
tran (\sa_count[1][0] , \sa_count[1].f.lower[0] );
tran (\sa_count[1][1] , \sa_count[1].r.part0[1] );
tran (\sa_count[1][1] , \sa_count[1].f.lower[1] );
tran (\sa_count[1][2] , \sa_count[1].r.part0[2] );
tran (\sa_count[1][2] , \sa_count[1].f.lower[2] );
tran (\sa_count[1][3] , \sa_count[1].r.part0[3] );
tran (\sa_count[1][3] , \sa_count[1].f.lower[3] );
tran (\sa_count[1][4] , \sa_count[1].r.part0[4] );
tran (\sa_count[1][4] , \sa_count[1].f.lower[4] );
tran (\sa_count[1][5] , \sa_count[1].r.part0[5] );
tran (\sa_count[1][5] , \sa_count[1].f.lower[5] );
tran (\sa_count[1][6] , \sa_count[1].r.part0[6] );
tran (\sa_count[1][6] , \sa_count[1].f.lower[6] );
tran (\sa_count[1][7] , \sa_count[1].r.part0[7] );
tran (\sa_count[1][7] , \sa_count[1].f.lower[7] );
tran (\sa_count[1][8] , \sa_count[1].r.part0[8] );
tran (\sa_count[1][8] , \sa_count[1].f.lower[8] );
tran (\sa_count[1][9] , \sa_count[1].r.part0[9] );
tran (\sa_count[1][9] , \sa_count[1].f.lower[9] );
tran (\sa_count[1][10] , \sa_count[1].r.part0[10] );
tran (\sa_count[1][10] , \sa_count[1].f.lower[10] );
tran (\sa_count[1][11] , \sa_count[1].r.part0[11] );
tran (\sa_count[1][11] , \sa_count[1].f.lower[11] );
tran (\sa_count[1][12] , \sa_count[1].r.part0[12] );
tran (\sa_count[1][12] , \sa_count[1].f.lower[12] );
tran (\sa_count[1][13] , \sa_count[1].r.part0[13] );
tran (\sa_count[1][13] , \sa_count[1].f.lower[13] );
tran (\sa_count[1][14] , \sa_count[1].r.part0[14] );
tran (\sa_count[1][14] , \sa_count[1].f.lower[14] );
tran (\sa_count[1][15] , \sa_count[1].r.part0[15] );
tran (\sa_count[1][15] , \sa_count[1].f.lower[15] );
tran (\sa_count[1][16] , \sa_count[1].r.part0[16] );
tran (\sa_count[1][16] , \sa_count[1].f.lower[16] );
tran (\sa_count[1][17] , \sa_count[1].r.part0[17] );
tran (\sa_count[1][17] , \sa_count[1].f.lower[17] );
tran (\sa_count[1][18] , \sa_count[1].r.part0[18] );
tran (\sa_count[1][18] , \sa_count[1].f.lower[18] );
tran (\sa_count[1][19] , \sa_count[1].r.part0[19] );
tran (\sa_count[1][19] , \sa_count[1].f.lower[19] );
tran (\sa_count[1][20] , \sa_count[1].r.part0[20] );
tran (\sa_count[1][20] , \sa_count[1].f.lower[20] );
tran (\sa_count[1][21] , \sa_count[1].r.part0[21] );
tran (\sa_count[1][21] , \sa_count[1].f.lower[21] );
tran (\sa_count[1][22] , \sa_count[1].r.part0[22] );
tran (\sa_count[1][22] , \sa_count[1].f.lower[22] );
tran (\sa_count[1][23] , \sa_count[1].r.part0[23] );
tran (\sa_count[1][23] , \sa_count[1].f.lower[23] );
tran (\sa_count[1][24] , \sa_count[1].r.part0[24] );
tran (\sa_count[1][24] , \sa_count[1].f.lower[24] );
tran (\sa_count[1][25] , \sa_count[1].r.part0[25] );
tran (\sa_count[1][25] , \sa_count[1].f.lower[25] );
tran (\sa_count[1][26] , \sa_count[1].r.part0[26] );
tran (\sa_count[1][26] , \sa_count[1].f.lower[26] );
tran (\sa_count[1][27] , \sa_count[1].r.part0[27] );
tran (\sa_count[1][27] , \sa_count[1].f.lower[27] );
tran (\sa_count[1][28] , \sa_count[1].r.part0[28] );
tran (\sa_count[1][28] , \sa_count[1].f.lower[28] );
tran (\sa_count[1][29] , \sa_count[1].r.part0[29] );
tran (\sa_count[1][29] , \sa_count[1].f.lower[29] );
tran (\sa_count[1][30] , \sa_count[1].r.part0[30] );
tran (\sa_count[1][30] , \sa_count[1].f.lower[30] );
tran (\sa_count[1][31] , \sa_count[1].r.part0[31] );
tran (\sa_count[1][31] , \sa_count[1].f.lower[31] );
tran (\sa_count[1][32] , \sa_count[1].r.part1[0] );
tran (\sa_count[1][32] , \sa_count[1].f.upper[0] );
tran (\sa_count[1][33] , \sa_count[1].r.part1[1] );
tran (\sa_count[1][33] , \sa_count[1].f.upper[1] );
tran (\sa_count[1][34] , \sa_count[1].r.part1[2] );
tran (\sa_count[1][34] , \sa_count[1].f.upper[2] );
tran (\sa_count[1][35] , \sa_count[1].r.part1[3] );
tran (\sa_count[1][35] , \sa_count[1].f.upper[3] );
tran (\sa_count[1][36] , \sa_count[1].r.part1[4] );
tran (\sa_count[1][36] , \sa_count[1].f.upper[4] );
tran (\sa_count[1][37] , \sa_count[1].r.part1[5] );
tran (\sa_count[1][37] , \sa_count[1].f.upper[5] );
tran (\sa_count[1][38] , \sa_count[1].r.part1[6] );
tran (\sa_count[1][38] , \sa_count[1].f.upper[6] );
tran (\sa_count[1][39] , \sa_count[1].r.part1[7] );
tran (\sa_count[1][39] , \sa_count[1].f.upper[7] );
tran (\sa_count[1][40] , \sa_count[1].r.part1[8] );
tran (\sa_count[1][40] , \sa_count[1].f.upper[8] );
tran (\sa_count[1][41] , \sa_count[1].r.part1[9] );
tran (\sa_count[1][41] , \sa_count[1].f.upper[9] );
tran (\sa_count[1][42] , \sa_count[1].r.part1[10] );
tran (\sa_count[1][42] , \sa_count[1].f.upper[10] );
tran (\sa_count[1][43] , \sa_count[1].r.part1[11] );
tran (\sa_count[1][43] , \sa_count[1].f.upper[11] );
tran (\sa_count[1][44] , \sa_count[1].r.part1[12] );
tran (\sa_count[1][44] , \sa_count[1].f.upper[12] );
tran (\sa_count[1][45] , \sa_count[1].r.part1[13] );
tran (\sa_count[1][45] , \sa_count[1].f.upper[13] );
tran (\sa_count[1][46] , \sa_count[1].r.part1[14] );
tran (\sa_count[1][46] , \sa_count[1].f.upper[14] );
tran (\sa_count[1][47] , \sa_count[1].r.part1[15] );
tran (\sa_count[1][47] , \sa_count[1].f.upper[15] );
tran (\sa_count[1][48] , \sa_count[1].r.part1[16] );
tran (\sa_count[1][48] , \sa_count[1].f.upper[16] );
tran (\sa_count[1][49] , \sa_count[1].r.part1[17] );
tran (\sa_count[1][49] , \sa_count[1].f.upper[17] );
tran (\sa_count[1][50] , \sa_count[1].r.part1[18] );
tran (\sa_count[1][50] , \sa_count[1].f.unused[0] );
tran (\sa_count[1][51] , \sa_count[1].r.part1[19] );
tran (\sa_count[1][51] , \sa_count[1].f.unused[1] );
tran (\sa_count[1][52] , \sa_count[1].r.part1[20] );
tran (\sa_count[1][52] , \sa_count[1].f.unused[2] );
tran (\sa_count[1][53] , \sa_count[1].r.part1[21] );
tran (\sa_count[1][53] , \sa_count[1].f.unused[3] );
tran (\sa_count[1][54] , \sa_count[1].r.part1[22] );
tran (\sa_count[1][54] , \sa_count[1].f.unused[4] );
tran (\sa_count[1][55] , \sa_count[1].r.part1[23] );
tran (\sa_count[1][55] , \sa_count[1].f.unused[5] );
tran (\sa_count[1][56] , \sa_count[1].r.part1[24] );
tran (\sa_count[1][56] , \sa_count[1].f.unused[6] );
tran (\sa_count[1][57] , \sa_count[1].r.part1[25] );
tran (\sa_count[1][57] , \sa_count[1].f.unused[7] );
tran (\sa_count[1][58] , \sa_count[1].r.part1[26] );
tran (\sa_count[1][58] , \sa_count[1].f.unused[8] );
tran (\sa_count[1][59] , \sa_count[1].r.part1[27] );
tran (\sa_count[1][59] , \sa_count[1].f.unused[9] );
tran (\sa_count[1][60] , \sa_count[1].r.part1[28] );
tran (\sa_count[1][60] , \sa_count[1].f.unused[10] );
tran (\sa_count[1][61] , \sa_count[1].r.part1[29] );
tran (\sa_count[1][61] , \sa_count[1].f.unused[11] );
tran (\sa_count[1][62] , \sa_count[1].r.part1[30] );
tran (\sa_count[1][62] , \sa_count[1].f.unused[12] );
tran (\sa_count[1][63] , \sa_count[1].r.part1[31] );
tran (\sa_count[1][63] , \sa_count[1].f.unused[13] );
tran (\sa_count[2][0] , \sa_count[2].r.part0[0] );
tran (\sa_count[2][0] , \sa_count[2].f.lower[0] );
tran (\sa_count[2][1] , \sa_count[2].r.part0[1] );
tran (\sa_count[2][1] , \sa_count[2].f.lower[1] );
tran (\sa_count[2][2] , \sa_count[2].r.part0[2] );
tran (\sa_count[2][2] , \sa_count[2].f.lower[2] );
tran (\sa_count[2][3] , \sa_count[2].r.part0[3] );
tran (\sa_count[2][3] , \sa_count[2].f.lower[3] );
tran (\sa_count[2][4] , \sa_count[2].r.part0[4] );
tran (\sa_count[2][4] , \sa_count[2].f.lower[4] );
tran (\sa_count[2][5] , \sa_count[2].r.part0[5] );
tran (\sa_count[2][5] , \sa_count[2].f.lower[5] );
tran (\sa_count[2][6] , \sa_count[2].r.part0[6] );
tran (\sa_count[2][6] , \sa_count[2].f.lower[6] );
tran (\sa_count[2][7] , \sa_count[2].r.part0[7] );
tran (\sa_count[2][7] , \sa_count[2].f.lower[7] );
tran (\sa_count[2][8] , \sa_count[2].r.part0[8] );
tran (\sa_count[2][8] , \sa_count[2].f.lower[8] );
tran (\sa_count[2][9] , \sa_count[2].r.part0[9] );
tran (\sa_count[2][9] , \sa_count[2].f.lower[9] );
tran (\sa_count[2][10] , \sa_count[2].r.part0[10] );
tran (\sa_count[2][10] , \sa_count[2].f.lower[10] );
tran (\sa_count[2][11] , \sa_count[2].r.part0[11] );
tran (\sa_count[2][11] , \sa_count[2].f.lower[11] );
tran (\sa_count[2][12] , \sa_count[2].r.part0[12] );
tran (\sa_count[2][12] , \sa_count[2].f.lower[12] );
tran (\sa_count[2][13] , \sa_count[2].r.part0[13] );
tran (\sa_count[2][13] , \sa_count[2].f.lower[13] );
tran (\sa_count[2][14] , \sa_count[2].r.part0[14] );
tran (\sa_count[2][14] , \sa_count[2].f.lower[14] );
tran (\sa_count[2][15] , \sa_count[2].r.part0[15] );
tran (\sa_count[2][15] , \sa_count[2].f.lower[15] );
tran (\sa_count[2][16] , \sa_count[2].r.part0[16] );
tran (\sa_count[2][16] , \sa_count[2].f.lower[16] );
tran (\sa_count[2][17] , \sa_count[2].r.part0[17] );
tran (\sa_count[2][17] , \sa_count[2].f.lower[17] );
tran (\sa_count[2][18] , \sa_count[2].r.part0[18] );
tran (\sa_count[2][18] , \sa_count[2].f.lower[18] );
tran (\sa_count[2][19] , \sa_count[2].r.part0[19] );
tran (\sa_count[2][19] , \sa_count[2].f.lower[19] );
tran (\sa_count[2][20] , \sa_count[2].r.part0[20] );
tran (\sa_count[2][20] , \sa_count[2].f.lower[20] );
tran (\sa_count[2][21] , \sa_count[2].r.part0[21] );
tran (\sa_count[2][21] , \sa_count[2].f.lower[21] );
tran (\sa_count[2][22] , \sa_count[2].r.part0[22] );
tran (\sa_count[2][22] , \sa_count[2].f.lower[22] );
tran (\sa_count[2][23] , \sa_count[2].r.part0[23] );
tran (\sa_count[2][23] , \sa_count[2].f.lower[23] );
tran (\sa_count[2][24] , \sa_count[2].r.part0[24] );
tran (\sa_count[2][24] , \sa_count[2].f.lower[24] );
tran (\sa_count[2][25] , \sa_count[2].r.part0[25] );
tran (\sa_count[2][25] , \sa_count[2].f.lower[25] );
tran (\sa_count[2][26] , \sa_count[2].r.part0[26] );
tran (\sa_count[2][26] , \sa_count[2].f.lower[26] );
tran (\sa_count[2][27] , \sa_count[2].r.part0[27] );
tran (\sa_count[2][27] , \sa_count[2].f.lower[27] );
tran (\sa_count[2][28] , \sa_count[2].r.part0[28] );
tran (\sa_count[2][28] , \sa_count[2].f.lower[28] );
tran (\sa_count[2][29] , \sa_count[2].r.part0[29] );
tran (\sa_count[2][29] , \sa_count[2].f.lower[29] );
tran (\sa_count[2][30] , \sa_count[2].r.part0[30] );
tran (\sa_count[2][30] , \sa_count[2].f.lower[30] );
tran (\sa_count[2][31] , \sa_count[2].r.part0[31] );
tran (\sa_count[2][31] , \sa_count[2].f.lower[31] );
tran (\sa_count[2][32] , \sa_count[2].r.part1[0] );
tran (\sa_count[2][32] , \sa_count[2].f.upper[0] );
tran (\sa_count[2][33] , \sa_count[2].r.part1[1] );
tran (\sa_count[2][33] , \sa_count[2].f.upper[1] );
tran (\sa_count[2][34] , \sa_count[2].r.part1[2] );
tran (\sa_count[2][34] , \sa_count[2].f.upper[2] );
tran (\sa_count[2][35] , \sa_count[2].r.part1[3] );
tran (\sa_count[2][35] , \sa_count[2].f.upper[3] );
tran (\sa_count[2][36] , \sa_count[2].r.part1[4] );
tran (\sa_count[2][36] , \sa_count[2].f.upper[4] );
tran (\sa_count[2][37] , \sa_count[2].r.part1[5] );
tran (\sa_count[2][37] , \sa_count[2].f.upper[5] );
tran (\sa_count[2][38] , \sa_count[2].r.part1[6] );
tran (\sa_count[2][38] , \sa_count[2].f.upper[6] );
tran (\sa_count[2][39] , \sa_count[2].r.part1[7] );
tran (\sa_count[2][39] , \sa_count[2].f.upper[7] );
tran (\sa_count[2][40] , \sa_count[2].r.part1[8] );
tran (\sa_count[2][40] , \sa_count[2].f.upper[8] );
tran (\sa_count[2][41] , \sa_count[2].r.part1[9] );
tran (\sa_count[2][41] , \sa_count[2].f.upper[9] );
tran (\sa_count[2][42] , \sa_count[2].r.part1[10] );
tran (\sa_count[2][42] , \sa_count[2].f.upper[10] );
tran (\sa_count[2][43] , \sa_count[2].r.part1[11] );
tran (\sa_count[2][43] , \sa_count[2].f.upper[11] );
tran (\sa_count[2][44] , \sa_count[2].r.part1[12] );
tran (\sa_count[2][44] , \sa_count[2].f.upper[12] );
tran (\sa_count[2][45] , \sa_count[2].r.part1[13] );
tran (\sa_count[2][45] , \sa_count[2].f.upper[13] );
tran (\sa_count[2][46] , \sa_count[2].r.part1[14] );
tran (\sa_count[2][46] , \sa_count[2].f.upper[14] );
tran (\sa_count[2][47] , \sa_count[2].r.part1[15] );
tran (\sa_count[2][47] , \sa_count[2].f.upper[15] );
tran (\sa_count[2][48] , \sa_count[2].r.part1[16] );
tran (\sa_count[2][48] , \sa_count[2].f.upper[16] );
tran (\sa_count[2][49] , \sa_count[2].r.part1[17] );
tran (\sa_count[2][49] , \sa_count[2].f.upper[17] );
tran (\sa_count[2][50] , \sa_count[2].r.part1[18] );
tran (\sa_count[2][50] , \sa_count[2].f.unused[0] );
tran (\sa_count[2][51] , \sa_count[2].r.part1[19] );
tran (\sa_count[2][51] , \sa_count[2].f.unused[1] );
tran (\sa_count[2][52] , \sa_count[2].r.part1[20] );
tran (\sa_count[2][52] , \sa_count[2].f.unused[2] );
tran (\sa_count[2][53] , \sa_count[2].r.part1[21] );
tran (\sa_count[2][53] , \sa_count[2].f.unused[3] );
tran (\sa_count[2][54] , \sa_count[2].r.part1[22] );
tran (\sa_count[2][54] , \sa_count[2].f.unused[4] );
tran (\sa_count[2][55] , \sa_count[2].r.part1[23] );
tran (\sa_count[2][55] , \sa_count[2].f.unused[5] );
tran (\sa_count[2][56] , \sa_count[2].r.part1[24] );
tran (\sa_count[2][56] , \sa_count[2].f.unused[6] );
tran (\sa_count[2][57] , \sa_count[2].r.part1[25] );
tran (\sa_count[2][57] , \sa_count[2].f.unused[7] );
tran (\sa_count[2][58] , \sa_count[2].r.part1[26] );
tran (\sa_count[2][58] , \sa_count[2].f.unused[8] );
tran (\sa_count[2][59] , \sa_count[2].r.part1[27] );
tran (\sa_count[2][59] , \sa_count[2].f.unused[9] );
tran (\sa_count[2][60] , \sa_count[2].r.part1[28] );
tran (\sa_count[2][60] , \sa_count[2].f.unused[10] );
tran (\sa_count[2][61] , \sa_count[2].r.part1[29] );
tran (\sa_count[2][61] , \sa_count[2].f.unused[11] );
tran (\sa_count[2][62] , \sa_count[2].r.part1[30] );
tran (\sa_count[2][62] , \sa_count[2].f.unused[12] );
tran (\sa_count[2][63] , \sa_count[2].r.part1[31] );
tran (\sa_count[2][63] , \sa_count[2].f.unused[13] );
tran (\sa_count[3][0] , \sa_count[3].r.part0[0] );
tran (\sa_count[3][0] , \sa_count[3].f.lower[0] );
tran (\sa_count[3][1] , \sa_count[3].r.part0[1] );
tran (\sa_count[3][1] , \sa_count[3].f.lower[1] );
tran (\sa_count[3][2] , \sa_count[3].r.part0[2] );
tran (\sa_count[3][2] , \sa_count[3].f.lower[2] );
tran (\sa_count[3][3] , \sa_count[3].r.part0[3] );
tran (\sa_count[3][3] , \sa_count[3].f.lower[3] );
tran (\sa_count[3][4] , \sa_count[3].r.part0[4] );
tran (\sa_count[3][4] , \sa_count[3].f.lower[4] );
tran (\sa_count[3][5] , \sa_count[3].r.part0[5] );
tran (\sa_count[3][5] , \sa_count[3].f.lower[5] );
tran (\sa_count[3][6] , \sa_count[3].r.part0[6] );
tran (\sa_count[3][6] , \sa_count[3].f.lower[6] );
tran (\sa_count[3][7] , \sa_count[3].r.part0[7] );
tran (\sa_count[3][7] , \sa_count[3].f.lower[7] );
tran (\sa_count[3][8] , \sa_count[3].r.part0[8] );
tran (\sa_count[3][8] , \sa_count[3].f.lower[8] );
tran (\sa_count[3][9] , \sa_count[3].r.part0[9] );
tran (\sa_count[3][9] , \sa_count[3].f.lower[9] );
tran (\sa_count[3][10] , \sa_count[3].r.part0[10] );
tran (\sa_count[3][10] , \sa_count[3].f.lower[10] );
tran (\sa_count[3][11] , \sa_count[3].r.part0[11] );
tran (\sa_count[3][11] , \sa_count[3].f.lower[11] );
tran (\sa_count[3][12] , \sa_count[3].r.part0[12] );
tran (\sa_count[3][12] , \sa_count[3].f.lower[12] );
tran (\sa_count[3][13] , \sa_count[3].r.part0[13] );
tran (\sa_count[3][13] , \sa_count[3].f.lower[13] );
tran (\sa_count[3][14] , \sa_count[3].r.part0[14] );
tran (\sa_count[3][14] , \sa_count[3].f.lower[14] );
tran (\sa_count[3][15] , \sa_count[3].r.part0[15] );
tran (\sa_count[3][15] , \sa_count[3].f.lower[15] );
tran (\sa_count[3][16] , \sa_count[3].r.part0[16] );
tran (\sa_count[3][16] , \sa_count[3].f.lower[16] );
tran (\sa_count[3][17] , \sa_count[3].r.part0[17] );
tran (\sa_count[3][17] , \sa_count[3].f.lower[17] );
tran (\sa_count[3][18] , \sa_count[3].r.part0[18] );
tran (\sa_count[3][18] , \sa_count[3].f.lower[18] );
tran (\sa_count[3][19] , \sa_count[3].r.part0[19] );
tran (\sa_count[3][19] , \sa_count[3].f.lower[19] );
tran (\sa_count[3][20] , \sa_count[3].r.part0[20] );
tran (\sa_count[3][20] , \sa_count[3].f.lower[20] );
tran (\sa_count[3][21] , \sa_count[3].r.part0[21] );
tran (\sa_count[3][21] , \sa_count[3].f.lower[21] );
tran (\sa_count[3][22] , \sa_count[3].r.part0[22] );
tran (\sa_count[3][22] , \sa_count[3].f.lower[22] );
tran (\sa_count[3][23] , \sa_count[3].r.part0[23] );
tran (\sa_count[3][23] , \sa_count[3].f.lower[23] );
tran (\sa_count[3][24] , \sa_count[3].r.part0[24] );
tran (\sa_count[3][24] , \sa_count[3].f.lower[24] );
tran (\sa_count[3][25] , \sa_count[3].r.part0[25] );
tran (\sa_count[3][25] , \sa_count[3].f.lower[25] );
tran (\sa_count[3][26] , \sa_count[3].r.part0[26] );
tran (\sa_count[3][26] , \sa_count[3].f.lower[26] );
tran (\sa_count[3][27] , \sa_count[3].r.part0[27] );
tran (\sa_count[3][27] , \sa_count[3].f.lower[27] );
tran (\sa_count[3][28] , \sa_count[3].r.part0[28] );
tran (\sa_count[3][28] , \sa_count[3].f.lower[28] );
tran (\sa_count[3][29] , \sa_count[3].r.part0[29] );
tran (\sa_count[3][29] , \sa_count[3].f.lower[29] );
tran (\sa_count[3][30] , \sa_count[3].r.part0[30] );
tran (\sa_count[3][30] , \sa_count[3].f.lower[30] );
tran (\sa_count[3][31] , \sa_count[3].r.part0[31] );
tran (\sa_count[3][31] , \sa_count[3].f.lower[31] );
tran (\sa_count[3][32] , \sa_count[3].r.part1[0] );
tran (\sa_count[3][32] , \sa_count[3].f.upper[0] );
tran (\sa_count[3][33] , \sa_count[3].r.part1[1] );
tran (\sa_count[3][33] , \sa_count[3].f.upper[1] );
tran (\sa_count[3][34] , \sa_count[3].r.part1[2] );
tran (\sa_count[3][34] , \sa_count[3].f.upper[2] );
tran (\sa_count[3][35] , \sa_count[3].r.part1[3] );
tran (\sa_count[3][35] , \sa_count[3].f.upper[3] );
tran (\sa_count[3][36] , \sa_count[3].r.part1[4] );
tran (\sa_count[3][36] , \sa_count[3].f.upper[4] );
tran (\sa_count[3][37] , \sa_count[3].r.part1[5] );
tran (\sa_count[3][37] , \sa_count[3].f.upper[5] );
tran (\sa_count[3][38] , \sa_count[3].r.part1[6] );
tran (\sa_count[3][38] , \sa_count[3].f.upper[6] );
tran (\sa_count[3][39] , \sa_count[3].r.part1[7] );
tran (\sa_count[3][39] , \sa_count[3].f.upper[7] );
tran (\sa_count[3][40] , \sa_count[3].r.part1[8] );
tran (\sa_count[3][40] , \sa_count[3].f.upper[8] );
tran (\sa_count[3][41] , \sa_count[3].r.part1[9] );
tran (\sa_count[3][41] , \sa_count[3].f.upper[9] );
tran (\sa_count[3][42] , \sa_count[3].r.part1[10] );
tran (\sa_count[3][42] , \sa_count[3].f.upper[10] );
tran (\sa_count[3][43] , \sa_count[3].r.part1[11] );
tran (\sa_count[3][43] , \sa_count[3].f.upper[11] );
tran (\sa_count[3][44] , \sa_count[3].r.part1[12] );
tran (\sa_count[3][44] , \sa_count[3].f.upper[12] );
tran (\sa_count[3][45] , \sa_count[3].r.part1[13] );
tran (\sa_count[3][45] , \sa_count[3].f.upper[13] );
tran (\sa_count[3][46] , \sa_count[3].r.part1[14] );
tran (\sa_count[3][46] , \sa_count[3].f.upper[14] );
tran (\sa_count[3][47] , \sa_count[3].r.part1[15] );
tran (\sa_count[3][47] , \sa_count[3].f.upper[15] );
tran (\sa_count[3][48] , \sa_count[3].r.part1[16] );
tran (\sa_count[3][48] , \sa_count[3].f.upper[16] );
tran (\sa_count[3][49] , \sa_count[3].r.part1[17] );
tran (\sa_count[3][49] , \sa_count[3].f.upper[17] );
tran (\sa_count[3][50] , \sa_count[3].r.part1[18] );
tran (\sa_count[3][50] , \sa_count[3].f.unused[0] );
tran (\sa_count[3][51] , \sa_count[3].r.part1[19] );
tran (\sa_count[3][51] , \sa_count[3].f.unused[1] );
tran (\sa_count[3][52] , \sa_count[3].r.part1[20] );
tran (\sa_count[3][52] , \sa_count[3].f.unused[2] );
tran (\sa_count[3][53] , \sa_count[3].r.part1[21] );
tran (\sa_count[3][53] , \sa_count[3].f.unused[3] );
tran (\sa_count[3][54] , \sa_count[3].r.part1[22] );
tran (\sa_count[3][54] , \sa_count[3].f.unused[4] );
tran (\sa_count[3][55] , \sa_count[3].r.part1[23] );
tran (\sa_count[3][55] , \sa_count[3].f.unused[5] );
tran (\sa_count[3][56] , \sa_count[3].r.part1[24] );
tran (\sa_count[3][56] , \sa_count[3].f.unused[6] );
tran (\sa_count[3][57] , \sa_count[3].r.part1[25] );
tran (\sa_count[3][57] , \sa_count[3].f.unused[7] );
tran (\sa_count[3][58] , \sa_count[3].r.part1[26] );
tran (\sa_count[3][58] , \sa_count[3].f.unused[8] );
tran (\sa_count[3][59] , \sa_count[3].r.part1[27] );
tran (\sa_count[3][59] , \sa_count[3].f.unused[9] );
tran (\sa_count[3][60] , \sa_count[3].r.part1[28] );
tran (\sa_count[3][60] , \sa_count[3].f.unused[10] );
tran (\sa_count[3][61] , \sa_count[3].r.part1[29] );
tran (\sa_count[3][61] , \sa_count[3].f.unused[11] );
tran (\sa_count[3][62] , \sa_count[3].r.part1[30] );
tran (\sa_count[3][62] , \sa_count[3].f.unused[12] );
tran (\sa_count[3][63] , \sa_count[3].r.part1[31] );
tran (\sa_count[3][63] , \sa_count[3].f.unused[13] );
tran (\sa_count[4][0] , \sa_count[4].r.part0[0] );
tran (\sa_count[4][0] , \sa_count[4].f.lower[0] );
tran (\sa_count[4][1] , \sa_count[4].r.part0[1] );
tran (\sa_count[4][1] , \sa_count[4].f.lower[1] );
tran (\sa_count[4][2] , \sa_count[4].r.part0[2] );
tran (\sa_count[4][2] , \sa_count[4].f.lower[2] );
tran (\sa_count[4][3] , \sa_count[4].r.part0[3] );
tran (\sa_count[4][3] , \sa_count[4].f.lower[3] );
tran (\sa_count[4][4] , \sa_count[4].r.part0[4] );
tran (\sa_count[4][4] , \sa_count[4].f.lower[4] );
tran (\sa_count[4][5] , \sa_count[4].r.part0[5] );
tran (\sa_count[4][5] , \sa_count[4].f.lower[5] );
tran (\sa_count[4][6] , \sa_count[4].r.part0[6] );
tran (\sa_count[4][6] , \sa_count[4].f.lower[6] );
tran (\sa_count[4][7] , \sa_count[4].r.part0[7] );
tran (\sa_count[4][7] , \sa_count[4].f.lower[7] );
tran (\sa_count[4][8] , \sa_count[4].r.part0[8] );
tran (\sa_count[4][8] , \sa_count[4].f.lower[8] );
tran (\sa_count[4][9] , \sa_count[4].r.part0[9] );
tran (\sa_count[4][9] , \sa_count[4].f.lower[9] );
tran (\sa_count[4][10] , \sa_count[4].r.part0[10] );
tran (\sa_count[4][10] , \sa_count[4].f.lower[10] );
tran (\sa_count[4][11] , \sa_count[4].r.part0[11] );
tran (\sa_count[4][11] , \sa_count[4].f.lower[11] );
tran (\sa_count[4][12] , \sa_count[4].r.part0[12] );
tran (\sa_count[4][12] , \sa_count[4].f.lower[12] );
tran (\sa_count[4][13] , \sa_count[4].r.part0[13] );
tran (\sa_count[4][13] , \sa_count[4].f.lower[13] );
tran (\sa_count[4][14] , \sa_count[4].r.part0[14] );
tran (\sa_count[4][14] , \sa_count[4].f.lower[14] );
tran (\sa_count[4][15] , \sa_count[4].r.part0[15] );
tran (\sa_count[4][15] , \sa_count[4].f.lower[15] );
tran (\sa_count[4][16] , \sa_count[4].r.part0[16] );
tran (\sa_count[4][16] , \sa_count[4].f.lower[16] );
tran (\sa_count[4][17] , \sa_count[4].r.part0[17] );
tran (\sa_count[4][17] , \sa_count[4].f.lower[17] );
tran (\sa_count[4][18] , \sa_count[4].r.part0[18] );
tran (\sa_count[4][18] , \sa_count[4].f.lower[18] );
tran (\sa_count[4][19] , \sa_count[4].r.part0[19] );
tran (\sa_count[4][19] , \sa_count[4].f.lower[19] );
tran (\sa_count[4][20] , \sa_count[4].r.part0[20] );
tran (\sa_count[4][20] , \sa_count[4].f.lower[20] );
tran (\sa_count[4][21] , \sa_count[4].r.part0[21] );
tran (\sa_count[4][21] , \sa_count[4].f.lower[21] );
tran (\sa_count[4][22] , \sa_count[4].r.part0[22] );
tran (\sa_count[4][22] , \sa_count[4].f.lower[22] );
tran (\sa_count[4][23] , \sa_count[4].r.part0[23] );
tran (\sa_count[4][23] , \sa_count[4].f.lower[23] );
tran (\sa_count[4][24] , \sa_count[4].r.part0[24] );
tran (\sa_count[4][24] , \sa_count[4].f.lower[24] );
tran (\sa_count[4][25] , \sa_count[4].r.part0[25] );
tran (\sa_count[4][25] , \sa_count[4].f.lower[25] );
tran (\sa_count[4][26] , \sa_count[4].r.part0[26] );
tran (\sa_count[4][26] , \sa_count[4].f.lower[26] );
tran (\sa_count[4][27] , \sa_count[4].r.part0[27] );
tran (\sa_count[4][27] , \sa_count[4].f.lower[27] );
tran (\sa_count[4][28] , \sa_count[4].r.part0[28] );
tran (\sa_count[4][28] , \sa_count[4].f.lower[28] );
tran (\sa_count[4][29] , \sa_count[4].r.part0[29] );
tran (\sa_count[4][29] , \sa_count[4].f.lower[29] );
tran (\sa_count[4][30] , \sa_count[4].r.part0[30] );
tran (\sa_count[4][30] , \sa_count[4].f.lower[30] );
tran (\sa_count[4][31] , \sa_count[4].r.part0[31] );
tran (\sa_count[4][31] , \sa_count[4].f.lower[31] );
tran (\sa_count[4][32] , \sa_count[4].r.part1[0] );
tran (\sa_count[4][32] , \sa_count[4].f.upper[0] );
tran (\sa_count[4][33] , \sa_count[4].r.part1[1] );
tran (\sa_count[4][33] , \sa_count[4].f.upper[1] );
tran (\sa_count[4][34] , \sa_count[4].r.part1[2] );
tran (\sa_count[4][34] , \sa_count[4].f.upper[2] );
tran (\sa_count[4][35] , \sa_count[4].r.part1[3] );
tran (\sa_count[4][35] , \sa_count[4].f.upper[3] );
tran (\sa_count[4][36] , \sa_count[4].r.part1[4] );
tran (\sa_count[4][36] , \sa_count[4].f.upper[4] );
tran (\sa_count[4][37] , \sa_count[4].r.part1[5] );
tran (\sa_count[4][37] , \sa_count[4].f.upper[5] );
tran (\sa_count[4][38] , \sa_count[4].r.part1[6] );
tran (\sa_count[4][38] , \sa_count[4].f.upper[6] );
tran (\sa_count[4][39] , \sa_count[4].r.part1[7] );
tran (\sa_count[4][39] , \sa_count[4].f.upper[7] );
tran (\sa_count[4][40] , \sa_count[4].r.part1[8] );
tran (\sa_count[4][40] , \sa_count[4].f.upper[8] );
tran (\sa_count[4][41] , \sa_count[4].r.part1[9] );
tran (\sa_count[4][41] , \sa_count[4].f.upper[9] );
tran (\sa_count[4][42] , \sa_count[4].r.part1[10] );
tran (\sa_count[4][42] , \sa_count[4].f.upper[10] );
tran (\sa_count[4][43] , \sa_count[4].r.part1[11] );
tran (\sa_count[4][43] , \sa_count[4].f.upper[11] );
tran (\sa_count[4][44] , \sa_count[4].r.part1[12] );
tran (\sa_count[4][44] , \sa_count[4].f.upper[12] );
tran (\sa_count[4][45] , \sa_count[4].r.part1[13] );
tran (\sa_count[4][45] , \sa_count[4].f.upper[13] );
tran (\sa_count[4][46] , \sa_count[4].r.part1[14] );
tran (\sa_count[4][46] , \sa_count[4].f.upper[14] );
tran (\sa_count[4][47] , \sa_count[4].r.part1[15] );
tran (\sa_count[4][47] , \sa_count[4].f.upper[15] );
tran (\sa_count[4][48] , \sa_count[4].r.part1[16] );
tran (\sa_count[4][48] , \sa_count[4].f.upper[16] );
tran (\sa_count[4][49] , \sa_count[4].r.part1[17] );
tran (\sa_count[4][49] , \sa_count[4].f.upper[17] );
tran (\sa_count[4][50] , \sa_count[4].r.part1[18] );
tran (\sa_count[4][50] , \sa_count[4].f.unused[0] );
tran (\sa_count[4][51] , \sa_count[4].r.part1[19] );
tran (\sa_count[4][51] , \sa_count[4].f.unused[1] );
tran (\sa_count[4][52] , \sa_count[4].r.part1[20] );
tran (\sa_count[4][52] , \sa_count[4].f.unused[2] );
tran (\sa_count[4][53] , \sa_count[4].r.part1[21] );
tran (\sa_count[4][53] , \sa_count[4].f.unused[3] );
tran (\sa_count[4][54] , \sa_count[4].r.part1[22] );
tran (\sa_count[4][54] , \sa_count[4].f.unused[4] );
tran (\sa_count[4][55] , \sa_count[4].r.part1[23] );
tran (\sa_count[4][55] , \sa_count[4].f.unused[5] );
tran (\sa_count[4][56] , \sa_count[4].r.part1[24] );
tran (\sa_count[4][56] , \sa_count[4].f.unused[6] );
tran (\sa_count[4][57] , \sa_count[4].r.part1[25] );
tran (\sa_count[4][57] , \sa_count[4].f.unused[7] );
tran (\sa_count[4][58] , \sa_count[4].r.part1[26] );
tran (\sa_count[4][58] , \sa_count[4].f.unused[8] );
tran (\sa_count[4][59] , \sa_count[4].r.part1[27] );
tran (\sa_count[4][59] , \sa_count[4].f.unused[9] );
tran (\sa_count[4][60] , \sa_count[4].r.part1[28] );
tran (\sa_count[4][60] , \sa_count[4].f.unused[10] );
tran (\sa_count[4][61] , \sa_count[4].r.part1[29] );
tran (\sa_count[4][61] , \sa_count[4].f.unused[11] );
tran (\sa_count[4][62] , \sa_count[4].r.part1[30] );
tran (\sa_count[4][62] , \sa_count[4].f.unused[12] );
tran (\sa_count[4][63] , \sa_count[4].r.part1[31] );
tran (\sa_count[4][63] , \sa_count[4].f.unused[13] );
tran (\sa_count[5][0] , \sa_count[5].r.part0[0] );
tran (\sa_count[5][0] , \sa_count[5].f.lower[0] );
tran (\sa_count[5][1] , \sa_count[5].r.part0[1] );
tran (\sa_count[5][1] , \sa_count[5].f.lower[1] );
tran (\sa_count[5][2] , \sa_count[5].r.part0[2] );
tran (\sa_count[5][2] , \sa_count[5].f.lower[2] );
tran (\sa_count[5][3] , \sa_count[5].r.part0[3] );
tran (\sa_count[5][3] , \sa_count[5].f.lower[3] );
tran (\sa_count[5][4] , \sa_count[5].r.part0[4] );
tran (\sa_count[5][4] , \sa_count[5].f.lower[4] );
tran (\sa_count[5][5] , \sa_count[5].r.part0[5] );
tran (\sa_count[5][5] , \sa_count[5].f.lower[5] );
tran (\sa_count[5][6] , \sa_count[5].r.part0[6] );
tran (\sa_count[5][6] , \sa_count[5].f.lower[6] );
tran (\sa_count[5][7] , \sa_count[5].r.part0[7] );
tran (\sa_count[5][7] , \sa_count[5].f.lower[7] );
tran (\sa_count[5][8] , \sa_count[5].r.part0[8] );
tran (\sa_count[5][8] , \sa_count[5].f.lower[8] );
tran (\sa_count[5][9] , \sa_count[5].r.part0[9] );
tran (\sa_count[5][9] , \sa_count[5].f.lower[9] );
tran (\sa_count[5][10] , \sa_count[5].r.part0[10] );
tran (\sa_count[5][10] , \sa_count[5].f.lower[10] );
tran (\sa_count[5][11] , \sa_count[5].r.part0[11] );
tran (\sa_count[5][11] , \sa_count[5].f.lower[11] );
tran (\sa_count[5][12] , \sa_count[5].r.part0[12] );
tran (\sa_count[5][12] , \sa_count[5].f.lower[12] );
tran (\sa_count[5][13] , \sa_count[5].r.part0[13] );
tran (\sa_count[5][13] , \sa_count[5].f.lower[13] );
tran (\sa_count[5][14] , \sa_count[5].r.part0[14] );
tran (\sa_count[5][14] , \sa_count[5].f.lower[14] );
tran (\sa_count[5][15] , \sa_count[5].r.part0[15] );
tran (\sa_count[5][15] , \sa_count[5].f.lower[15] );
tran (\sa_count[5][16] , \sa_count[5].r.part0[16] );
tran (\sa_count[5][16] , \sa_count[5].f.lower[16] );
tran (\sa_count[5][17] , \sa_count[5].r.part0[17] );
tran (\sa_count[5][17] , \sa_count[5].f.lower[17] );
tran (\sa_count[5][18] , \sa_count[5].r.part0[18] );
tran (\sa_count[5][18] , \sa_count[5].f.lower[18] );
tran (\sa_count[5][19] , \sa_count[5].r.part0[19] );
tran (\sa_count[5][19] , \sa_count[5].f.lower[19] );
tran (\sa_count[5][20] , \sa_count[5].r.part0[20] );
tran (\sa_count[5][20] , \sa_count[5].f.lower[20] );
tran (\sa_count[5][21] , \sa_count[5].r.part0[21] );
tran (\sa_count[5][21] , \sa_count[5].f.lower[21] );
tran (\sa_count[5][22] , \sa_count[5].r.part0[22] );
tran (\sa_count[5][22] , \sa_count[5].f.lower[22] );
tran (\sa_count[5][23] , \sa_count[5].r.part0[23] );
tran (\sa_count[5][23] , \sa_count[5].f.lower[23] );
tran (\sa_count[5][24] , \sa_count[5].r.part0[24] );
tran (\sa_count[5][24] , \sa_count[5].f.lower[24] );
tran (\sa_count[5][25] , \sa_count[5].r.part0[25] );
tran (\sa_count[5][25] , \sa_count[5].f.lower[25] );
tran (\sa_count[5][26] , \sa_count[5].r.part0[26] );
tran (\sa_count[5][26] , \sa_count[5].f.lower[26] );
tran (\sa_count[5][27] , \sa_count[5].r.part0[27] );
tran (\sa_count[5][27] , \sa_count[5].f.lower[27] );
tran (\sa_count[5][28] , \sa_count[5].r.part0[28] );
tran (\sa_count[5][28] , \sa_count[5].f.lower[28] );
tran (\sa_count[5][29] , \sa_count[5].r.part0[29] );
tran (\sa_count[5][29] , \sa_count[5].f.lower[29] );
tran (\sa_count[5][30] , \sa_count[5].r.part0[30] );
tran (\sa_count[5][30] , \sa_count[5].f.lower[30] );
tran (\sa_count[5][31] , \sa_count[5].r.part0[31] );
tran (\sa_count[5][31] , \sa_count[5].f.lower[31] );
tran (\sa_count[5][32] , \sa_count[5].r.part1[0] );
tran (\sa_count[5][32] , \sa_count[5].f.upper[0] );
tran (\sa_count[5][33] , \sa_count[5].r.part1[1] );
tran (\sa_count[5][33] , \sa_count[5].f.upper[1] );
tran (\sa_count[5][34] , \sa_count[5].r.part1[2] );
tran (\sa_count[5][34] , \sa_count[5].f.upper[2] );
tran (\sa_count[5][35] , \sa_count[5].r.part1[3] );
tran (\sa_count[5][35] , \sa_count[5].f.upper[3] );
tran (\sa_count[5][36] , \sa_count[5].r.part1[4] );
tran (\sa_count[5][36] , \sa_count[5].f.upper[4] );
tran (\sa_count[5][37] , \sa_count[5].r.part1[5] );
tran (\sa_count[5][37] , \sa_count[5].f.upper[5] );
tran (\sa_count[5][38] , \sa_count[5].r.part1[6] );
tran (\sa_count[5][38] , \sa_count[5].f.upper[6] );
tran (\sa_count[5][39] , \sa_count[5].r.part1[7] );
tran (\sa_count[5][39] , \sa_count[5].f.upper[7] );
tran (\sa_count[5][40] , \sa_count[5].r.part1[8] );
tran (\sa_count[5][40] , \sa_count[5].f.upper[8] );
tran (\sa_count[5][41] , \sa_count[5].r.part1[9] );
tran (\sa_count[5][41] , \sa_count[5].f.upper[9] );
tran (\sa_count[5][42] , \sa_count[5].r.part1[10] );
tran (\sa_count[5][42] , \sa_count[5].f.upper[10] );
tran (\sa_count[5][43] , \sa_count[5].r.part1[11] );
tran (\sa_count[5][43] , \sa_count[5].f.upper[11] );
tran (\sa_count[5][44] , \sa_count[5].r.part1[12] );
tran (\sa_count[5][44] , \sa_count[5].f.upper[12] );
tran (\sa_count[5][45] , \sa_count[5].r.part1[13] );
tran (\sa_count[5][45] , \sa_count[5].f.upper[13] );
tran (\sa_count[5][46] , \sa_count[5].r.part1[14] );
tran (\sa_count[5][46] , \sa_count[5].f.upper[14] );
tran (\sa_count[5][47] , \sa_count[5].r.part1[15] );
tran (\sa_count[5][47] , \sa_count[5].f.upper[15] );
tran (\sa_count[5][48] , \sa_count[5].r.part1[16] );
tran (\sa_count[5][48] , \sa_count[5].f.upper[16] );
tran (\sa_count[5][49] , \sa_count[5].r.part1[17] );
tran (\sa_count[5][49] , \sa_count[5].f.upper[17] );
tran (\sa_count[5][50] , \sa_count[5].r.part1[18] );
tran (\sa_count[5][50] , \sa_count[5].f.unused[0] );
tran (\sa_count[5][51] , \sa_count[5].r.part1[19] );
tran (\sa_count[5][51] , \sa_count[5].f.unused[1] );
tran (\sa_count[5][52] , \sa_count[5].r.part1[20] );
tran (\sa_count[5][52] , \sa_count[5].f.unused[2] );
tran (\sa_count[5][53] , \sa_count[5].r.part1[21] );
tran (\sa_count[5][53] , \sa_count[5].f.unused[3] );
tran (\sa_count[5][54] , \sa_count[5].r.part1[22] );
tran (\sa_count[5][54] , \sa_count[5].f.unused[4] );
tran (\sa_count[5][55] , \sa_count[5].r.part1[23] );
tran (\sa_count[5][55] , \sa_count[5].f.unused[5] );
tran (\sa_count[5][56] , \sa_count[5].r.part1[24] );
tran (\sa_count[5][56] , \sa_count[5].f.unused[6] );
tran (\sa_count[5][57] , \sa_count[5].r.part1[25] );
tran (\sa_count[5][57] , \sa_count[5].f.unused[7] );
tran (\sa_count[5][58] , \sa_count[5].r.part1[26] );
tran (\sa_count[5][58] , \sa_count[5].f.unused[8] );
tran (\sa_count[5][59] , \sa_count[5].r.part1[27] );
tran (\sa_count[5][59] , \sa_count[5].f.unused[9] );
tran (\sa_count[5][60] , \sa_count[5].r.part1[28] );
tran (\sa_count[5][60] , \sa_count[5].f.unused[10] );
tran (\sa_count[5][61] , \sa_count[5].r.part1[29] );
tran (\sa_count[5][61] , \sa_count[5].f.unused[11] );
tran (\sa_count[5][62] , \sa_count[5].r.part1[30] );
tran (\sa_count[5][62] , \sa_count[5].f.unused[12] );
tran (\sa_count[5][63] , \sa_count[5].r.part1[31] );
tran (\sa_count[5][63] , \sa_count[5].f.unused[13] );
tran (\sa_count[6][0] , \sa_count[6].r.part0[0] );
tran (\sa_count[6][0] , \sa_count[6].f.lower[0] );
tran (\sa_count[6][1] , \sa_count[6].r.part0[1] );
tran (\sa_count[6][1] , \sa_count[6].f.lower[1] );
tran (\sa_count[6][2] , \sa_count[6].r.part0[2] );
tran (\sa_count[6][2] , \sa_count[6].f.lower[2] );
tran (\sa_count[6][3] , \sa_count[6].r.part0[3] );
tran (\sa_count[6][3] , \sa_count[6].f.lower[3] );
tran (\sa_count[6][4] , \sa_count[6].r.part0[4] );
tran (\sa_count[6][4] , \sa_count[6].f.lower[4] );
tran (\sa_count[6][5] , \sa_count[6].r.part0[5] );
tran (\sa_count[6][5] , \sa_count[6].f.lower[5] );
tran (\sa_count[6][6] , \sa_count[6].r.part0[6] );
tran (\sa_count[6][6] , \sa_count[6].f.lower[6] );
tran (\sa_count[6][7] , \sa_count[6].r.part0[7] );
tran (\sa_count[6][7] , \sa_count[6].f.lower[7] );
tran (\sa_count[6][8] , \sa_count[6].r.part0[8] );
tran (\sa_count[6][8] , \sa_count[6].f.lower[8] );
tran (\sa_count[6][9] , \sa_count[6].r.part0[9] );
tran (\sa_count[6][9] , \sa_count[6].f.lower[9] );
tran (\sa_count[6][10] , \sa_count[6].r.part0[10] );
tran (\sa_count[6][10] , \sa_count[6].f.lower[10] );
tran (\sa_count[6][11] , \sa_count[6].r.part0[11] );
tran (\sa_count[6][11] , \sa_count[6].f.lower[11] );
tran (\sa_count[6][12] , \sa_count[6].r.part0[12] );
tran (\sa_count[6][12] , \sa_count[6].f.lower[12] );
tran (\sa_count[6][13] , \sa_count[6].r.part0[13] );
tran (\sa_count[6][13] , \sa_count[6].f.lower[13] );
tran (\sa_count[6][14] , \sa_count[6].r.part0[14] );
tran (\sa_count[6][14] , \sa_count[6].f.lower[14] );
tran (\sa_count[6][15] , \sa_count[6].r.part0[15] );
tran (\sa_count[6][15] , \sa_count[6].f.lower[15] );
tran (\sa_count[6][16] , \sa_count[6].r.part0[16] );
tran (\sa_count[6][16] , \sa_count[6].f.lower[16] );
tran (\sa_count[6][17] , \sa_count[6].r.part0[17] );
tran (\sa_count[6][17] , \sa_count[6].f.lower[17] );
tran (\sa_count[6][18] , \sa_count[6].r.part0[18] );
tran (\sa_count[6][18] , \sa_count[6].f.lower[18] );
tran (\sa_count[6][19] , \sa_count[6].r.part0[19] );
tran (\sa_count[6][19] , \sa_count[6].f.lower[19] );
tran (\sa_count[6][20] , \sa_count[6].r.part0[20] );
tran (\sa_count[6][20] , \sa_count[6].f.lower[20] );
tran (\sa_count[6][21] , \sa_count[6].r.part0[21] );
tran (\sa_count[6][21] , \sa_count[6].f.lower[21] );
tran (\sa_count[6][22] , \sa_count[6].r.part0[22] );
tran (\sa_count[6][22] , \sa_count[6].f.lower[22] );
tran (\sa_count[6][23] , \sa_count[6].r.part0[23] );
tran (\sa_count[6][23] , \sa_count[6].f.lower[23] );
tran (\sa_count[6][24] , \sa_count[6].r.part0[24] );
tran (\sa_count[6][24] , \sa_count[6].f.lower[24] );
tran (\sa_count[6][25] , \sa_count[6].r.part0[25] );
tran (\sa_count[6][25] , \sa_count[6].f.lower[25] );
tran (\sa_count[6][26] , \sa_count[6].r.part0[26] );
tran (\sa_count[6][26] , \sa_count[6].f.lower[26] );
tran (\sa_count[6][27] , \sa_count[6].r.part0[27] );
tran (\sa_count[6][27] , \sa_count[6].f.lower[27] );
tran (\sa_count[6][28] , \sa_count[6].r.part0[28] );
tran (\sa_count[6][28] , \sa_count[6].f.lower[28] );
tran (\sa_count[6][29] , \sa_count[6].r.part0[29] );
tran (\sa_count[6][29] , \sa_count[6].f.lower[29] );
tran (\sa_count[6][30] , \sa_count[6].r.part0[30] );
tran (\sa_count[6][30] , \sa_count[6].f.lower[30] );
tran (\sa_count[6][31] , \sa_count[6].r.part0[31] );
tran (\sa_count[6][31] , \sa_count[6].f.lower[31] );
tran (\sa_count[6][32] , \sa_count[6].r.part1[0] );
tran (\sa_count[6][32] , \sa_count[6].f.upper[0] );
tran (\sa_count[6][33] , \sa_count[6].r.part1[1] );
tran (\sa_count[6][33] , \sa_count[6].f.upper[1] );
tran (\sa_count[6][34] , \sa_count[6].r.part1[2] );
tran (\sa_count[6][34] , \sa_count[6].f.upper[2] );
tran (\sa_count[6][35] , \sa_count[6].r.part1[3] );
tran (\sa_count[6][35] , \sa_count[6].f.upper[3] );
tran (\sa_count[6][36] , \sa_count[6].r.part1[4] );
tran (\sa_count[6][36] , \sa_count[6].f.upper[4] );
tran (\sa_count[6][37] , \sa_count[6].r.part1[5] );
tran (\sa_count[6][37] , \sa_count[6].f.upper[5] );
tran (\sa_count[6][38] , \sa_count[6].r.part1[6] );
tran (\sa_count[6][38] , \sa_count[6].f.upper[6] );
tran (\sa_count[6][39] , \sa_count[6].r.part1[7] );
tran (\sa_count[6][39] , \sa_count[6].f.upper[7] );
tran (\sa_count[6][40] , \sa_count[6].r.part1[8] );
tran (\sa_count[6][40] , \sa_count[6].f.upper[8] );
tran (\sa_count[6][41] , \sa_count[6].r.part1[9] );
tran (\sa_count[6][41] , \sa_count[6].f.upper[9] );
tran (\sa_count[6][42] , \sa_count[6].r.part1[10] );
tran (\sa_count[6][42] , \sa_count[6].f.upper[10] );
tran (\sa_count[6][43] , \sa_count[6].r.part1[11] );
tran (\sa_count[6][43] , \sa_count[6].f.upper[11] );
tran (\sa_count[6][44] , \sa_count[6].r.part1[12] );
tran (\sa_count[6][44] , \sa_count[6].f.upper[12] );
tran (\sa_count[6][45] , \sa_count[6].r.part1[13] );
tran (\sa_count[6][45] , \sa_count[6].f.upper[13] );
tran (\sa_count[6][46] , \sa_count[6].r.part1[14] );
tran (\sa_count[6][46] , \sa_count[6].f.upper[14] );
tran (\sa_count[6][47] , \sa_count[6].r.part1[15] );
tran (\sa_count[6][47] , \sa_count[6].f.upper[15] );
tran (\sa_count[6][48] , \sa_count[6].r.part1[16] );
tran (\sa_count[6][48] , \sa_count[6].f.upper[16] );
tran (\sa_count[6][49] , \sa_count[6].r.part1[17] );
tran (\sa_count[6][49] , \sa_count[6].f.upper[17] );
tran (\sa_count[6][50] , \sa_count[6].r.part1[18] );
tran (\sa_count[6][50] , \sa_count[6].f.unused[0] );
tran (\sa_count[6][51] , \sa_count[6].r.part1[19] );
tran (\sa_count[6][51] , \sa_count[6].f.unused[1] );
tran (\sa_count[6][52] , \sa_count[6].r.part1[20] );
tran (\sa_count[6][52] , \sa_count[6].f.unused[2] );
tran (\sa_count[6][53] , \sa_count[6].r.part1[21] );
tran (\sa_count[6][53] , \sa_count[6].f.unused[3] );
tran (\sa_count[6][54] , \sa_count[6].r.part1[22] );
tran (\sa_count[6][54] , \sa_count[6].f.unused[4] );
tran (\sa_count[6][55] , \sa_count[6].r.part1[23] );
tran (\sa_count[6][55] , \sa_count[6].f.unused[5] );
tran (\sa_count[6][56] , \sa_count[6].r.part1[24] );
tran (\sa_count[6][56] , \sa_count[6].f.unused[6] );
tran (\sa_count[6][57] , \sa_count[6].r.part1[25] );
tran (\sa_count[6][57] , \sa_count[6].f.unused[7] );
tran (\sa_count[6][58] , \sa_count[6].r.part1[26] );
tran (\sa_count[6][58] , \sa_count[6].f.unused[8] );
tran (\sa_count[6][59] , \sa_count[6].r.part1[27] );
tran (\sa_count[6][59] , \sa_count[6].f.unused[9] );
tran (\sa_count[6][60] , \sa_count[6].r.part1[28] );
tran (\sa_count[6][60] , \sa_count[6].f.unused[10] );
tran (\sa_count[6][61] , \sa_count[6].r.part1[29] );
tran (\sa_count[6][61] , \sa_count[6].f.unused[11] );
tran (\sa_count[6][62] , \sa_count[6].r.part1[30] );
tran (\sa_count[6][62] , \sa_count[6].f.unused[12] );
tran (\sa_count[6][63] , \sa_count[6].r.part1[31] );
tran (\sa_count[6][63] , \sa_count[6].f.unused[13] );
tran (\sa_count[7][0] , \sa_count[7].r.part0[0] );
tran (\sa_count[7][0] , \sa_count[7].f.lower[0] );
tran (\sa_count[7][1] , \sa_count[7].r.part0[1] );
tran (\sa_count[7][1] , \sa_count[7].f.lower[1] );
tran (\sa_count[7][2] , \sa_count[7].r.part0[2] );
tran (\sa_count[7][2] , \sa_count[7].f.lower[2] );
tran (\sa_count[7][3] , \sa_count[7].r.part0[3] );
tran (\sa_count[7][3] , \sa_count[7].f.lower[3] );
tran (\sa_count[7][4] , \sa_count[7].r.part0[4] );
tran (\sa_count[7][4] , \sa_count[7].f.lower[4] );
tran (\sa_count[7][5] , \sa_count[7].r.part0[5] );
tran (\sa_count[7][5] , \sa_count[7].f.lower[5] );
tran (\sa_count[7][6] , \sa_count[7].r.part0[6] );
tran (\sa_count[7][6] , \sa_count[7].f.lower[6] );
tran (\sa_count[7][7] , \sa_count[7].r.part0[7] );
tran (\sa_count[7][7] , \sa_count[7].f.lower[7] );
tran (\sa_count[7][8] , \sa_count[7].r.part0[8] );
tran (\sa_count[7][8] , \sa_count[7].f.lower[8] );
tran (\sa_count[7][9] , \sa_count[7].r.part0[9] );
tran (\sa_count[7][9] , \sa_count[7].f.lower[9] );
tran (\sa_count[7][10] , \sa_count[7].r.part0[10] );
tran (\sa_count[7][10] , \sa_count[7].f.lower[10] );
tran (\sa_count[7][11] , \sa_count[7].r.part0[11] );
tran (\sa_count[7][11] , \sa_count[7].f.lower[11] );
tran (\sa_count[7][12] , \sa_count[7].r.part0[12] );
tran (\sa_count[7][12] , \sa_count[7].f.lower[12] );
tran (\sa_count[7][13] , \sa_count[7].r.part0[13] );
tran (\sa_count[7][13] , \sa_count[7].f.lower[13] );
tran (\sa_count[7][14] , \sa_count[7].r.part0[14] );
tran (\sa_count[7][14] , \sa_count[7].f.lower[14] );
tran (\sa_count[7][15] , \sa_count[7].r.part0[15] );
tran (\sa_count[7][15] , \sa_count[7].f.lower[15] );
tran (\sa_count[7][16] , \sa_count[7].r.part0[16] );
tran (\sa_count[7][16] , \sa_count[7].f.lower[16] );
tran (\sa_count[7][17] , \sa_count[7].r.part0[17] );
tran (\sa_count[7][17] , \sa_count[7].f.lower[17] );
tran (\sa_count[7][18] , \sa_count[7].r.part0[18] );
tran (\sa_count[7][18] , \sa_count[7].f.lower[18] );
tran (\sa_count[7][19] , \sa_count[7].r.part0[19] );
tran (\sa_count[7][19] , \sa_count[7].f.lower[19] );
tran (\sa_count[7][20] , \sa_count[7].r.part0[20] );
tran (\sa_count[7][20] , \sa_count[7].f.lower[20] );
tran (\sa_count[7][21] , \sa_count[7].r.part0[21] );
tran (\sa_count[7][21] , \sa_count[7].f.lower[21] );
tran (\sa_count[7][22] , \sa_count[7].r.part0[22] );
tran (\sa_count[7][22] , \sa_count[7].f.lower[22] );
tran (\sa_count[7][23] , \sa_count[7].r.part0[23] );
tran (\sa_count[7][23] , \sa_count[7].f.lower[23] );
tran (\sa_count[7][24] , \sa_count[7].r.part0[24] );
tran (\sa_count[7][24] , \sa_count[7].f.lower[24] );
tran (\sa_count[7][25] , \sa_count[7].r.part0[25] );
tran (\sa_count[7][25] , \sa_count[7].f.lower[25] );
tran (\sa_count[7][26] , \sa_count[7].r.part0[26] );
tran (\sa_count[7][26] , \sa_count[7].f.lower[26] );
tran (\sa_count[7][27] , \sa_count[7].r.part0[27] );
tran (\sa_count[7][27] , \sa_count[7].f.lower[27] );
tran (\sa_count[7][28] , \sa_count[7].r.part0[28] );
tran (\sa_count[7][28] , \sa_count[7].f.lower[28] );
tran (\sa_count[7][29] , \sa_count[7].r.part0[29] );
tran (\sa_count[7][29] , \sa_count[7].f.lower[29] );
tran (\sa_count[7][30] , \sa_count[7].r.part0[30] );
tran (\sa_count[7][30] , \sa_count[7].f.lower[30] );
tran (\sa_count[7][31] , \sa_count[7].r.part0[31] );
tran (\sa_count[7][31] , \sa_count[7].f.lower[31] );
tran (\sa_count[7][32] , \sa_count[7].r.part1[0] );
tran (\sa_count[7][32] , \sa_count[7].f.upper[0] );
tran (\sa_count[7][33] , \sa_count[7].r.part1[1] );
tran (\sa_count[7][33] , \sa_count[7].f.upper[1] );
tran (\sa_count[7][34] , \sa_count[7].r.part1[2] );
tran (\sa_count[7][34] , \sa_count[7].f.upper[2] );
tran (\sa_count[7][35] , \sa_count[7].r.part1[3] );
tran (\sa_count[7][35] , \sa_count[7].f.upper[3] );
tran (\sa_count[7][36] , \sa_count[7].r.part1[4] );
tran (\sa_count[7][36] , \sa_count[7].f.upper[4] );
tran (\sa_count[7][37] , \sa_count[7].r.part1[5] );
tran (\sa_count[7][37] , \sa_count[7].f.upper[5] );
tran (\sa_count[7][38] , \sa_count[7].r.part1[6] );
tran (\sa_count[7][38] , \sa_count[7].f.upper[6] );
tran (\sa_count[7][39] , \sa_count[7].r.part1[7] );
tran (\sa_count[7][39] , \sa_count[7].f.upper[7] );
tran (\sa_count[7][40] , \sa_count[7].r.part1[8] );
tran (\sa_count[7][40] , \sa_count[7].f.upper[8] );
tran (\sa_count[7][41] , \sa_count[7].r.part1[9] );
tran (\sa_count[7][41] , \sa_count[7].f.upper[9] );
tran (\sa_count[7][42] , \sa_count[7].r.part1[10] );
tran (\sa_count[7][42] , \sa_count[7].f.upper[10] );
tran (\sa_count[7][43] , \sa_count[7].r.part1[11] );
tran (\sa_count[7][43] , \sa_count[7].f.upper[11] );
tran (\sa_count[7][44] , \sa_count[7].r.part1[12] );
tran (\sa_count[7][44] , \sa_count[7].f.upper[12] );
tran (\sa_count[7][45] , \sa_count[7].r.part1[13] );
tran (\sa_count[7][45] , \sa_count[7].f.upper[13] );
tran (\sa_count[7][46] , \sa_count[7].r.part1[14] );
tran (\sa_count[7][46] , \sa_count[7].f.upper[14] );
tran (\sa_count[7][47] , \sa_count[7].r.part1[15] );
tran (\sa_count[7][47] , \sa_count[7].f.upper[15] );
tran (\sa_count[7][48] , \sa_count[7].r.part1[16] );
tran (\sa_count[7][48] , \sa_count[7].f.upper[16] );
tran (\sa_count[7][49] , \sa_count[7].r.part1[17] );
tran (\sa_count[7][49] , \sa_count[7].f.upper[17] );
tran (\sa_count[7][50] , \sa_count[7].r.part1[18] );
tran (\sa_count[7][50] , \sa_count[7].f.unused[0] );
tran (\sa_count[7][51] , \sa_count[7].r.part1[19] );
tran (\sa_count[7][51] , \sa_count[7].f.unused[1] );
tran (\sa_count[7][52] , \sa_count[7].r.part1[20] );
tran (\sa_count[7][52] , \sa_count[7].f.unused[2] );
tran (\sa_count[7][53] , \sa_count[7].r.part1[21] );
tran (\sa_count[7][53] , \sa_count[7].f.unused[3] );
tran (\sa_count[7][54] , \sa_count[7].r.part1[22] );
tran (\sa_count[7][54] , \sa_count[7].f.unused[4] );
tran (\sa_count[7][55] , \sa_count[7].r.part1[23] );
tran (\sa_count[7][55] , \sa_count[7].f.unused[5] );
tran (\sa_count[7][56] , \sa_count[7].r.part1[24] );
tran (\sa_count[7][56] , \sa_count[7].f.unused[6] );
tran (\sa_count[7][57] , \sa_count[7].r.part1[25] );
tran (\sa_count[7][57] , \sa_count[7].f.unused[7] );
tran (\sa_count[7][58] , \sa_count[7].r.part1[26] );
tran (\sa_count[7][58] , \sa_count[7].f.unused[8] );
tran (\sa_count[7][59] , \sa_count[7].r.part1[27] );
tran (\sa_count[7][59] , \sa_count[7].f.unused[9] );
tran (\sa_count[7][60] , \sa_count[7].r.part1[28] );
tran (\sa_count[7][60] , \sa_count[7].f.unused[10] );
tran (\sa_count[7][61] , \sa_count[7].r.part1[29] );
tran (\sa_count[7][61] , \sa_count[7].f.unused[11] );
tran (\sa_count[7][62] , \sa_count[7].r.part1[30] );
tran (\sa_count[7][62] , \sa_count[7].f.unused[12] );
tran (\sa_count[7][63] , \sa_count[7].r.part1[31] );
tran (\sa_count[7][63] , \sa_count[7].f.unused[13] );
tran (\sa_count[8][0] , \sa_count[8].r.part0[0] );
tran (\sa_count[8][0] , \sa_count[8].f.lower[0] );
tran (\sa_count[8][1] , \sa_count[8].r.part0[1] );
tran (\sa_count[8][1] , \sa_count[8].f.lower[1] );
tran (\sa_count[8][2] , \sa_count[8].r.part0[2] );
tran (\sa_count[8][2] , \sa_count[8].f.lower[2] );
tran (\sa_count[8][3] , \sa_count[8].r.part0[3] );
tran (\sa_count[8][3] , \sa_count[8].f.lower[3] );
tran (\sa_count[8][4] , \sa_count[8].r.part0[4] );
tran (\sa_count[8][4] , \sa_count[8].f.lower[4] );
tran (\sa_count[8][5] , \sa_count[8].r.part0[5] );
tran (\sa_count[8][5] , \sa_count[8].f.lower[5] );
tran (\sa_count[8][6] , \sa_count[8].r.part0[6] );
tran (\sa_count[8][6] , \sa_count[8].f.lower[6] );
tran (\sa_count[8][7] , \sa_count[8].r.part0[7] );
tran (\sa_count[8][7] , \sa_count[8].f.lower[7] );
tran (\sa_count[8][8] , \sa_count[8].r.part0[8] );
tran (\sa_count[8][8] , \sa_count[8].f.lower[8] );
tran (\sa_count[8][9] , \sa_count[8].r.part0[9] );
tran (\sa_count[8][9] , \sa_count[8].f.lower[9] );
tran (\sa_count[8][10] , \sa_count[8].r.part0[10] );
tran (\sa_count[8][10] , \sa_count[8].f.lower[10] );
tran (\sa_count[8][11] , \sa_count[8].r.part0[11] );
tran (\sa_count[8][11] , \sa_count[8].f.lower[11] );
tran (\sa_count[8][12] , \sa_count[8].r.part0[12] );
tran (\sa_count[8][12] , \sa_count[8].f.lower[12] );
tran (\sa_count[8][13] , \sa_count[8].r.part0[13] );
tran (\sa_count[8][13] , \sa_count[8].f.lower[13] );
tran (\sa_count[8][14] , \sa_count[8].r.part0[14] );
tran (\sa_count[8][14] , \sa_count[8].f.lower[14] );
tran (\sa_count[8][15] , \sa_count[8].r.part0[15] );
tran (\sa_count[8][15] , \sa_count[8].f.lower[15] );
tran (\sa_count[8][16] , \sa_count[8].r.part0[16] );
tran (\sa_count[8][16] , \sa_count[8].f.lower[16] );
tran (\sa_count[8][17] , \sa_count[8].r.part0[17] );
tran (\sa_count[8][17] , \sa_count[8].f.lower[17] );
tran (\sa_count[8][18] , \sa_count[8].r.part0[18] );
tran (\sa_count[8][18] , \sa_count[8].f.lower[18] );
tran (\sa_count[8][19] , \sa_count[8].r.part0[19] );
tran (\sa_count[8][19] , \sa_count[8].f.lower[19] );
tran (\sa_count[8][20] , \sa_count[8].r.part0[20] );
tran (\sa_count[8][20] , \sa_count[8].f.lower[20] );
tran (\sa_count[8][21] , \sa_count[8].r.part0[21] );
tran (\sa_count[8][21] , \sa_count[8].f.lower[21] );
tran (\sa_count[8][22] , \sa_count[8].r.part0[22] );
tran (\sa_count[8][22] , \sa_count[8].f.lower[22] );
tran (\sa_count[8][23] , \sa_count[8].r.part0[23] );
tran (\sa_count[8][23] , \sa_count[8].f.lower[23] );
tran (\sa_count[8][24] , \sa_count[8].r.part0[24] );
tran (\sa_count[8][24] , \sa_count[8].f.lower[24] );
tran (\sa_count[8][25] , \sa_count[8].r.part0[25] );
tran (\sa_count[8][25] , \sa_count[8].f.lower[25] );
tran (\sa_count[8][26] , \sa_count[8].r.part0[26] );
tran (\sa_count[8][26] , \sa_count[8].f.lower[26] );
tran (\sa_count[8][27] , \sa_count[8].r.part0[27] );
tran (\sa_count[8][27] , \sa_count[8].f.lower[27] );
tran (\sa_count[8][28] , \sa_count[8].r.part0[28] );
tran (\sa_count[8][28] , \sa_count[8].f.lower[28] );
tran (\sa_count[8][29] , \sa_count[8].r.part0[29] );
tran (\sa_count[8][29] , \sa_count[8].f.lower[29] );
tran (\sa_count[8][30] , \sa_count[8].r.part0[30] );
tran (\sa_count[8][30] , \sa_count[8].f.lower[30] );
tran (\sa_count[8][31] , \sa_count[8].r.part0[31] );
tran (\sa_count[8][31] , \sa_count[8].f.lower[31] );
tran (\sa_count[8][32] , \sa_count[8].r.part1[0] );
tran (\sa_count[8][32] , \sa_count[8].f.upper[0] );
tran (\sa_count[8][33] , \sa_count[8].r.part1[1] );
tran (\sa_count[8][33] , \sa_count[8].f.upper[1] );
tran (\sa_count[8][34] , \sa_count[8].r.part1[2] );
tran (\sa_count[8][34] , \sa_count[8].f.upper[2] );
tran (\sa_count[8][35] , \sa_count[8].r.part1[3] );
tran (\sa_count[8][35] , \sa_count[8].f.upper[3] );
tran (\sa_count[8][36] , \sa_count[8].r.part1[4] );
tran (\sa_count[8][36] , \sa_count[8].f.upper[4] );
tran (\sa_count[8][37] , \sa_count[8].r.part1[5] );
tran (\sa_count[8][37] , \sa_count[8].f.upper[5] );
tran (\sa_count[8][38] , \sa_count[8].r.part1[6] );
tran (\sa_count[8][38] , \sa_count[8].f.upper[6] );
tran (\sa_count[8][39] , \sa_count[8].r.part1[7] );
tran (\sa_count[8][39] , \sa_count[8].f.upper[7] );
tran (\sa_count[8][40] , \sa_count[8].r.part1[8] );
tran (\sa_count[8][40] , \sa_count[8].f.upper[8] );
tran (\sa_count[8][41] , \sa_count[8].r.part1[9] );
tran (\sa_count[8][41] , \sa_count[8].f.upper[9] );
tran (\sa_count[8][42] , \sa_count[8].r.part1[10] );
tran (\sa_count[8][42] , \sa_count[8].f.upper[10] );
tran (\sa_count[8][43] , \sa_count[8].r.part1[11] );
tran (\sa_count[8][43] , \sa_count[8].f.upper[11] );
tran (\sa_count[8][44] , \sa_count[8].r.part1[12] );
tran (\sa_count[8][44] , \sa_count[8].f.upper[12] );
tran (\sa_count[8][45] , \sa_count[8].r.part1[13] );
tran (\sa_count[8][45] , \sa_count[8].f.upper[13] );
tran (\sa_count[8][46] , \sa_count[8].r.part1[14] );
tran (\sa_count[8][46] , \sa_count[8].f.upper[14] );
tran (\sa_count[8][47] , \sa_count[8].r.part1[15] );
tran (\sa_count[8][47] , \sa_count[8].f.upper[15] );
tran (\sa_count[8][48] , \sa_count[8].r.part1[16] );
tran (\sa_count[8][48] , \sa_count[8].f.upper[16] );
tran (\sa_count[8][49] , \sa_count[8].r.part1[17] );
tran (\sa_count[8][49] , \sa_count[8].f.upper[17] );
tran (\sa_count[8][50] , \sa_count[8].r.part1[18] );
tran (\sa_count[8][50] , \sa_count[8].f.unused[0] );
tran (\sa_count[8][51] , \sa_count[8].r.part1[19] );
tran (\sa_count[8][51] , \sa_count[8].f.unused[1] );
tran (\sa_count[8][52] , \sa_count[8].r.part1[20] );
tran (\sa_count[8][52] , \sa_count[8].f.unused[2] );
tran (\sa_count[8][53] , \sa_count[8].r.part1[21] );
tran (\sa_count[8][53] , \sa_count[8].f.unused[3] );
tran (\sa_count[8][54] , \sa_count[8].r.part1[22] );
tran (\sa_count[8][54] , \sa_count[8].f.unused[4] );
tran (\sa_count[8][55] , \sa_count[8].r.part1[23] );
tran (\sa_count[8][55] , \sa_count[8].f.unused[5] );
tran (\sa_count[8][56] , \sa_count[8].r.part1[24] );
tran (\sa_count[8][56] , \sa_count[8].f.unused[6] );
tran (\sa_count[8][57] , \sa_count[8].r.part1[25] );
tran (\sa_count[8][57] , \sa_count[8].f.unused[7] );
tran (\sa_count[8][58] , \sa_count[8].r.part1[26] );
tran (\sa_count[8][58] , \sa_count[8].f.unused[8] );
tran (\sa_count[8][59] , \sa_count[8].r.part1[27] );
tran (\sa_count[8][59] , \sa_count[8].f.unused[9] );
tran (\sa_count[8][60] , \sa_count[8].r.part1[28] );
tran (\sa_count[8][60] , \sa_count[8].f.unused[10] );
tran (\sa_count[8][61] , \sa_count[8].r.part1[29] );
tran (\sa_count[8][61] , \sa_count[8].f.unused[11] );
tran (\sa_count[8][62] , \sa_count[8].r.part1[30] );
tran (\sa_count[8][62] , \sa_count[8].f.unused[12] );
tran (\sa_count[8][63] , \sa_count[8].r.part1[31] );
tran (\sa_count[8][63] , \sa_count[8].f.unused[13] );
tran (\sa_count[9][0] , \sa_count[9].r.part0[0] );
tran (\sa_count[9][0] , \sa_count[9].f.lower[0] );
tran (\sa_count[9][1] , \sa_count[9].r.part0[1] );
tran (\sa_count[9][1] , \sa_count[9].f.lower[1] );
tran (\sa_count[9][2] , \sa_count[9].r.part0[2] );
tran (\sa_count[9][2] , \sa_count[9].f.lower[2] );
tran (\sa_count[9][3] , \sa_count[9].r.part0[3] );
tran (\sa_count[9][3] , \sa_count[9].f.lower[3] );
tran (\sa_count[9][4] , \sa_count[9].r.part0[4] );
tran (\sa_count[9][4] , \sa_count[9].f.lower[4] );
tran (\sa_count[9][5] , \sa_count[9].r.part0[5] );
tran (\sa_count[9][5] , \sa_count[9].f.lower[5] );
tran (\sa_count[9][6] , \sa_count[9].r.part0[6] );
tran (\sa_count[9][6] , \sa_count[9].f.lower[6] );
tran (\sa_count[9][7] , \sa_count[9].r.part0[7] );
tran (\sa_count[9][7] , \sa_count[9].f.lower[7] );
tran (\sa_count[9][8] , \sa_count[9].r.part0[8] );
tran (\sa_count[9][8] , \sa_count[9].f.lower[8] );
tran (\sa_count[9][9] , \sa_count[9].r.part0[9] );
tran (\sa_count[9][9] , \sa_count[9].f.lower[9] );
tran (\sa_count[9][10] , \sa_count[9].r.part0[10] );
tran (\sa_count[9][10] , \sa_count[9].f.lower[10] );
tran (\sa_count[9][11] , \sa_count[9].r.part0[11] );
tran (\sa_count[9][11] , \sa_count[9].f.lower[11] );
tran (\sa_count[9][12] , \sa_count[9].r.part0[12] );
tran (\sa_count[9][12] , \sa_count[9].f.lower[12] );
tran (\sa_count[9][13] , \sa_count[9].r.part0[13] );
tran (\sa_count[9][13] , \sa_count[9].f.lower[13] );
tran (\sa_count[9][14] , \sa_count[9].r.part0[14] );
tran (\sa_count[9][14] , \sa_count[9].f.lower[14] );
tran (\sa_count[9][15] , \sa_count[9].r.part0[15] );
tran (\sa_count[9][15] , \sa_count[9].f.lower[15] );
tran (\sa_count[9][16] , \sa_count[9].r.part0[16] );
tran (\sa_count[9][16] , \sa_count[9].f.lower[16] );
tran (\sa_count[9][17] , \sa_count[9].r.part0[17] );
tran (\sa_count[9][17] , \sa_count[9].f.lower[17] );
tran (\sa_count[9][18] , \sa_count[9].r.part0[18] );
tran (\sa_count[9][18] , \sa_count[9].f.lower[18] );
tran (\sa_count[9][19] , \sa_count[9].r.part0[19] );
tran (\sa_count[9][19] , \sa_count[9].f.lower[19] );
tran (\sa_count[9][20] , \sa_count[9].r.part0[20] );
tran (\sa_count[9][20] , \sa_count[9].f.lower[20] );
tran (\sa_count[9][21] , \sa_count[9].r.part0[21] );
tran (\sa_count[9][21] , \sa_count[9].f.lower[21] );
tran (\sa_count[9][22] , \sa_count[9].r.part0[22] );
tran (\sa_count[9][22] , \sa_count[9].f.lower[22] );
tran (\sa_count[9][23] , \sa_count[9].r.part0[23] );
tran (\sa_count[9][23] , \sa_count[9].f.lower[23] );
tran (\sa_count[9][24] , \sa_count[9].r.part0[24] );
tran (\sa_count[9][24] , \sa_count[9].f.lower[24] );
tran (\sa_count[9][25] , \sa_count[9].r.part0[25] );
tran (\sa_count[9][25] , \sa_count[9].f.lower[25] );
tran (\sa_count[9][26] , \sa_count[9].r.part0[26] );
tran (\sa_count[9][26] , \sa_count[9].f.lower[26] );
tran (\sa_count[9][27] , \sa_count[9].r.part0[27] );
tran (\sa_count[9][27] , \sa_count[9].f.lower[27] );
tran (\sa_count[9][28] , \sa_count[9].r.part0[28] );
tran (\sa_count[9][28] , \sa_count[9].f.lower[28] );
tran (\sa_count[9][29] , \sa_count[9].r.part0[29] );
tran (\sa_count[9][29] , \sa_count[9].f.lower[29] );
tran (\sa_count[9][30] , \sa_count[9].r.part0[30] );
tran (\sa_count[9][30] , \sa_count[9].f.lower[30] );
tran (\sa_count[9][31] , \sa_count[9].r.part0[31] );
tran (\sa_count[9][31] , \sa_count[9].f.lower[31] );
tran (\sa_count[9][32] , \sa_count[9].r.part1[0] );
tran (\sa_count[9][32] , \sa_count[9].f.upper[0] );
tran (\sa_count[9][33] , \sa_count[9].r.part1[1] );
tran (\sa_count[9][33] , \sa_count[9].f.upper[1] );
tran (\sa_count[9][34] , \sa_count[9].r.part1[2] );
tran (\sa_count[9][34] , \sa_count[9].f.upper[2] );
tran (\sa_count[9][35] , \sa_count[9].r.part1[3] );
tran (\sa_count[9][35] , \sa_count[9].f.upper[3] );
tran (\sa_count[9][36] , \sa_count[9].r.part1[4] );
tran (\sa_count[9][36] , \sa_count[9].f.upper[4] );
tran (\sa_count[9][37] , \sa_count[9].r.part1[5] );
tran (\sa_count[9][37] , \sa_count[9].f.upper[5] );
tran (\sa_count[9][38] , \sa_count[9].r.part1[6] );
tran (\sa_count[9][38] , \sa_count[9].f.upper[6] );
tran (\sa_count[9][39] , \sa_count[9].r.part1[7] );
tran (\sa_count[9][39] , \sa_count[9].f.upper[7] );
tran (\sa_count[9][40] , \sa_count[9].r.part1[8] );
tran (\sa_count[9][40] , \sa_count[9].f.upper[8] );
tran (\sa_count[9][41] , \sa_count[9].r.part1[9] );
tran (\sa_count[9][41] , \sa_count[9].f.upper[9] );
tran (\sa_count[9][42] , \sa_count[9].r.part1[10] );
tran (\sa_count[9][42] , \sa_count[9].f.upper[10] );
tran (\sa_count[9][43] , \sa_count[9].r.part1[11] );
tran (\sa_count[9][43] , \sa_count[9].f.upper[11] );
tran (\sa_count[9][44] , \sa_count[9].r.part1[12] );
tran (\sa_count[9][44] , \sa_count[9].f.upper[12] );
tran (\sa_count[9][45] , \sa_count[9].r.part1[13] );
tran (\sa_count[9][45] , \sa_count[9].f.upper[13] );
tran (\sa_count[9][46] , \sa_count[9].r.part1[14] );
tran (\sa_count[9][46] , \sa_count[9].f.upper[14] );
tran (\sa_count[9][47] , \sa_count[9].r.part1[15] );
tran (\sa_count[9][47] , \sa_count[9].f.upper[15] );
tran (\sa_count[9][48] , \sa_count[9].r.part1[16] );
tran (\sa_count[9][48] , \sa_count[9].f.upper[16] );
tran (\sa_count[9][49] , \sa_count[9].r.part1[17] );
tran (\sa_count[9][49] , \sa_count[9].f.upper[17] );
tran (\sa_count[9][50] , \sa_count[9].r.part1[18] );
tran (\sa_count[9][50] , \sa_count[9].f.unused[0] );
tran (\sa_count[9][51] , \sa_count[9].r.part1[19] );
tran (\sa_count[9][51] , \sa_count[9].f.unused[1] );
tran (\sa_count[9][52] , \sa_count[9].r.part1[20] );
tran (\sa_count[9][52] , \sa_count[9].f.unused[2] );
tran (\sa_count[9][53] , \sa_count[9].r.part1[21] );
tran (\sa_count[9][53] , \sa_count[9].f.unused[3] );
tran (\sa_count[9][54] , \sa_count[9].r.part1[22] );
tran (\sa_count[9][54] , \sa_count[9].f.unused[4] );
tran (\sa_count[9][55] , \sa_count[9].r.part1[23] );
tran (\sa_count[9][55] , \sa_count[9].f.unused[5] );
tran (\sa_count[9][56] , \sa_count[9].r.part1[24] );
tran (\sa_count[9][56] , \sa_count[9].f.unused[6] );
tran (\sa_count[9][57] , \sa_count[9].r.part1[25] );
tran (\sa_count[9][57] , \sa_count[9].f.unused[7] );
tran (\sa_count[9][58] , \sa_count[9].r.part1[26] );
tran (\sa_count[9][58] , \sa_count[9].f.unused[8] );
tran (\sa_count[9][59] , \sa_count[9].r.part1[27] );
tran (\sa_count[9][59] , \sa_count[9].f.unused[9] );
tran (\sa_count[9][60] , \sa_count[9].r.part1[28] );
tran (\sa_count[9][60] , \sa_count[9].f.unused[10] );
tran (\sa_count[9][61] , \sa_count[9].r.part1[29] );
tran (\sa_count[9][61] , \sa_count[9].f.unused[11] );
tran (\sa_count[9][62] , \sa_count[9].r.part1[30] );
tran (\sa_count[9][62] , \sa_count[9].f.unused[12] );
tran (\sa_count[9][63] , \sa_count[9].r.part1[31] );
tran (\sa_count[9][63] , \sa_count[9].f.unused[13] );
tran (\sa_count[10][0] , \sa_count[10].r.part0[0] );
tran (\sa_count[10][0] , \sa_count[10].f.lower[0] );
tran (\sa_count[10][1] , \sa_count[10].r.part0[1] );
tran (\sa_count[10][1] , \sa_count[10].f.lower[1] );
tran (\sa_count[10][2] , \sa_count[10].r.part0[2] );
tran (\sa_count[10][2] , \sa_count[10].f.lower[2] );
tran (\sa_count[10][3] , \sa_count[10].r.part0[3] );
tran (\sa_count[10][3] , \sa_count[10].f.lower[3] );
tran (\sa_count[10][4] , \sa_count[10].r.part0[4] );
tran (\sa_count[10][4] , \sa_count[10].f.lower[4] );
tran (\sa_count[10][5] , \sa_count[10].r.part0[5] );
tran (\sa_count[10][5] , \sa_count[10].f.lower[5] );
tran (\sa_count[10][6] , \sa_count[10].r.part0[6] );
tran (\sa_count[10][6] , \sa_count[10].f.lower[6] );
tran (\sa_count[10][7] , \sa_count[10].r.part0[7] );
tran (\sa_count[10][7] , \sa_count[10].f.lower[7] );
tran (\sa_count[10][8] , \sa_count[10].r.part0[8] );
tran (\sa_count[10][8] , \sa_count[10].f.lower[8] );
tran (\sa_count[10][9] , \sa_count[10].r.part0[9] );
tran (\sa_count[10][9] , \sa_count[10].f.lower[9] );
tran (\sa_count[10][10] , \sa_count[10].r.part0[10] );
tran (\sa_count[10][10] , \sa_count[10].f.lower[10] );
tran (\sa_count[10][11] , \sa_count[10].r.part0[11] );
tran (\sa_count[10][11] , \sa_count[10].f.lower[11] );
tran (\sa_count[10][12] , \sa_count[10].r.part0[12] );
tran (\sa_count[10][12] , \sa_count[10].f.lower[12] );
tran (\sa_count[10][13] , \sa_count[10].r.part0[13] );
tran (\sa_count[10][13] , \sa_count[10].f.lower[13] );
tran (\sa_count[10][14] , \sa_count[10].r.part0[14] );
tran (\sa_count[10][14] , \sa_count[10].f.lower[14] );
tran (\sa_count[10][15] , \sa_count[10].r.part0[15] );
tran (\sa_count[10][15] , \sa_count[10].f.lower[15] );
tran (\sa_count[10][16] , \sa_count[10].r.part0[16] );
tran (\sa_count[10][16] , \sa_count[10].f.lower[16] );
tran (\sa_count[10][17] , \sa_count[10].r.part0[17] );
tran (\sa_count[10][17] , \sa_count[10].f.lower[17] );
tran (\sa_count[10][18] , \sa_count[10].r.part0[18] );
tran (\sa_count[10][18] , \sa_count[10].f.lower[18] );
tran (\sa_count[10][19] , \sa_count[10].r.part0[19] );
tran (\sa_count[10][19] , \sa_count[10].f.lower[19] );
tran (\sa_count[10][20] , \sa_count[10].r.part0[20] );
tran (\sa_count[10][20] , \sa_count[10].f.lower[20] );
tran (\sa_count[10][21] , \sa_count[10].r.part0[21] );
tran (\sa_count[10][21] , \sa_count[10].f.lower[21] );
tran (\sa_count[10][22] , \sa_count[10].r.part0[22] );
tran (\sa_count[10][22] , \sa_count[10].f.lower[22] );
tran (\sa_count[10][23] , \sa_count[10].r.part0[23] );
tran (\sa_count[10][23] , \sa_count[10].f.lower[23] );
tran (\sa_count[10][24] , \sa_count[10].r.part0[24] );
tran (\sa_count[10][24] , \sa_count[10].f.lower[24] );
tran (\sa_count[10][25] , \sa_count[10].r.part0[25] );
tran (\sa_count[10][25] , \sa_count[10].f.lower[25] );
tran (\sa_count[10][26] , \sa_count[10].r.part0[26] );
tran (\sa_count[10][26] , \sa_count[10].f.lower[26] );
tran (\sa_count[10][27] , \sa_count[10].r.part0[27] );
tran (\sa_count[10][27] , \sa_count[10].f.lower[27] );
tran (\sa_count[10][28] , \sa_count[10].r.part0[28] );
tran (\sa_count[10][28] , \sa_count[10].f.lower[28] );
tran (\sa_count[10][29] , \sa_count[10].r.part0[29] );
tran (\sa_count[10][29] , \sa_count[10].f.lower[29] );
tran (\sa_count[10][30] , \sa_count[10].r.part0[30] );
tran (\sa_count[10][30] , \sa_count[10].f.lower[30] );
tran (\sa_count[10][31] , \sa_count[10].r.part0[31] );
tran (\sa_count[10][31] , \sa_count[10].f.lower[31] );
tran (\sa_count[10][32] , \sa_count[10].r.part1[0] );
tran (\sa_count[10][32] , \sa_count[10].f.upper[0] );
tran (\sa_count[10][33] , \sa_count[10].r.part1[1] );
tran (\sa_count[10][33] , \sa_count[10].f.upper[1] );
tran (\sa_count[10][34] , \sa_count[10].r.part1[2] );
tran (\sa_count[10][34] , \sa_count[10].f.upper[2] );
tran (\sa_count[10][35] , \sa_count[10].r.part1[3] );
tran (\sa_count[10][35] , \sa_count[10].f.upper[3] );
tran (\sa_count[10][36] , \sa_count[10].r.part1[4] );
tran (\sa_count[10][36] , \sa_count[10].f.upper[4] );
tran (\sa_count[10][37] , \sa_count[10].r.part1[5] );
tran (\sa_count[10][37] , \sa_count[10].f.upper[5] );
tran (\sa_count[10][38] , \sa_count[10].r.part1[6] );
tran (\sa_count[10][38] , \sa_count[10].f.upper[6] );
tran (\sa_count[10][39] , \sa_count[10].r.part1[7] );
tran (\sa_count[10][39] , \sa_count[10].f.upper[7] );
tran (\sa_count[10][40] , \sa_count[10].r.part1[8] );
tran (\sa_count[10][40] , \sa_count[10].f.upper[8] );
tran (\sa_count[10][41] , \sa_count[10].r.part1[9] );
tran (\sa_count[10][41] , \sa_count[10].f.upper[9] );
tran (\sa_count[10][42] , \sa_count[10].r.part1[10] );
tran (\sa_count[10][42] , \sa_count[10].f.upper[10] );
tran (\sa_count[10][43] , \sa_count[10].r.part1[11] );
tran (\sa_count[10][43] , \sa_count[10].f.upper[11] );
tran (\sa_count[10][44] , \sa_count[10].r.part1[12] );
tran (\sa_count[10][44] , \sa_count[10].f.upper[12] );
tran (\sa_count[10][45] , \sa_count[10].r.part1[13] );
tran (\sa_count[10][45] , \sa_count[10].f.upper[13] );
tran (\sa_count[10][46] , \sa_count[10].r.part1[14] );
tran (\sa_count[10][46] , \sa_count[10].f.upper[14] );
tran (\sa_count[10][47] , \sa_count[10].r.part1[15] );
tran (\sa_count[10][47] , \sa_count[10].f.upper[15] );
tran (\sa_count[10][48] , \sa_count[10].r.part1[16] );
tran (\sa_count[10][48] , \sa_count[10].f.upper[16] );
tran (\sa_count[10][49] , \sa_count[10].r.part1[17] );
tran (\sa_count[10][49] , \sa_count[10].f.upper[17] );
tran (\sa_count[10][50] , \sa_count[10].r.part1[18] );
tran (\sa_count[10][50] , \sa_count[10].f.unused[0] );
tran (\sa_count[10][51] , \sa_count[10].r.part1[19] );
tran (\sa_count[10][51] , \sa_count[10].f.unused[1] );
tran (\sa_count[10][52] , \sa_count[10].r.part1[20] );
tran (\sa_count[10][52] , \sa_count[10].f.unused[2] );
tran (\sa_count[10][53] , \sa_count[10].r.part1[21] );
tran (\sa_count[10][53] , \sa_count[10].f.unused[3] );
tran (\sa_count[10][54] , \sa_count[10].r.part1[22] );
tran (\sa_count[10][54] , \sa_count[10].f.unused[4] );
tran (\sa_count[10][55] , \sa_count[10].r.part1[23] );
tran (\sa_count[10][55] , \sa_count[10].f.unused[5] );
tran (\sa_count[10][56] , \sa_count[10].r.part1[24] );
tran (\sa_count[10][56] , \sa_count[10].f.unused[6] );
tran (\sa_count[10][57] , \sa_count[10].r.part1[25] );
tran (\sa_count[10][57] , \sa_count[10].f.unused[7] );
tran (\sa_count[10][58] , \sa_count[10].r.part1[26] );
tran (\sa_count[10][58] , \sa_count[10].f.unused[8] );
tran (\sa_count[10][59] , \sa_count[10].r.part1[27] );
tran (\sa_count[10][59] , \sa_count[10].f.unused[9] );
tran (\sa_count[10][60] , \sa_count[10].r.part1[28] );
tran (\sa_count[10][60] , \sa_count[10].f.unused[10] );
tran (\sa_count[10][61] , \sa_count[10].r.part1[29] );
tran (\sa_count[10][61] , \sa_count[10].f.unused[11] );
tran (\sa_count[10][62] , \sa_count[10].r.part1[30] );
tran (\sa_count[10][62] , \sa_count[10].f.unused[12] );
tran (\sa_count[10][63] , \sa_count[10].r.part1[31] );
tran (\sa_count[10][63] , \sa_count[10].f.unused[13] );
tran (\sa_count[11][0] , \sa_count[11].r.part0[0] );
tran (\sa_count[11][0] , \sa_count[11].f.lower[0] );
tran (\sa_count[11][1] , \sa_count[11].r.part0[1] );
tran (\sa_count[11][1] , \sa_count[11].f.lower[1] );
tran (\sa_count[11][2] , \sa_count[11].r.part0[2] );
tran (\sa_count[11][2] , \sa_count[11].f.lower[2] );
tran (\sa_count[11][3] , \sa_count[11].r.part0[3] );
tran (\sa_count[11][3] , \sa_count[11].f.lower[3] );
tran (\sa_count[11][4] , \sa_count[11].r.part0[4] );
tran (\sa_count[11][4] , \sa_count[11].f.lower[4] );
tran (\sa_count[11][5] , \sa_count[11].r.part0[5] );
tran (\sa_count[11][5] , \sa_count[11].f.lower[5] );
tran (\sa_count[11][6] , \sa_count[11].r.part0[6] );
tran (\sa_count[11][6] , \sa_count[11].f.lower[6] );
tran (\sa_count[11][7] , \sa_count[11].r.part0[7] );
tran (\sa_count[11][7] , \sa_count[11].f.lower[7] );
tran (\sa_count[11][8] , \sa_count[11].r.part0[8] );
tran (\sa_count[11][8] , \sa_count[11].f.lower[8] );
tran (\sa_count[11][9] , \sa_count[11].r.part0[9] );
tran (\sa_count[11][9] , \sa_count[11].f.lower[9] );
tran (\sa_count[11][10] , \sa_count[11].r.part0[10] );
tran (\sa_count[11][10] , \sa_count[11].f.lower[10] );
tran (\sa_count[11][11] , \sa_count[11].r.part0[11] );
tran (\sa_count[11][11] , \sa_count[11].f.lower[11] );
tran (\sa_count[11][12] , \sa_count[11].r.part0[12] );
tran (\sa_count[11][12] , \sa_count[11].f.lower[12] );
tran (\sa_count[11][13] , \sa_count[11].r.part0[13] );
tran (\sa_count[11][13] , \sa_count[11].f.lower[13] );
tran (\sa_count[11][14] , \sa_count[11].r.part0[14] );
tran (\sa_count[11][14] , \sa_count[11].f.lower[14] );
tran (\sa_count[11][15] , \sa_count[11].r.part0[15] );
tran (\sa_count[11][15] , \sa_count[11].f.lower[15] );
tran (\sa_count[11][16] , \sa_count[11].r.part0[16] );
tran (\sa_count[11][16] , \sa_count[11].f.lower[16] );
tran (\sa_count[11][17] , \sa_count[11].r.part0[17] );
tran (\sa_count[11][17] , \sa_count[11].f.lower[17] );
tran (\sa_count[11][18] , \sa_count[11].r.part0[18] );
tran (\sa_count[11][18] , \sa_count[11].f.lower[18] );
tran (\sa_count[11][19] , \sa_count[11].r.part0[19] );
tran (\sa_count[11][19] , \sa_count[11].f.lower[19] );
tran (\sa_count[11][20] , \sa_count[11].r.part0[20] );
tran (\sa_count[11][20] , \sa_count[11].f.lower[20] );
tran (\sa_count[11][21] , \sa_count[11].r.part0[21] );
tran (\sa_count[11][21] , \sa_count[11].f.lower[21] );
tran (\sa_count[11][22] , \sa_count[11].r.part0[22] );
tran (\sa_count[11][22] , \sa_count[11].f.lower[22] );
tran (\sa_count[11][23] , \sa_count[11].r.part0[23] );
tran (\sa_count[11][23] , \sa_count[11].f.lower[23] );
tran (\sa_count[11][24] , \sa_count[11].r.part0[24] );
tran (\sa_count[11][24] , \sa_count[11].f.lower[24] );
tran (\sa_count[11][25] , \sa_count[11].r.part0[25] );
tran (\sa_count[11][25] , \sa_count[11].f.lower[25] );
tran (\sa_count[11][26] , \sa_count[11].r.part0[26] );
tran (\sa_count[11][26] , \sa_count[11].f.lower[26] );
tran (\sa_count[11][27] , \sa_count[11].r.part0[27] );
tran (\sa_count[11][27] , \sa_count[11].f.lower[27] );
tran (\sa_count[11][28] , \sa_count[11].r.part0[28] );
tran (\sa_count[11][28] , \sa_count[11].f.lower[28] );
tran (\sa_count[11][29] , \sa_count[11].r.part0[29] );
tran (\sa_count[11][29] , \sa_count[11].f.lower[29] );
tran (\sa_count[11][30] , \sa_count[11].r.part0[30] );
tran (\sa_count[11][30] , \sa_count[11].f.lower[30] );
tran (\sa_count[11][31] , \sa_count[11].r.part0[31] );
tran (\sa_count[11][31] , \sa_count[11].f.lower[31] );
tran (\sa_count[11][32] , \sa_count[11].r.part1[0] );
tran (\sa_count[11][32] , \sa_count[11].f.upper[0] );
tran (\sa_count[11][33] , \sa_count[11].r.part1[1] );
tran (\sa_count[11][33] , \sa_count[11].f.upper[1] );
tran (\sa_count[11][34] , \sa_count[11].r.part1[2] );
tran (\sa_count[11][34] , \sa_count[11].f.upper[2] );
tran (\sa_count[11][35] , \sa_count[11].r.part1[3] );
tran (\sa_count[11][35] , \sa_count[11].f.upper[3] );
tran (\sa_count[11][36] , \sa_count[11].r.part1[4] );
tran (\sa_count[11][36] , \sa_count[11].f.upper[4] );
tran (\sa_count[11][37] , \sa_count[11].r.part1[5] );
tran (\sa_count[11][37] , \sa_count[11].f.upper[5] );
tran (\sa_count[11][38] , \sa_count[11].r.part1[6] );
tran (\sa_count[11][38] , \sa_count[11].f.upper[6] );
tran (\sa_count[11][39] , \sa_count[11].r.part1[7] );
tran (\sa_count[11][39] , \sa_count[11].f.upper[7] );
tran (\sa_count[11][40] , \sa_count[11].r.part1[8] );
tran (\sa_count[11][40] , \sa_count[11].f.upper[8] );
tran (\sa_count[11][41] , \sa_count[11].r.part1[9] );
tran (\sa_count[11][41] , \sa_count[11].f.upper[9] );
tran (\sa_count[11][42] , \sa_count[11].r.part1[10] );
tran (\sa_count[11][42] , \sa_count[11].f.upper[10] );
tran (\sa_count[11][43] , \sa_count[11].r.part1[11] );
tran (\sa_count[11][43] , \sa_count[11].f.upper[11] );
tran (\sa_count[11][44] , \sa_count[11].r.part1[12] );
tran (\sa_count[11][44] , \sa_count[11].f.upper[12] );
tran (\sa_count[11][45] , \sa_count[11].r.part1[13] );
tran (\sa_count[11][45] , \sa_count[11].f.upper[13] );
tran (\sa_count[11][46] , \sa_count[11].r.part1[14] );
tran (\sa_count[11][46] , \sa_count[11].f.upper[14] );
tran (\sa_count[11][47] , \sa_count[11].r.part1[15] );
tran (\sa_count[11][47] , \sa_count[11].f.upper[15] );
tran (\sa_count[11][48] , \sa_count[11].r.part1[16] );
tran (\sa_count[11][48] , \sa_count[11].f.upper[16] );
tran (\sa_count[11][49] , \sa_count[11].r.part1[17] );
tran (\sa_count[11][49] , \sa_count[11].f.upper[17] );
tran (\sa_count[11][50] , \sa_count[11].r.part1[18] );
tran (\sa_count[11][50] , \sa_count[11].f.unused[0] );
tran (\sa_count[11][51] , \sa_count[11].r.part1[19] );
tran (\sa_count[11][51] , \sa_count[11].f.unused[1] );
tran (\sa_count[11][52] , \sa_count[11].r.part1[20] );
tran (\sa_count[11][52] , \sa_count[11].f.unused[2] );
tran (\sa_count[11][53] , \sa_count[11].r.part1[21] );
tran (\sa_count[11][53] , \sa_count[11].f.unused[3] );
tran (\sa_count[11][54] , \sa_count[11].r.part1[22] );
tran (\sa_count[11][54] , \sa_count[11].f.unused[4] );
tran (\sa_count[11][55] , \sa_count[11].r.part1[23] );
tran (\sa_count[11][55] , \sa_count[11].f.unused[5] );
tran (\sa_count[11][56] , \sa_count[11].r.part1[24] );
tran (\sa_count[11][56] , \sa_count[11].f.unused[6] );
tran (\sa_count[11][57] , \sa_count[11].r.part1[25] );
tran (\sa_count[11][57] , \sa_count[11].f.unused[7] );
tran (\sa_count[11][58] , \sa_count[11].r.part1[26] );
tran (\sa_count[11][58] , \sa_count[11].f.unused[8] );
tran (\sa_count[11][59] , \sa_count[11].r.part1[27] );
tran (\sa_count[11][59] , \sa_count[11].f.unused[9] );
tran (\sa_count[11][60] , \sa_count[11].r.part1[28] );
tran (\sa_count[11][60] , \sa_count[11].f.unused[10] );
tran (\sa_count[11][61] , \sa_count[11].r.part1[29] );
tran (\sa_count[11][61] , \sa_count[11].f.unused[11] );
tran (\sa_count[11][62] , \sa_count[11].r.part1[30] );
tran (\sa_count[11][62] , \sa_count[11].f.unused[12] );
tran (\sa_count[11][63] , \sa_count[11].r.part1[31] );
tran (\sa_count[11][63] , \sa_count[11].f.unused[13] );
tran (\sa_count[12][0] , \sa_count[12].r.part0[0] );
tran (\sa_count[12][0] , \sa_count[12].f.lower[0] );
tran (\sa_count[12][1] , \sa_count[12].r.part0[1] );
tran (\sa_count[12][1] , \sa_count[12].f.lower[1] );
tran (\sa_count[12][2] , \sa_count[12].r.part0[2] );
tran (\sa_count[12][2] , \sa_count[12].f.lower[2] );
tran (\sa_count[12][3] , \sa_count[12].r.part0[3] );
tran (\sa_count[12][3] , \sa_count[12].f.lower[3] );
tran (\sa_count[12][4] , \sa_count[12].r.part0[4] );
tran (\sa_count[12][4] , \sa_count[12].f.lower[4] );
tran (\sa_count[12][5] , \sa_count[12].r.part0[5] );
tran (\sa_count[12][5] , \sa_count[12].f.lower[5] );
tran (\sa_count[12][6] , \sa_count[12].r.part0[6] );
tran (\sa_count[12][6] , \sa_count[12].f.lower[6] );
tran (\sa_count[12][7] , \sa_count[12].r.part0[7] );
tran (\sa_count[12][7] , \sa_count[12].f.lower[7] );
tran (\sa_count[12][8] , \sa_count[12].r.part0[8] );
tran (\sa_count[12][8] , \sa_count[12].f.lower[8] );
tran (\sa_count[12][9] , \sa_count[12].r.part0[9] );
tran (\sa_count[12][9] , \sa_count[12].f.lower[9] );
tran (\sa_count[12][10] , \sa_count[12].r.part0[10] );
tran (\sa_count[12][10] , \sa_count[12].f.lower[10] );
tran (\sa_count[12][11] , \sa_count[12].r.part0[11] );
tran (\sa_count[12][11] , \sa_count[12].f.lower[11] );
tran (\sa_count[12][12] , \sa_count[12].r.part0[12] );
tran (\sa_count[12][12] , \sa_count[12].f.lower[12] );
tran (\sa_count[12][13] , \sa_count[12].r.part0[13] );
tran (\sa_count[12][13] , \sa_count[12].f.lower[13] );
tran (\sa_count[12][14] , \sa_count[12].r.part0[14] );
tran (\sa_count[12][14] , \sa_count[12].f.lower[14] );
tran (\sa_count[12][15] , \sa_count[12].r.part0[15] );
tran (\sa_count[12][15] , \sa_count[12].f.lower[15] );
tran (\sa_count[12][16] , \sa_count[12].r.part0[16] );
tran (\sa_count[12][16] , \sa_count[12].f.lower[16] );
tran (\sa_count[12][17] , \sa_count[12].r.part0[17] );
tran (\sa_count[12][17] , \sa_count[12].f.lower[17] );
tran (\sa_count[12][18] , \sa_count[12].r.part0[18] );
tran (\sa_count[12][18] , \sa_count[12].f.lower[18] );
tran (\sa_count[12][19] , \sa_count[12].r.part0[19] );
tran (\sa_count[12][19] , \sa_count[12].f.lower[19] );
tran (\sa_count[12][20] , \sa_count[12].r.part0[20] );
tran (\sa_count[12][20] , \sa_count[12].f.lower[20] );
tran (\sa_count[12][21] , \sa_count[12].r.part0[21] );
tran (\sa_count[12][21] , \sa_count[12].f.lower[21] );
tran (\sa_count[12][22] , \sa_count[12].r.part0[22] );
tran (\sa_count[12][22] , \sa_count[12].f.lower[22] );
tran (\sa_count[12][23] , \sa_count[12].r.part0[23] );
tran (\sa_count[12][23] , \sa_count[12].f.lower[23] );
tran (\sa_count[12][24] , \sa_count[12].r.part0[24] );
tran (\sa_count[12][24] , \sa_count[12].f.lower[24] );
tran (\sa_count[12][25] , \sa_count[12].r.part0[25] );
tran (\sa_count[12][25] , \sa_count[12].f.lower[25] );
tran (\sa_count[12][26] , \sa_count[12].r.part0[26] );
tran (\sa_count[12][26] , \sa_count[12].f.lower[26] );
tran (\sa_count[12][27] , \sa_count[12].r.part0[27] );
tran (\sa_count[12][27] , \sa_count[12].f.lower[27] );
tran (\sa_count[12][28] , \sa_count[12].r.part0[28] );
tran (\sa_count[12][28] , \sa_count[12].f.lower[28] );
tran (\sa_count[12][29] , \sa_count[12].r.part0[29] );
tran (\sa_count[12][29] , \sa_count[12].f.lower[29] );
tran (\sa_count[12][30] , \sa_count[12].r.part0[30] );
tran (\sa_count[12][30] , \sa_count[12].f.lower[30] );
tran (\sa_count[12][31] , \sa_count[12].r.part0[31] );
tran (\sa_count[12][31] , \sa_count[12].f.lower[31] );
tran (\sa_count[12][32] , \sa_count[12].r.part1[0] );
tran (\sa_count[12][32] , \sa_count[12].f.upper[0] );
tran (\sa_count[12][33] , \sa_count[12].r.part1[1] );
tran (\sa_count[12][33] , \sa_count[12].f.upper[1] );
tran (\sa_count[12][34] , \sa_count[12].r.part1[2] );
tran (\sa_count[12][34] , \sa_count[12].f.upper[2] );
tran (\sa_count[12][35] , \sa_count[12].r.part1[3] );
tran (\sa_count[12][35] , \sa_count[12].f.upper[3] );
tran (\sa_count[12][36] , \sa_count[12].r.part1[4] );
tran (\sa_count[12][36] , \sa_count[12].f.upper[4] );
tran (\sa_count[12][37] , \sa_count[12].r.part1[5] );
tran (\sa_count[12][37] , \sa_count[12].f.upper[5] );
tran (\sa_count[12][38] , \sa_count[12].r.part1[6] );
tran (\sa_count[12][38] , \sa_count[12].f.upper[6] );
tran (\sa_count[12][39] , \sa_count[12].r.part1[7] );
tran (\sa_count[12][39] , \sa_count[12].f.upper[7] );
tran (\sa_count[12][40] , \sa_count[12].r.part1[8] );
tran (\sa_count[12][40] , \sa_count[12].f.upper[8] );
tran (\sa_count[12][41] , \sa_count[12].r.part1[9] );
tran (\sa_count[12][41] , \sa_count[12].f.upper[9] );
tran (\sa_count[12][42] , \sa_count[12].r.part1[10] );
tran (\sa_count[12][42] , \sa_count[12].f.upper[10] );
tran (\sa_count[12][43] , \sa_count[12].r.part1[11] );
tran (\sa_count[12][43] , \sa_count[12].f.upper[11] );
tran (\sa_count[12][44] , \sa_count[12].r.part1[12] );
tran (\sa_count[12][44] , \sa_count[12].f.upper[12] );
tran (\sa_count[12][45] , \sa_count[12].r.part1[13] );
tran (\sa_count[12][45] , \sa_count[12].f.upper[13] );
tran (\sa_count[12][46] , \sa_count[12].r.part1[14] );
tran (\sa_count[12][46] , \sa_count[12].f.upper[14] );
tran (\sa_count[12][47] , \sa_count[12].r.part1[15] );
tran (\sa_count[12][47] , \sa_count[12].f.upper[15] );
tran (\sa_count[12][48] , \sa_count[12].r.part1[16] );
tran (\sa_count[12][48] , \sa_count[12].f.upper[16] );
tran (\sa_count[12][49] , \sa_count[12].r.part1[17] );
tran (\sa_count[12][49] , \sa_count[12].f.upper[17] );
tran (\sa_count[12][50] , \sa_count[12].r.part1[18] );
tran (\sa_count[12][50] , \sa_count[12].f.unused[0] );
tran (\sa_count[12][51] , \sa_count[12].r.part1[19] );
tran (\sa_count[12][51] , \sa_count[12].f.unused[1] );
tran (\sa_count[12][52] , \sa_count[12].r.part1[20] );
tran (\sa_count[12][52] , \sa_count[12].f.unused[2] );
tran (\sa_count[12][53] , \sa_count[12].r.part1[21] );
tran (\sa_count[12][53] , \sa_count[12].f.unused[3] );
tran (\sa_count[12][54] , \sa_count[12].r.part1[22] );
tran (\sa_count[12][54] , \sa_count[12].f.unused[4] );
tran (\sa_count[12][55] , \sa_count[12].r.part1[23] );
tran (\sa_count[12][55] , \sa_count[12].f.unused[5] );
tran (\sa_count[12][56] , \sa_count[12].r.part1[24] );
tran (\sa_count[12][56] , \sa_count[12].f.unused[6] );
tran (\sa_count[12][57] , \sa_count[12].r.part1[25] );
tran (\sa_count[12][57] , \sa_count[12].f.unused[7] );
tran (\sa_count[12][58] , \sa_count[12].r.part1[26] );
tran (\sa_count[12][58] , \sa_count[12].f.unused[8] );
tran (\sa_count[12][59] , \sa_count[12].r.part1[27] );
tran (\sa_count[12][59] , \sa_count[12].f.unused[9] );
tran (\sa_count[12][60] , \sa_count[12].r.part1[28] );
tran (\sa_count[12][60] , \sa_count[12].f.unused[10] );
tran (\sa_count[12][61] , \sa_count[12].r.part1[29] );
tran (\sa_count[12][61] , \sa_count[12].f.unused[11] );
tran (\sa_count[12][62] , \sa_count[12].r.part1[30] );
tran (\sa_count[12][62] , \sa_count[12].f.unused[12] );
tran (\sa_count[12][63] , \sa_count[12].r.part1[31] );
tran (\sa_count[12][63] , \sa_count[12].f.unused[13] );
tran (\sa_count[13][0] , \sa_count[13].r.part0[0] );
tran (\sa_count[13][0] , \sa_count[13].f.lower[0] );
tran (\sa_count[13][1] , \sa_count[13].r.part0[1] );
tran (\sa_count[13][1] , \sa_count[13].f.lower[1] );
tran (\sa_count[13][2] , \sa_count[13].r.part0[2] );
tran (\sa_count[13][2] , \sa_count[13].f.lower[2] );
tran (\sa_count[13][3] , \sa_count[13].r.part0[3] );
tran (\sa_count[13][3] , \sa_count[13].f.lower[3] );
tran (\sa_count[13][4] , \sa_count[13].r.part0[4] );
tran (\sa_count[13][4] , \sa_count[13].f.lower[4] );
tran (\sa_count[13][5] , \sa_count[13].r.part0[5] );
tran (\sa_count[13][5] , \sa_count[13].f.lower[5] );
tran (\sa_count[13][6] , \sa_count[13].r.part0[6] );
tran (\sa_count[13][6] , \sa_count[13].f.lower[6] );
tran (\sa_count[13][7] , \sa_count[13].r.part0[7] );
tran (\sa_count[13][7] , \sa_count[13].f.lower[7] );
tran (\sa_count[13][8] , \sa_count[13].r.part0[8] );
tran (\sa_count[13][8] , \sa_count[13].f.lower[8] );
tran (\sa_count[13][9] , \sa_count[13].r.part0[9] );
tran (\sa_count[13][9] , \sa_count[13].f.lower[9] );
tran (\sa_count[13][10] , \sa_count[13].r.part0[10] );
tran (\sa_count[13][10] , \sa_count[13].f.lower[10] );
tran (\sa_count[13][11] , \sa_count[13].r.part0[11] );
tran (\sa_count[13][11] , \sa_count[13].f.lower[11] );
tran (\sa_count[13][12] , \sa_count[13].r.part0[12] );
tran (\sa_count[13][12] , \sa_count[13].f.lower[12] );
tran (\sa_count[13][13] , \sa_count[13].r.part0[13] );
tran (\sa_count[13][13] , \sa_count[13].f.lower[13] );
tran (\sa_count[13][14] , \sa_count[13].r.part0[14] );
tran (\sa_count[13][14] , \sa_count[13].f.lower[14] );
tran (\sa_count[13][15] , \sa_count[13].r.part0[15] );
tran (\sa_count[13][15] , \sa_count[13].f.lower[15] );
tran (\sa_count[13][16] , \sa_count[13].r.part0[16] );
tran (\sa_count[13][16] , \sa_count[13].f.lower[16] );
tran (\sa_count[13][17] , \sa_count[13].r.part0[17] );
tran (\sa_count[13][17] , \sa_count[13].f.lower[17] );
tran (\sa_count[13][18] , \sa_count[13].r.part0[18] );
tran (\sa_count[13][18] , \sa_count[13].f.lower[18] );
tran (\sa_count[13][19] , \sa_count[13].r.part0[19] );
tran (\sa_count[13][19] , \sa_count[13].f.lower[19] );
tran (\sa_count[13][20] , \sa_count[13].r.part0[20] );
tran (\sa_count[13][20] , \sa_count[13].f.lower[20] );
tran (\sa_count[13][21] , \sa_count[13].r.part0[21] );
tran (\sa_count[13][21] , \sa_count[13].f.lower[21] );
tran (\sa_count[13][22] , \sa_count[13].r.part0[22] );
tran (\sa_count[13][22] , \sa_count[13].f.lower[22] );
tran (\sa_count[13][23] , \sa_count[13].r.part0[23] );
tran (\sa_count[13][23] , \sa_count[13].f.lower[23] );
tran (\sa_count[13][24] , \sa_count[13].r.part0[24] );
tran (\sa_count[13][24] , \sa_count[13].f.lower[24] );
tran (\sa_count[13][25] , \sa_count[13].r.part0[25] );
tran (\sa_count[13][25] , \sa_count[13].f.lower[25] );
tran (\sa_count[13][26] , \sa_count[13].r.part0[26] );
tran (\sa_count[13][26] , \sa_count[13].f.lower[26] );
tran (\sa_count[13][27] , \sa_count[13].r.part0[27] );
tran (\sa_count[13][27] , \sa_count[13].f.lower[27] );
tran (\sa_count[13][28] , \sa_count[13].r.part0[28] );
tran (\sa_count[13][28] , \sa_count[13].f.lower[28] );
tran (\sa_count[13][29] , \sa_count[13].r.part0[29] );
tran (\sa_count[13][29] , \sa_count[13].f.lower[29] );
tran (\sa_count[13][30] , \sa_count[13].r.part0[30] );
tran (\sa_count[13][30] , \sa_count[13].f.lower[30] );
tran (\sa_count[13][31] , \sa_count[13].r.part0[31] );
tran (\sa_count[13][31] , \sa_count[13].f.lower[31] );
tran (\sa_count[13][32] , \sa_count[13].r.part1[0] );
tran (\sa_count[13][32] , \sa_count[13].f.upper[0] );
tran (\sa_count[13][33] , \sa_count[13].r.part1[1] );
tran (\sa_count[13][33] , \sa_count[13].f.upper[1] );
tran (\sa_count[13][34] , \sa_count[13].r.part1[2] );
tran (\sa_count[13][34] , \sa_count[13].f.upper[2] );
tran (\sa_count[13][35] , \sa_count[13].r.part1[3] );
tran (\sa_count[13][35] , \sa_count[13].f.upper[3] );
tran (\sa_count[13][36] , \sa_count[13].r.part1[4] );
tran (\sa_count[13][36] , \sa_count[13].f.upper[4] );
tran (\sa_count[13][37] , \sa_count[13].r.part1[5] );
tran (\sa_count[13][37] , \sa_count[13].f.upper[5] );
tran (\sa_count[13][38] , \sa_count[13].r.part1[6] );
tran (\sa_count[13][38] , \sa_count[13].f.upper[6] );
tran (\sa_count[13][39] , \sa_count[13].r.part1[7] );
tran (\sa_count[13][39] , \sa_count[13].f.upper[7] );
tran (\sa_count[13][40] , \sa_count[13].r.part1[8] );
tran (\sa_count[13][40] , \sa_count[13].f.upper[8] );
tran (\sa_count[13][41] , \sa_count[13].r.part1[9] );
tran (\sa_count[13][41] , \sa_count[13].f.upper[9] );
tran (\sa_count[13][42] , \sa_count[13].r.part1[10] );
tran (\sa_count[13][42] , \sa_count[13].f.upper[10] );
tran (\sa_count[13][43] , \sa_count[13].r.part1[11] );
tran (\sa_count[13][43] , \sa_count[13].f.upper[11] );
tran (\sa_count[13][44] , \sa_count[13].r.part1[12] );
tran (\sa_count[13][44] , \sa_count[13].f.upper[12] );
tran (\sa_count[13][45] , \sa_count[13].r.part1[13] );
tran (\sa_count[13][45] , \sa_count[13].f.upper[13] );
tran (\sa_count[13][46] , \sa_count[13].r.part1[14] );
tran (\sa_count[13][46] , \sa_count[13].f.upper[14] );
tran (\sa_count[13][47] , \sa_count[13].r.part1[15] );
tran (\sa_count[13][47] , \sa_count[13].f.upper[15] );
tran (\sa_count[13][48] , \sa_count[13].r.part1[16] );
tran (\sa_count[13][48] , \sa_count[13].f.upper[16] );
tran (\sa_count[13][49] , \sa_count[13].r.part1[17] );
tran (\sa_count[13][49] , \sa_count[13].f.upper[17] );
tran (\sa_count[13][50] , \sa_count[13].r.part1[18] );
tran (\sa_count[13][50] , \sa_count[13].f.unused[0] );
tran (\sa_count[13][51] , \sa_count[13].r.part1[19] );
tran (\sa_count[13][51] , \sa_count[13].f.unused[1] );
tran (\sa_count[13][52] , \sa_count[13].r.part1[20] );
tran (\sa_count[13][52] , \sa_count[13].f.unused[2] );
tran (\sa_count[13][53] , \sa_count[13].r.part1[21] );
tran (\sa_count[13][53] , \sa_count[13].f.unused[3] );
tran (\sa_count[13][54] , \sa_count[13].r.part1[22] );
tran (\sa_count[13][54] , \sa_count[13].f.unused[4] );
tran (\sa_count[13][55] , \sa_count[13].r.part1[23] );
tran (\sa_count[13][55] , \sa_count[13].f.unused[5] );
tran (\sa_count[13][56] , \sa_count[13].r.part1[24] );
tran (\sa_count[13][56] , \sa_count[13].f.unused[6] );
tran (\sa_count[13][57] , \sa_count[13].r.part1[25] );
tran (\sa_count[13][57] , \sa_count[13].f.unused[7] );
tran (\sa_count[13][58] , \sa_count[13].r.part1[26] );
tran (\sa_count[13][58] , \sa_count[13].f.unused[8] );
tran (\sa_count[13][59] , \sa_count[13].r.part1[27] );
tran (\sa_count[13][59] , \sa_count[13].f.unused[9] );
tran (\sa_count[13][60] , \sa_count[13].r.part1[28] );
tran (\sa_count[13][60] , \sa_count[13].f.unused[10] );
tran (\sa_count[13][61] , \sa_count[13].r.part1[29] );
tran (\sa_count[13][61] , \sa_count[13].f.unused[11] );
tran (\sa_count[13][62] , \sa_count[13].r.part1[30] );
tran (\sa_count[13][62] , \sa_count[13].f.unused[12] );
tran (\sa_count[13][63] , \sa_count[13].r.part1[31] );
tran (\sa_count[13][63] , \sa_count[13].f.unused[13] );
tran (\sa_count[14][0] , \sa_count[14].r.part0[0] );
tran (\sa_count[14][0] , \sa_count[14].f.lower[0] );
tran (\sa_count[14][1] , \sa_count[14].r.part0[1] );
tran (\sa_count[14][1] , \sa_count[14].f.lower[1] );
tran (\sa_count[14][2] , \sa_count[14].r.part0[2] );
tran (\sa_count[14][2] , \sa_count[14].f.lower[2] );
tran (\sa_count[14][3] , \sa_count[14].r.part0[3] );
tran (\sa_count[14][3] , \sa_count[14].f.lower[3] );
tran (\sa_count[14][4] , \sa_count[14].r.part0[4] );
tran (\sa_count[14][4] , \sa_count[14].f.lower[4] );
tran (\sa_count[14][5] , \sa_count[14].r.part0[5] );
tran (\sa_count[14][5] , \sa_count[14].f.lower[5] );
tran (\sa_count[14][6] , \sa_count[14].r.part0[6] );
tran (\sa_count[14][6] , \sa_count[14].f.lower[6] );
tran (\sa_count[14][7] , \sa_count[14].r.part0[7] );
tran (\sa_count[14][7] , \sa_count[14].f.lower[7] );
tran (\sa_count[14][8] , \sa_count[14].r.part0[8] );
tran (\sa_count[14][8] , \sa_count[14].f.lower[8] );
tran (\sa_count[14][9] , \sa_count[14].r.part0[9] );
tran (\sa_count[14][9] , \sa_count[14].f.lower[9] );
tran (\sa_count[14][10] , \sa_count[14].r.part0[10] );
tran (\sa_count[14][10] , \sa_count[14].f.lower[10] );
tran (\sa_count[14][11] , \sa_count[14].r.part0[11] );
tran (\sa_count[14][11] , \sa_count[14].f.lower[11] );
tran (\sa_count[14][12] , \sa_count[14].r.part0[12] );
tran (\sa_count[14][12] , \sa_count[14].f.lower[12] );
tran (\sa_count[14][13] , \sa_count[14].r.part0[13] );
tran (\sa_count[14][13] , \sa_count[14].f.lower[13] );
tran (\sa_count[14][14] , \sa_count[14].r.part0[14] );
tran (\sa_count[14][14] , \sa_count[14].f.lower[14] );
tran (\sa_count[14][15] , \sa_count[14].r.part0[15] );
tran (\sa_count[14][15] , \sa_count[14].f.lower[15] );
tran (\sa_count[14][16] , \sa_count[14].r.part0[16] );
tran (\sa_count[14][16] , \sa_count[14].f.lower[16] );
tran (\sa_count[14][17] , \sa_count[14].r.part0[17] );
tran (\sa_count[14][17] , \sa_count[14].f.lower[17] );
tran (\sa_count[14][18] , \sa_count[14].r.part0[18] );
tran (\sa_count[14][18] , \sa_count[14].f.lower[18] );
tran (\sa_count[14][19] , \sa_count[14].r.part0[19] );
tran (\sa_count[14][19] , \sa_count[14].f.lower[19] );
tran (\sa_count[14][20] , \sa_count[14].r.part0[20] );
tran (\sa_count[14][20] , \sa_count[14].f.lower[20] );
tran (\sa_count[14][21] , \sa_count[14].r.part0[21] );
tran (\sa_count[14][21] , \sa_count[14].f.lower[21] );
tran (\sa_count[14][22] , \sa_count[14].r.part0[22] );
tran (\sa_count[14][22] , \sa_count[14].f.lower[22] );
tran (\sa_count[14][23] , \sa_count[14].r.part0[23] );
tran (\sa_count[14][23] , \sa_count[14].f.lower[23] );
tran (\sa_count[14][24] , \sa_count[14].r.part0[24] );
tran (\sa_count[14][24] , \sa_count[14].f.lower[24] );
tran (\sa_count[14][25] , \sa_count[14].r.part0[25] );
tran (\sa_count[14][25] , \sa_count[14].f.lower[25] );
tran (\sa_count[14][26] , \sa_count[14].r.part0[26] );
tran (\sa_count[14][26] , \sa_count[14].f.lower[26] );
tran (\sa_count[14][27] , \sa_count[14].r.part0[27] );
tran (\sa_count[14][27] , \sa_count[14].f.lower[27] );
tran (\sa_count[14][28] , \sa_count[14].r.part0[28] );
tran (\sa_count[14][28] , \sa_count[14].f.lower[28] );
tran (\sa_count[14][29] , \sa_count[14].r.part0[29] );
tran (\sa_count[14][29] , \sa_count[14].f.lower[29] );
tran (\sa_count[14][30] , \sa_count[14].r.part0[30] );
tran (\sa_count[14][30] , \sa_count[14].f.lower[30] );
tran (\sa_count[14][31] , \sa_count[14].r.part0[31] );
tran (\sa_count[14][31] , \sa_count[14].f.lower[31] );
tran (\sa_count[14][32] , \sa_count[14].r.part1[0] );
tran (\sa_count[14][32] , \sa_count[14].f.upper[0] );
tran (\sa_count[14][33] , \sa_count[14].r.part1[1] );
tran (\sa_count[14][33] , \sa_count[14].f.upper[1] );
tran (\sa_count[14][34] , \sa_count[14].r.part1[2] );
tran (\sa_count[14][34] , \sa_count[14].f.upper[2] );
tran (\sa_count[14][35] , \sa_count[14].r.part1[3] );
tran (\sa_count[14][35] , \sa_count[14].f.upper[3] );
tran (\sa_count[14][36] , \sa_count[14].r.part1[4] );
tran (\sa_count[14][36] , \sa_count[14].f.upper[4] );
tran (\sa_count[14][37] , \sa_count[14].r.part1[5] );
tran (\sa_count[14][37] , \sa_count[14].f.upper[5] );
tran (\sa_count[14][38] , \sa_count[14].r.part1[6] );
tran (\sa_count[14][38] , \sa_count[14].f.upper[6] );
tran (\sa_count[14][39] , \sa_count[14].r.part1[7] );
tran (\sa_count[14][39] , \sa_count[14].f.upper[7] );
tran (\sa_count[14][40] , \sa_count[14].r.part1[8] );
tran (\sa_count[14][40] , \sa_count[14].f.upper[8] );
tran (\sa_count[14][41] , \sa_count[14].r.part1[9] );
tran (\sa_count[14][41] , \sa_count[14].f.upper[9] );
tran (\sa_count[14][42] , \sa_count[14].r.part1[10] );
tran (\sa_count[14][42] , \sa_count[14].f.upper[10] );
tran (\sa_count[14][43] , \sa_count[14].r.part1[11] );
tran (\sa_count[14][43] , \sa_count[14].f.upper[11] );
tran (\sa_count[14][44] , \sa_count[14].r.part1[12] );
tran (\sa_count[14][44] , \sa_count[14].f.upper[12] );
tran (\sa_count[14][45] , \sa_count[14].r.part1[13] );
tran (\sa_count[14][45] , \sa_count[14].f.upper[13] );
tran (\sa_count[14][46] , \sa_count[14].r.part1[14] );
tran (\sa_count[14][46] , \sa_count[14].f.upper[14] );
tran (\sa_count[14][47] , \sa_count[14].r.part1[15] );
tran (\sa_count[14][47] , \sa_count[14].f.upper[15] );
tran (\sa_count[14][48] , \sa_count[14].r.part1[16] );
tran (\sa_count[14][48] , \sa_count[14].f.upper[16] );
tran (\sa_count[14][49] , \sa_count[14].r.part1[17] );
tran (\sa_count[14][49] , \sa_count[14].f.upper[17] );
tran (\sa_count[14][50] , \sa_count[14].r.part1[18] );
tran (\sa_count[14][50] , \sa_count[14].f.unused[0] );
tran (\sa_count[14][51] , \sa_count[14].r.part1[19] );
tran (\sa_count[14][51] , \sa_count[14].f.unused[1] );
tran (\sa_count[14][52] , \sa_count[14].r.part1[20] );
tran (\sa_count[14][52] , \sa_count[14].f.unused[2] );
tran (\sa_count[14][53] , \sa_count[14].r.part1[21] );
tran (\sa_count[14][53] , \sa_count[14].f.unused[3] );
tran (\sa_count[14][54] , \sa_count[14].r.part1[22] );
tran (\sa_count[14][54] , \sa_count[14].f.unused[4] );
tran (\sa_count[14][55] , \sa_count[14].r.part1[23] );
tran (\sa_count[14][55] , \sa_count[14].f.unused[5] );
tran (\sa_count[14][56] , \sa_count[14].r.part1[24] );
tran (\sa_count[14][56] , \sa_count[14].f.unused[6] );
tran (\sa_count[14][57] , \sa_count[14].r.part1[25] );
tran (\sa_count[14][57] , \sa_count[14].f.unused[7] );
tran (\sa_count[14][58] , \sa_count[14].r.part1[26] );
tran (\sa_count[14][58] , \sa_count[14].f.unused[8] );
tran (\sa_count[14][59] , \sa_count[14].r.part1[27] );
tran (\sa_count[14][59] , \sa_count[14].f.unused[9] );
tran (\sa_count[14][60] , \sa_count[14].r.part1[28] );
tran (\sa_count[14][60] , \sa_count[14].f.unused[10] );
tran (\sa_count[14][61] , \sa_count[14].r.part1[29] );
tran (\sa_count[14][61] , \sa_count[14].f.unused[11] );
tran (\sa_count[14][62] , \sa_count[14].r.part1[30] );
tran (\sa_count[14][62] , \sa_count[14].f.unused[12] );
tran (\sa_count[14][63] , \sa_count[14].r.part1[31] );
tran (\sa_count[14][63] , \sa_count[14].f.unused[13] );
tran (\sa_count[15][0] , \sa_count[15].r.part0[0] );
tran (\sa_count[15][0] , \sa_count[15].f.lower[0] );
tran (\sa_count[15][1] , \sa_count[15].r.part0[1] );
tran (\sa_count[15][1] , \sa_count[15].f.lower[1] );
tran (\sa_count[15][2] , \sa_count[15].r.part0[2] );
tran (\sa_count[15][2] , \sa_count[15].f.lower[2] );
tran (\sa_count[15][3] , \sa_count[15].r.part0[3] );
tran (\sa_count[15][3] , \sa_count[15].f.lower[3] );
tran (\sa_count[15][4] , \sa_count[15].r.part0[4] );
tran (\sa_count[15][4] , \sa_count[15].f.lower[4] );
tran (\sa_count[15][5] , \sa_count[15].r.part0[5] );
tran (\sa_count[15][5] , \sa_count[15].f.lower[5] );
tran (\sa_count[15][6] , \sa_count[15].r.part0[6] );
tran (\sa_count[15][6] , \sa_count[15].f.lower[6] );
tran (\sa_count[15][7] , \sa_count[15].r.part0[7] );
tran (\sa_count[15][7] , \sa_count[15].f.lower[7] );
tran (\sa_count[15][8] , \sa_count[15].r.part0[8] );
tran (\sa_count[15][8] , \sa_count[15].f.lower[8] );
tran (\sa_count[15][9] , \sa_count[15].r.part0[9] );
tran (\sa_count[15][9] , \sa_count[15].f.lower[9] );
tran (\sa_count[15][10] , \sa_count[15].r.part0[10] );
tran (\sa_count[15][10] , \sa_count[15].f.lower[10] );
tran (\sa_count[15][11] , \sa_count[15].r.part0[11] );
tran (\sa_count[15][11] , \sa_count[15].f.lower[11] );
tran (\sa_count[15][12] , \sa_count[15].r.part0[12] );
tran (\sa_count[15][12] , \sa_count[15].f.lower[12] );
tran (\sa_count[15][13] , \sa_count[15].r.part0[13] );
tran (\sa_count[15][13] , \sa_count[15].f.lower[13] );
tran (\sa_count[15][14] , \sa_count[15].r.part0[14] );
tran (\sa_count[15][14] , \sa_count[15].f.lower[14] );
tran (\sa_count[15][15] , \sa_count[15].r.part0[15] );
tran (\sa_count[15][15] , \sa_count[15].f.lower[15] );
tran (\sa_count[15][16] , \sa_count[15].r.part0[16] );
tran (\sa_count[15][16] , \sa_count[15].f.lower[16] );
tran (\sa_count[15][17] , \sa_count[15].r.part0[17] );
tran (\sa_count[15][17] , \sa_count[15].f.lower[17] );
tran (\sa_count[15][18] , \sa_count[15].r.part0[18] );
tran (\sa_count[15][18] , \sa_count[15].f.lower[18] );
tran (\sa_count[15][19] , \sa_count[15].r.part0[19] );
tran (\sa_count[15][19] , \sa_count[15].f.lower[19] );
tran (\sa_count[15][20] , \sa_count[15].r.part0[20] );
tran (\sa_count[15][20] , \sa_count[15].f.lower[20] );
tran (\sa_count[15][21] , \sa_count[15].r.part0[21] );
tran (\sa_count[15][21] , \sa_count[15].f.lower[21] );
tran (\sa_count[15][22] , \sa_count[15].r.part0[22] );
tran (\sa_count[15][22] , \sa_count[15].f.lower[22] );
tran (\sa_count[15][23] , \sa_count[15].r.part0[23] );
tran (\sa_count[15][23] , \sa_count[15].f.lower[23] );
tran (\sa_count[15][24] , \sa_count[15].r.part0[24] );
tran (\sa_count[15][24] , \sa_count[15].f.lower[24] );
tran (\sa_count[15][25] , \sa_count[15].r.part0[25] );
tran (\sa_count[15][25] , \sa_count[15].f.lower[25] );
tran (\sa_count[15][26] , \sa_count[15].r.part0[26] );
tran (\sa_count[15][26] , \sa_count[15].f.lower[26] );
tran (\sa_count[15][27] , \sa_count[15].r.part0[27] );
tran (\sa_count[15][27] , \sa_count[15].f.lower[27] );
tran (\sa_count[15][28] , \sa_count[15].r.part0[28] );
tran (\sa_count[15][28] , \sa_count[15].f.lower[28] );
tran (\sa_count[15][29] , \sa_count[15].r.part0[29] );
tran (\sa_count[15][29] , \sa_count[15].f.lower[29] );
tran (\sa_count[15][30] , \sa_count[15].r.part0[30] );
tran (\sa_count[15][30] , \sa_count[15].f.lower[30] );
tran (\sa_count[15][31] , \sa_count[15].r.part0[31] );
tran (\sa_count[15][31] , \sa_count[15].f.lower[31] );
tran (\sa_count[15][32] , \sa_count[15].r.part1[0] );
tran (\sa_count[15][32] , \sa_count[15].f.upper[0] );
tran (\sa_count[15][33] , \sa_count[15].r.part1[1] );
tran (\sa_count[15][33] , \sa_count[15].f.upper[1] );
tran (\sa_count[15][34] , \sa_count[15].r.part1[2] );
tran (\sa_count[15][34] , \sa_count[15].f.upper[2] );
tran (\sa_count[15][35] , \sa_count[15].r.part1[3] );
tran (\sa_count[15][35] , \sa_count[15].f.upper[3] );
tran (\sa_count[15][36] , \sa_count[15].r.part1[4] );
tran (\sa_count[15][36] , \sa_count[15].f.upper[4] );
tran (\sa_count[15][37] , \sa_count[15].r.part1[5] );
tran (\sa_count[15][37] , \sa_count[15].f.upper[5] );
tran (\sa_count[15][38] , \sa_count[15].r.part1[6] );
tran (\sa_count[15][38] , \sa_count[15].f.upper[6] );
tran (\sa_count[15][39] , \sa_count[15].r.part1[7] );
tran (\sa_count[15][39] , \sa_count[15].f.upper[7] );
tran (\sa_count[15][40] , \sa_count[15].r.part1[8] );
tran (\sa_count[15][40] , \sa_count[15].f.upper[8] );
tran (\sa_count[15][41] , \sa_count[15].r.part1[9] );
tran (\sa_count[15][41] , \sa_count[15].f.upper[9] );
tran (\sa_count[15][42] , \sa_count[15].r.part1[10] );
tran (\sa_count[15][42] , \sa_count[15].f.upper[10] );
tran (\sa_count[15][43] , \sa_count[15].r.part1[11] );
tran (\sa_count[15][43] , \sa_count[15].f.upper[11] );
tran (\sa_count[15][44] , \sa_count[15].r.part1[12] );
tran (\sa_count[15][44] , \sa_count[15].f.upper[12] );
tran (\sa_count[15][45] , \sa_count[15].r.part1[13] );
tran (\sa_count[15][45] , \sa_count[15].f.upper[13] );
tran (\sa_count[15][46] , \sa_count[15].r.part1[14] );
tran (\sa_count[15][46] , \sa_count[15].f.upper[14] );
tran (\sa_count[15][47] , \sa_count[15].r.part1[15] );
tran (\sa_count[15][47] , \sa_count[15].f.upper[15] );
tran (\sa_count[15][48] , \sa_count[15].r.part1[16] );
tran (\sa_count[15][48] , \sa_count[15].f.upper[16] );
tran (\sa_count[15][49] , \sa_count[15].r.part1[17] );
tran (\sa_count[15][49] , \sa_count[15].f.upper[17] );
tran (\sa_count[15][50] , \sa_count[15].r.part1[18] );
tran (\sa_count[15][50] , \sa_count[15].f.unused[0] );
tran (\sa_count[15][51] , \sa_count[15].r.part1[19] );
tran (\sa_count[15][51] , \sa_count[15].f.unused[1] );
tran (\sa_count[15][52] , \sa_count[15].r.part1[20] );
tran (\sa_count[15][52] , \sa_count[15].f.unused[2] );
tran (\sa_count[15][53] , \sa_count[15].r.part1[21] );
tran (\sa_count[15][53] , \sa_count[15].f.unused[3] );
tran (\sa_count[15][54] , \sa_count[15].r.part1[22] );
tran (\sa_count[15][54] , \sa_count[15].f.unused[4] );
tran (\sa_count[15][55] , \sa_count[15].r.part1[23] );
tran (\sa_count[15][55] , \sa_count[15].f.unused[5] );
tran (\sa_count[15][56] , \sa_count[15].r.part1[24] );
tran (\sa_count[15][56] , \sa_count[15].f.unused[6] );
tran (\sa_count[15][57] , \sa_count[15].r.part1[25] );
tran (\sa_count[15][57] , \sa_count[15].f.unused[7] );
tran (\sa_count[15][58] , \sa_count[15].r.part1[26] );
tran (\sa_count[15][58] , \sa_count[15].f.unused[8] );
tran (\sa_count[15][59] , \sa_count[15].r.part1[27] );
tran (\sa_count[15][59] , \sa_count[15].f.unused[9] );
tran (\sa_count[15][60] , \sa_count[15].r.part1[28] );
tran (\sa_count[15][60] , \sa_count[15].f.unused[10] );
tran (\sa_count[15][61] , \sa_count[15].r.part1[29] );
tran (\sa_count[15][61] , \sa_count[15].f.unused[11] );
tran (\sa_count[15][62] , \sa_count[15].r.part1[30] );
tran (\sa_count[15][62] , \sa_count[15].f.unused[12] );
tran (\sa_count[15][63] , \sa_count[15].r.part1[31] );
tran (\sa_count[15][63] , \sa_count[15].f.unused[13] );
tran (\sa_count[16][0] , \sa_count[16].r.part0[0] );
tran (\sa_count[16][0] , \sa_count[16].f.lower[0] );
tran (\sa_count[16][1] , \sa_count[16].r.part0[1] );
tran (\sa_count[16][1] , \sa_count[16].f.lower[1] );
tran (\sa_count[16][2] , \sa_count[16].r.part0[2] );
tran (\sa_count[16][2] , \sa_count[16].f.lower[2] );
tran (\sa_count[16][3] , \sa_count[16].r.part0[3] );
tran (\sa_count[16][3] , \sa_count[16].f.lower[3] );
tran (\sa_count[16][4] , \sa_count[16].r.part0[4] );
tran (\sa_count[16][4] , \sa_count[16].f.lower[4] );
tran (\sa_count[16][5] , \sa_count[16].r.part0[5] );
tran (\sa_count[16][5] , \sa_count[16].f.lower[5] );
tran (\sa_count[16][6] , \sa_count[16].r.part0[6] );
tran (\sa_count[16][6] , \sa_count[16].f.lower[6] );
tran (\sa_count[16][7] , \sa_count[16].r.part0[7] );
tran (\sa_count[16][7] , \sa_count[16].f.lower[7] );
tran (\sa_count[16][8] , \sa_count[16].r.part0[8] );
tran (\sa_count[16][8] , \sa_count[16].f.lower[8] );
tran (\sa_count[16][9] , \sa_count[16].r.part0[9] );
tran (\sa_count[16][9] , \sa_count[16].f.lower[9] );
tran (\sa_count[16][10] , \sa_count[16].r.part0[10] );
tran (\sa_count[16][10] , \sa_count[16].f.lower[10] );
tran (\sa_count[16][11] , \sa_count[16].r.part0[11] );
tran (\sa_count[16][11] , \sa_count[16].f.lower[11] );
tran (\sa_count[16][12] , \sa_count[16].r.part0[12] );
tran (\sa_count[16][12] , \sa_count[16].f.lower[12] );
tran (\sa_count[16][13] , \sa_count[16].r.part0[13] );
tran (\sa_count[16][13] , \sa_count[16].f.lower[13] );
tran (\sa_count[16][14] , \sa_count[16].r.part0[14] );
tran (\sa_count[16][14] , \sa_count[16].f.lower[14] );
tran (\sa_count[16][15] , \sa_count[16].r.part0[15] );
tran (\sa_count[16][15] , \sa_count[16].f.lower[15] );
tran (\sa_count[16][16] , \sa_count[16].r.part0[16] );
tran (\sa_count[16][16] , \sa_count[16].f.lower[16] );
tran (\sa_count[16][17] , \sa_count[16].r.part0[17] );
tran (\sa_count[16][17] , \sa_count[16].f.lower[17] );
tran (\sa_count[16][18] , \sa_count[16].r.part0[18] );
tran (\sa_count[16][18] , \sa_count[16].f.lower[18] );
tran (\sa_count[16][19] , \sa_count[16].r.part0[19] );
tran (\sa_count[16][19] , \sa_count[16].f.lower[19] );
tran (\sa_count[16][20] , \sa_count[16].r.part0[20] );
tran (\sa_count[16][20] , \sa_count[16].f.lower[20] );
tran (\sa_count[16][21] , \sa_count[16].r.part0[21] );
tran (\sa_count[16][21] , \sa_count[16].f.lower[21] );
tran (\sa_count[16][22] , \sa_count[16].r.part0[22] );
tran (\sa_count[16][22] , \sa_count[16].f.lower[22] );
tran (\sa_count[16][23] , \sa_count[16].r.part0[23] );
tran (\sa_count[16][23] , \sa_count[16].f.lower[23] );
tran (\sa_count[16][24] , \sa_count[16].r.part0[24] );
tran (\sa_count[16][24] , \sa_count[16].f.lower[24] );
tran (\sa_count[16][25] , \sa_count[16].r.part0[25] );
tran (\sa_count[16][25] , \sa_count[16].f.lower[25] );
tran (\sa_count[16][26] , \sa_count[16].r.part0[26] );
tran (\sa_count[16][26] , \sa_count[16].f.lower[26] );
tran (\sa_count[16][27] , \sa_count[16].r.part0[27] );
tran (\sa_count[16][27] , \sa_count[16].f.lower[27] );
tran (\sa_count[16][28] , \sa_count[16].r.part0[28] );
tran (\sa_count[16][28] , \sa_count[16].f.lower[28] );
tran (\sa_count[16][29] , \sa_count[16].r.part0[29] );
tran (\sa_count[16][29] , \sa_count[16].f.lower[29] );
tran (\sa_count[16][30] , \sa_count[16].r.part0[30] );
tran (\sa_count[16][30] , \sa_count[16].f.lower[30] );
tran (\sa_count[16][31] , \sa_count[16].r.part0[31] );
tran (\sa_count[16][31] , \sa_count[16].f.lower[31] );
tran (\sa_count[16][32] , \sa_count[16].r.part1[0] );
tran (\sa_count[16][32] , \sa_count[16].f.upper[0] );
tran (\sa_count[16][33] , \sa_count[16].r.part1[1] );
tran (\sa_count[16][33] , \sa_count[16].f.upper[1] );
tran (\sa_count[16][34] , \sa_count[16].r.part1[2] );
tran (\sa_count[16][34] , \sa_count[16].f.upper[2] );
tran (\sa_count[16][35] , \sa_count[16].r.part1[3] );
tran (\sa_count[16][35] , \sa_count[16].f.upper[3] );
tran (\sa_count[16][36] , \sa_count[16].r.part1[4] );
tran (\sa_count[16][36] , \sa_count[16].f.upper[4] );
tran (\sa_count[16][37] , \sa_count[16].r.part1[5] );
tran (\sa_count[16][37] , \sa_count[16].f.upper[5] );
tran (\sa_count[16][38] , \sa_count[16].r.part1[6] );
tran (\sa_count[16][38] , \sa_count[16].f.upper[6] );
tran (\sa_count[16][39] , \sa_count[16].r.part1[7] );
tran (\sa_count[16][39] , \sa_count[16].f.upper[7] );
tran (\sa_count[16][40] , \sa_count[16].r.part1[8] );
tran (\sa_count[16][40] , \sa_count[16].f.upper[8] );
tran (\sa_count[16][41] , \sa_count[16].r.part1[9] );
tran (\sa_count[16][41] , \sa_count[16].f.upper[9] );
tran (\sa_count[16][42] , \sa_count[16].r.part1[10] );
tran (\sa_count[16][42] , \sa_count[16].f.upper[10] );
tran (\sa_count[16][43] , \sa_count[16].r.part1[11] );
tran (\sa_count[16][43] , \sa_count[16].f.upper[11] );
tran (\sa_count[16][44] , \sa_count[16].r.part1[12] );
tran (\sa_count[16][44] , \sa_count[16].f.upper[12] );
tran (\sa_count[16][45] , \sa_count[16].r.part1[13] );
tran (\sa_count[16][45] , \sa_count[16].f.upper[13] );
tran (\sa_count[16][46] , \sa_count[16].r.part1[14] );
tran (\sa_count[16][46] , \sa_count[16].f.upper[14] );
tran (\sa_count[16][47] , \sa_count[16].r.part1[15] );
tran (\sa_count[16][47] , \sa_count[16].f.upper[15] );
tran (\sa_count[16][48] , \sa_count[16].r.part1[16] );
tran (\sa_count[16][48] , \sa_count[16].f.upper[16] );
tran (\sa_count[16][49] , \sa_count[16].r.part1[17] );
tran (\sa_count[16][49] , \sa_count[16].f.upper[17] );
tran (\sa_count[16][50] , \sa_count[16].r.part1[18] );
tran (\sa_count[16][50] , \sa_count[16].f.unused[0] );
tran (\sa_count[16][51] , \sa_count[16].r.part1[19] );
tran (\sa_count[16][51] , \sa_count[16].f.unused[1] );
tran (\sa_count[16][52] , \sa_count[16].r.part1[20] );
tran (\sa_count[16][52] , \sa_count[16].f.unused[2] );
tran (\sa_count[16][53] , \sa_count[16].r.part1[21] );
tran (\sa_count[16][53] , \sa_count[16].f.unused[3] );
tran (\sa_count[16][54] , \sa_count[16].r.part1[22] );
tran (\sa_count[16][54] , \sa_count[16].f.unused[4] );
tran (\sa_count[16][55] , \sa_count[16].r.part1[23] );
tran (\sa_count[16][55] , \sa_count[16].f.unused[5] );
tran (\sa_count[16][56] , \sa_count[16].r.part1[24] );
tran (\sa_count[16][56] , \sa_count[16].f.unused[6] );
tran (\sa_count[16][57] , \sa_count[16].r.part1[25] );
tran (\sa_count[16][57] , \sa_count[16].f.unused[7] );
tran (\sa_count[16][58] , \sa_count[16].r.part1[26] );
tran (\sa_count[16][58] , \sa_count[16].f.unused[8] );
tran (\sa_count[16][59] , \sa_count[16].r.part1[27] );
tran (\sa_count[16][59] , \sa_count[16].f.unused[9] );
tran (\sa_count[16][60] , \sa_count[16].r.part1[28] );
tran (\sa_count[16][60] , \sa_count[16].f.unused[10] );
tran (\sa_count[16][61] , \sa_count[16].r.part1[29] );
tran (\sa_count[16][61] , \sa_count[16].f.unused[11] );
tran (\sa_count[16][62] , \sa_count[16].r.part1[30] );
tran (\sa_count[16][62] , \sa_count[16].f.unused[12] );
tran (\sa_count[16][63] , \sa_count[16].r.part1[31] );
tran (\sa_count[16][63] , \sa_count[16].f.unused[13] );
tran (\sa_count[17][0] , \sa_count[17].r.part0[0] );
tran (\sa_count[17][0] , \sa_count[17].f.lower[0] );
tran (\sa_count[17][1] , \sa_count[17].r.part0[1] );
tran (\sa_count[17][1] , \sa_count[17].f.lower[1] );
tran (\sa_count[17][2] , \sa_count[17].r.part0[2] );
tran (\sa_count[17][2] , \sa_count[17].f.lower[2] );
tran (\sa_count[17][3] , \sa_count[17].r.part0[3] );
tran (\sa_count[17][3] , \sa_count[17].f.lower[3] );
tran (\sa_count[17][4] , \sa_count[17].r.part0[4] );
tran (\sa_count[17][4] , \sa_count[17].f.lower[4] );
tran (\sa_count[17][5] , \sa_count[17].r.part0[5] );
tran (\sa_count[17][5] , \sa_count[17].f.lower[5] );
tran (\sa_count[17][6] , \sa_count[17].r.part0[6] );
tran (\sa_count[17][6] , \sa_count[17].f.lower[6] );
tran (\sa_count[17][7] , \sa_count[17].r.part0[7] );
tran (\sa_count[17][7] , \sa_count[17].f.lower[7] );
tran (\sa_count[17][8] , \sa_count[17].r.part0[8] );
tran (\sa_count[17][8] , \sa_count[17].f.lower[8] );
tran (\sa_count[17][9] , \sa_count[17].r.part0[9] );
tran (\sa_count[17][9] , \sa_count[17].f.lower[9] );
tran (\sa_count[17][10] , \sa_count[17].r.part0[10] );
tran (\sa_count[17][10] , \sa_count[17].f.lower[10] );
tran (\sa_count[17][11] , \sa_count[17].r.part0[11] );
tran (\sa_count[17][11] , \sa_count[17].f.lower[11] );
tran (\sa_count[17][12] , \sa_count[17].r.part0[12] );
tran (\sa_count[17][12] , \sa_count[17].f.lower[12] );
tran (\sa_count[17][13] , \sa_count[17].r.part0[13] );
tran (\sa_count[17][13] , \sa_count[17].f.lower[13] );
tran (\sa_count[17][14] , \sa_count[17].r.part0[14] );
tran (\sa_count[17][14] , \sa_count[17].f.lower[14] );
tran (\sa_count[17][15] , \sa_count[17].r.part0[15] );
tran (\sa_count[17][15] , \sa_count[17].f.lower[15] );
tran (\sa_count[17][16] , \sa_count[17].r.part0[16] );
tran (\sa_count[17][16] , \sa_count[17].f.lower[16] );
tran (\sa_count[17][17] , \sa_count[17].r.part0[17] );
tran (\sa_count[17][17] , \sa_count[17].f.lower[17] );
tran (\sa_count[17][18] , \sa_count[17].r.part0[18] );
tran (\sa_count[17][18] , \sa_count[17].f.lower[18] );
tran (\sa_count[17][19] , \sa_count[17].r.part0[19] );
tran (\sa_count[17][19] , \sa_count[17].f.lower[19] );
tran (\sa_count[17][20] , \sa_count[17].r.part0[20] );
tran (\sa_count[17][20] , \sa_count[17].f.lower[20] );
tran (\sa_count[17][21] , \sa_count[17].r.part0[21] );
tran (\sa_count[17][21] , \sa_count[17].f.lower[21] );
tran (\sa_count[17][22] , \sa_count[17].r.part0[22] );
tran (\sa_count[17][22] , \sa_count[17].f.lower[22] );
tran (\sa_count[17][23] , \sa_count[17].r.part0[23] );
tran (\sa_count[17][23] , \sa_count[17].f.lower[23] );
tran (\sa_count[17][24] , \sa_count[17].r.part0[24] );
tran (\sa_count[17][24] , \sa_count[17].f.lower[24] );
tran (\sa_count[17][25] , \sa_count[17].r.part0[25] );
tran (\sa_count[17][25] , \sa_count[17].f.lower[25] );
tran (\sa_count[17][26] , \sa_count[17].r.part0[26] );
tran (\sa_count[17][26] , \sa_count[17].f.lower[26] );
tran (\sa_count[17][27] , \sa_count[17].r.part0[27] );
tran (\sa_count[17][27] , \sa_count[17].f.lower[27] );
tran (\sa_count[17][28] , \sa_count[17].r.part0[28] );
tran (\sa_count[17][28] , \sa_count[17].f.lower[28] );
tran (\sa_count[17][29] , \sa_count[17].r.part0[29] );
tran (\sa_count[17][29] , \sa_count[17].f.lower[29] );
tran (\sa_count[17][30] , \sa_count[17].r.part0[30] );
tran (\sa_count[17][30] , \sa_count[17].f.lower[30] );
tran (\sa_count[17][31] , \sa_count[17].r.part0[31] );
tran (\sa_count[17][31] , \sa_count[17].f.lower[31] );
tran (\sa_count[17][32] , \sa_count[17].r.part1[0] );
tran (\sa_count[17][32] , \sa_count[17].f.upper[0] );
tran (\sa_count[17][33] , \sa_count[17].r.part1[1] );
tran (\sa_count[17][33] , \sa_count[17].f.upper[1] );
tran (\sa_count[17][34] , \sa_count[17].r.part1[2] );
tran (\sa_count[17][34] , \sa_count[17].f.upper[2] );
tran (\sa_count[17][35] , \sa_count[17].r.part1[3] );
tran (\sa_count[17][35] , \sa_count[17].f.upper[3] );
tran (\sa_count[17][36] , \sa_count[17].r.part1[4] );
tran (\sa_count[17][36] , \sa_count[17].f.upper[4] );
tran (\sa_count[17][37] , \sa_count[17].r.part1[5] );
tran (\sa_count[17][37] , \sa_count[17].f.upper[5] );
tran (\sa_count[17][38] , \sa_count[17].r.part1[6] );
tran (\sa_count[17][38] , \sa_count[17].f.upper[6] );
tran (\sa_count[17][39] , \sa_count[17].r.part1[7] );
tran (\sa_count[17][39] , \sa_count[17].f.upper[7] );
tran (\sa_count[17][40] , \sa_count[17].r.part1[8] );
tran (\sa_count[17][40] , \sa_count[17].f.upper[8] );
tran (\sa_count[17][41] , \sa_count[17].r.part1[9] );
tran (\sa_count[17][41] , \sa_count[17].f.upper[9] );
tran (\sa_count[17][42] , \sa_count[17].r.part1[10] );
tran (\sa_count[17][42] , \sa_count[17].f.upper[10] );
tran (\sa_count[17][43] , \sa_count[17].r.part1[11] );
tran (\sa_count[17][43] , \sa_count[17].f.upper[11] );
tran (\sa_count[17][44] , \sa_count[17].r.part1[12] );
tran (\sa_count[17][44] , \sa_count[17].f.upper[12] );
tran (\sa_count[17][45] , \sa_count[17].r.part1[13] );
tran (\sa_count[17][45] , \sa_count[17].f.upper[13] );
tran (\sa_count[17][46] , \sa_count[17].r.part1[14] );
tran (\sa_count[17][46] , \sa_count[17].f.upper[14] );
tran (\sa_count[17][47] , \sa_count[17].r.part1[15] );
tran (\sa_count[17][47] , \sa_count[17].f.upper[15] );
tran (\sa_count[17][48] , \sa_count[17].r.part1[16] );
tran (\sa_count[17][48] , \sa_count[17].f.upper[16] );
tran (\sa_count[17][49] , \sa_count[17].r.part1[17] );
tran (\sa_count[17][49] , \sa_count[17].f.upper[17] );
tran (\sa_count[17][50] , \sa_count[17].r.part1[18] );
tran (\sa_count[17][50] , \sa_count[17].f.unused[0] );
tran (\sa_count[17][51] , \sa_count[17].r.part1[19] );
tran (\sa_count[17][51] , \sa_count[17].f.unused[1] );
tran (\sa_count[17][52] , \sa_count[17].r.part1[20] );
tran (\sa_count[17][52] , \sa_count[17].f.unused[2] );
tran (\sa_count[17][53] , \sa_count[17].r.part1[21] );
tran (\sa_count[17][53] , \sa_count[17].f.unused[3] );
tran (\sa_count[17][54] , \sa_count[17].r.part1[22] );
tran (\sa_count[17][54] , \sa_count[17].f.unused[4] );
tran (\sa_count[17][55] , \sa_count[17].r.part1[23] );
tran (\sa_count[17][55] , \sa_count[17].f.unused[5] );
tran (\sa_count[17][56] , \sa_count[17].r.part1[24] );
tran (\sa_count[17][56] , \sa_count[17].f.unused[6] );
tran (\sa_count[17][57] , \sa_count[17].r.part1[25] );
tran (\sa_count[17][57] , \sa_count[17].f.unused[7] );
tran (\sa_count[17][58] , \sa_count[17].r.part1[26] );
tran (\sa_count[17][58] , \sa_count[17].f.unused[8] );
tran (\sa_count[17][59] , \sa_count[17].r.part1[27] );
tran (\sa_count[17][59] , \sa_count[17].f.unused[9] );
tran (\sa_count[17][60] , \sa_count[17].r.part1[28] );
tran (\sa_count[17][60] , \sa_count[17].f.unused[10] );
tran (\sa_count[17][61] , \sa_count[17].r.part1[29] );
tran (\sa_count[17][61] , \sa_count[17].f.unused[11] );
tran (\sa_count[17][62] , \sa_count[17].r.part1[30] );
tran (\sa_count[17][62] , \sa_count[17].f.unused[12] );
tran (\sa_count[17][63] , \sa_count[17].r.part1[31] );
tran (\sa_count[17][63] , \sa_count[17].f.unused[13] );
tran (\sa_count[18][0] , \sa_count[18].r.part0[0] );
tran (\sa_count[18][0] , \sa_count[18].f.lower[0] );
tran (\sa_count[18][1] , \sa_count[18].r.part0[1] );
tran (\sa_count[18][1] , \sa_count[18].f.lower[1] );
tran (\sa_count[18][2] , \sa_count[18].r.part0[2] );
tran (\sa_count[18][2] , \sa_count[18].f.lower[2] );
tran (\sa_count[18][3] , \sa_count[18].r.part0[3] );
tran (\sa_count[18][3] , \sa_count[18].f.lower[3] );
tran (\sa_count[18][4] , \sa_count[18].r.part0[4] );
tran (\sa_count[18][4] , \sa_count[18].f.lower[4] );
tran (\sa_count[18][5] , \sa_count[18].r.part0[5] );
tran (\sa_count[18][5] , \sa_count[18].f.lower[5] );
tran (\sa_count[18][6] , \sa_count[18].r.part0[6] );
tran (\sa_count[18][6] , \sa_count[18].f.lower[6] );
tran (\sa_count[18][7] , \sa_count[18].r.part0[7] );
tran (\sa_count[18][7] , \sa_count[18].f.lower[7] );
tran (\sa_count[18][8] , \sa_count[18].r.part0[8] );
tran (\sa_count[18][8] , \sa_count[18].f.lower[8] );
tran (\sa_count[18][9] , \sa_count[18].r.part0[9] );
tran (\sa_count[18][9] , \sa_count[18].f.lower[9] );
tran (\sa_count[18][10] , \sa_count[18].r.part0[10] );
tran (\sa_count[18][10] , \sa_count[18].f.lower[10] );
tran (\sa_count[18][11] , \sa_count[18].r.part0[11] );
tran (\sa_count[18][11] , \sa_count[18].f.lower[11] );
tran (\sa_count[18][12] , \sa_count[18].r.part0[12] );
tran (\sa_count[18][12] , \sa_count[18].f.lower[12] );
tran (\sa_count[18][13] , \sa_count[18].r.part0[13] );
tran (\sa_count[18][13] , \sa_count[18].f.lower[13] );
tran (\sa_count[18][14] , \sa_count[18].r.part0[14] );
tran (\sa_count[18][14] , \sa_count[18].f.lower[14] );
tran (\sa_count[18][15] , \sa_count[18].r.part0[15] );
tran (\sa_count[18][15] , \sa_count[18].f.lower[15] );
tran (\sa_count[18][16] , \sa_count[18].r.part0[16] );
tran (\sa_count[18][16] , \sa_count[18].f.lower[16] );
tran (\sa_count[18][17] , \sa_count[18].r.part0[17] );
tran (\sa_count[18][17] , \sa_count[18].f.lower[17] );
tran (\sa_count[18][18] , \sa_count[18].r.part0[18] );
tran (\sa_count[18][18] , \sa_count[18].f.lower[18] );
tran (\sa_count[18][19] , \sa_count[18].r.part0[19] );
tran (\sa_count[18][19] , \sa_count[18].f.lower[19] );
tran (\sa_count[18][20] , \sa_count[18].r.part0[20] );
tran (\sa_count[18][20] , \sa_count[18].f.lower[20] );
tran (\sa_count[18][21] , \sa_count[18].r.part0[21] );
tran (\sa_count[18][21] , \sa_count[18].f.lower[21] );
tran (\sa_count[18][22] , \sa_count[18].r.part0[22] );
tran (\sa_count[18][22] , \sa_count[18].f.lower[22] );
tran (\sa_count[18][23] , \sa_count[18].r.part0[23] );
tran (\sa_count[18][23] , \sa_count[18].f.lower[23] );
tran (\sa_count[18][24] , \sa_count[18].r.part0[24] );
tran (\sa_count[18][24] , \sa_count[18].f.lower[24] );
tran (\sa_count[18][25] , \sa_count[18].r.part0[25] );
tran (\sa_count[18][25] , \sa_count[18].f.lower[25] );
tran (\sa_count[18][26] , \sa_count[18].r.part0[26] );
tran (\sa_count[18][26] , \sa_count[18].f.lower[26] );
tran (\sa_count[18][27] , \sa_count[18].r.part0[27] );
tran (\sa_count[18][27] , \sa_count[18].f.lower[27] );
tran (\sa_count[18][28] , \sa_count[18].r.part0[28] );
tran (\sa_count[18][28] , \sa_count[18].f.lower[28] );
tran (\sa_count[18][29] , \sa_count[18].r.part0[29] );
tran (\sa_count[18][29] , \sa_count[18].f.lower[29] );
tran (\sa_count[18][30] , \sa_count[18].r.part0[30] );
tran (\sa_count[18][30] , \sa_count[18].f.lower[30] );
tran (\sa_count[18][31] , \sa_count[18].r.part0[31] );
tran (\sa_count[18][31] , \sa_count[18].f.lower[31] );
tran (\sa_count[18][32] , \sa_count[18].r.part1[0] );
tran (\sa_count[18][32] , \sa_count[18].f.upper[0] );
tran (\sa_count[18][33] , \sa_count[18].r.part1[1] );
tran (\sa_count[18][33] , \sa_count[18].f.upper[1] );
tran (\sa_count[18][34] , \sa_count[18].r.part1[2] );
tran (\sa_count[18][34] , \sa_count[18].f.upper[2] );
tran (\sa_count[18][35] , \sa_count[18].r.part1[3] );
tran (\sa_count[18][35] , \sa_count[18].f.upper[3] );
tran (\sa_count[18][36] , \sa_count[18].r.part1[4] );
tran (\sa_count[18][36] , \sa_count[18].f.upper[4] );
tran (\sa_count[18][37] , \sa_count[18].r.part1[5] );
tran (\sa_count[18][37] , \sa_count[18].f.upper[5] );
tran (\sa_count[18][38] , \sa_count[18].r.part1[6] );
tran (\sa_count[18][38] , \sa_count[18].f.upper[6] );
tran (\sa_count[18][39] , \sa_count[18].r.part1[7] );
tran (\sa_count[18][39] , \sa_count[18].f.upper[7] );
tran (\sa_count[18][40] , \sa_count[18].r.part1[8] );
tran (\sa_count[18][40] , \sa_count[18].f.upper[8] );
tran (\sa_count[18][41] , \sa_count[18].r.part1[9] );
tran (\sa_count[18][41] , \sa_count[18].f.upper[9] );
tran (\sa_count[18][42] , \sa_count[18].r.part1[10] );
tran (\sa_count[18][42] , \sa_count[18].f.upper[10] );
tran (\sa_count[18][43] , \sa_count[18].r.part1[11] );
tran (\sa_count[18][43] , \sa_count[18].f.upper[11] );
tran (\sa_count[18][44] , \sa_count[18].r.part1[12] );
tran (\sa_count[18][44] , \sa_count[18].f.upper[12] );
tran (\sa_count[18][45] , \sa_count[18].r.part1[13] );
tran (\sa_count[18][45] , \sa_count[18].f.upper[13] );
tran (\sa_count[18][46] , \sa_count[18].r.part1[14] );
tran (\sa_count[18][46] , \sa_count[18].f.upper[14] );
tran (\sa_count[18][47] , \sa_count[18].r.part1[15] );
tran (\sa_count[18][47] , \sa_count[18].f.upper[15] );
tran (\sa_count[18][48] , \sa_count[18].r.part1[16] );
tran (\sa_count[18][48] , \sa_count[18].f.upper[16] );
tran (\sa_count[18][49] , \sa_count[18].r.part1[17] );
tran (\sa_count[18][49] , \sa_count[18].f.upper[17] );
tran (\sa_count[18][50] , \sa_count[18].r.part1[18] );
tran (\sa_count[18][50] , \sa_count[18].f.unused[0] );
tran (\sa_count[18][51] , \sa_count[18].r.part1[19] );
tran (\sa_count[18][51] , \sa_count[18].f.unused[1] );
tran (\sa_count[18][52] , \sa_count[18].r.part1[20] );
tran (\sa_count[18][52] , \sa_count[18].f.unused[2] );
tran (\sa_count[18][53] , \sa_count[18].r.part1[21] );
tran (\sa_count[18][53] , \sa_count[18].f.unused[3] );
tran (\sa_count[18][54] , \sa_count[18].r.part1[22] );
tran (\sa_count[18][54] , \sa_count[18].f.unused[4] );
tran (\sa_count[18][55] , \sa_count[18].r.part1[23] );
tran (\sa_count[18][55] , \sa_count[18].f.unused[5] );
tran (\sa_count[18][56] , \sa_count[18].r.part1[24] );
tran (\sa_count[18][56] , \sa_count[18].f.unused[6] );
tran (\sa_count[18][57] , \sa_count[18].r.part1[25] );
tran (\sa_count[18][57] , \sa_count[18].f.unused[7] );
tran (\sa_count[18][58] , \sa_count[18].r.part1[26] );
tran (\sa_count[18][58] , \sa_count[18].f.unused[8] );
tran (\sa_count[18][59] , \sa_count[18].r.part1[27] );
tran (\sa_count[18][59] , \sa_count[18].f.unused[9] );
tran (\sa_count[18][60] , \sa_count[18].r.part1[28] );
tran (\sa_count[18][60] , \sa_count[18].f.unused[10] );
tran (\sa_count[18][61] , \sa_count[18].r.part1[29] );
tran (\sa_count[18][61] , \sa_count[18].f.unused[11] );
tran (\sa_count[18][62] , \sa_count[18].r.part1[30] );
tran (\sa_count[18][62] , \sa_count[18].f.unused[12] );
tran (\sa_count[18][63] , \sa_count[18].r.part1[31] );
tran (\sa_count[18][63] , \sa_count[18].f.unused[13] );
tran (\sa_count[19][0] , \sa_count[19].r.part0[0] );
tran (\sa_count[19][0] , \sa_count[19].f.lower[0] );
tran (\sa_count[19][1] , \sa_count[19].r.part0[1] );
tran (\sa_count[19][1] , \sa_count[19].f.lower[1] );
tran (\sa_count[19][2] , \sa_count[19].r.part0[2] );
tran (\sa_count[19][2] , \sa_count[19].f.lower[2] );
tran (\sa_count[19][3] , \sa_count[19].r.part0[3] );
tran (\sa_count[19][3] , \sa_count[19].f.lower[3] );
tran (\sa_count[19][4] , \sa_count[19].r.part0[4] );
tran (\sa_count[19][4] , \sa_count[19].f.lower[4] );
tran (\sa_count[19][5] , \sa_count[19].r.part0[5] );
tran (\sa_count[19][5] , \sa_count[19].f.lower[5] );
tran (\sa_count[19][6] , \sa_count[19].r.part0[6] );
tran (\sa_count[19][6] , \sa_count[19].f.lower[6] );
tran (\sa_count[19][7] , \sa_count[19].r.part0[7] );
tran (\sa_count[19][7] , \sa_count[19].f.lower[7] );
tran (\sa_count[19][8] , \sa_count[19].r.part0[8] );
tran (\sa_count[19][8] , \sa_count[19].f.lower[8] );
tran (\sa_count[19][9] , \sa_count[19].r.part0[9] );
tran (\sa_count[19][9] , \sa_count[19].f.lower[9] );
tran (\sa_count[19][10] , \sa_count[19].r.part0[10] );
tran (\sa_count[19][10] , \sa_count[19].f.lower[10] );
tran (\sa_count[19][11] , \sa_count[19].r.part0[11] );
tran (\sa_count[19][11] , \sa_count[19].f.lower[11] );
tran (\sa_count[19][12] , \sa_count[19].r.part0[12] );
tran (\sa_count[19][12] , \sa_count[19].f.lower[12] );
tran (\sa_count[19][13] , \sa_count[19].r.part0[13] );
tran (\sa_count[19][13] , \sa_count[19].f.lower[13] );
tran (\sa_count[19][14] , \sa_count[19].r.part0[14] );
tran (\sa_count[19][14] , \sa_count[19].f.lower[14] );
tran (\sa_count[19][15] , \sa_count[19].r.part0[15] );
tran (\sa_count[19][15] , \sa_count[19].f.lower[15] );
tran (\sa_count[19][16] , \sa_count[19].r.part0[16] );
tran (\sa_count[19][16] , \sa_count[19].f.lower[16] );
tran (\sa_count[19][17] , \sa_count[19].r.part0[17] );
tran (\sa_count[19][17] , \sa_count[19].f.lower[17] );
tran (\sa_count[19][18] , \sa_count[19].r.part0[18] );
tran (\sa_count[19][18] , \sa_count[19].f.lower[18] );
tran (\sa_count[19][19] , \sa_count[19].r.part0[19] );
tran (\sa_count[19][19] , \sa_count[19].f.lower[19] );
tran (\sa_count[19][20] , \sa_count[19].r.part0[20] );
tran (\sa_count[19][20] , \sa_count[19].f.lower[20] );
tran (\sa_count[19][21] , \sa_count[19].r.part0[21] );
tran (\sa_count[19][21] , \sa_count[19].f.lower[21] );
tran (\sa_count[19][22] , \sa_count[19].r.part0[22] );
tran (\sa_count[19][22] , \sa_count[19].f.lower[22] );
tran (\sa_count[19][23] , \sa_count[19].r.part0[23] );
tran (\sa_count[19][23] , \sa_count[19].f.lower[23] );
tran (\sa_count[19][24] , \sa_count[19].r.part0[24] );
tran (\sa_count[19][24] , \sa_count[19].f.lower[24] );
tran (\sa_count[19][25] , \sa_count[19].r.part0[25] );
tran (\sa_count[19][25] , \sa_count[19].f.lower[25] );
tran (\sa_count[19][26] , \sa_count[19].r.part0[26] );
tran (\sa_count[19][26] , \sa_count[19].f.lower[26] );
tran (\sa_count[19][27] , \sa_count[19].r.part0[27] );
tran (\sa_count[19][27] , \sa_count[19].f.lower[27] );
tran (\sa_count[19][28] , \sa_count[19].r.part0[28] );
tran (\sa_count[19][28] , \sa_count[19].f.lower[28] );
tran (\sa_count[19][29] , \sa_count[19].r.part0[29] );
tran (\sa_count[19][29] , \sa_count[19].f.lower[29] );
tran (\sa_count[19][30] , \sa_count[19].r.part0[30] );
tran (\sa_count[19][30] , \sa_count[19].f.lower[30] );
tran (\sa_count[19][31] , \sa_count[19].r.part0[31] );
tran (\sa_count[19][31] , \sa_count[19].f.lower[31] );
tran (\sa_count[19][32] , \sa_count[19].r.part1[0] );
tran (\sa_count[19][32] , \sa_count[19].f.upper[0] );
tran (\sa_count[19][33] , \sa_count[19].r.part1[1] );
tran (\sa_count[19][33] , \sa_count[19].f.upper[1] );
tran (\sa_count[19][34] , \sa_count[19].r.part1[2] );
tran (\sa_count[19][34] , \sa_count[19].f.upper[2] );
tran (\sa_count[19][35] , \sa_count[19].r.part1[3] );
tran (\sa_count[19][35] , \sa_count[19].f.upper[3] );
tran (\sa_count[19][36] , \sa_count[19].r.part1[4] );
tran (\sa_count[19][36] , \sa_count[19].f.upper[4] );
tran (\sa_count[19][37] , \sa_count[19].r.part1[5] );
tran (\sa_count[19][37] , \sa_count[19].f.upper[5] );
tran (\sa_count[19][38] , \sa_count[19].r.part1[6] );
tran (\sa_count[19][38] , \sa_count[19].f.upper[6] );
tran (\sa_count[19][39] , \sa_count[19].r.part1[7] );
tran (\sa_count[19][39] , \sa_count[19].f.upper[7] );
tran (\sa_count[19][40] , \sa_count[19].r.part1[8] );
tran (\sa_count[19][40] , \sa_count[19].f.upper[8] );
tran (\sa_count[19][41] , \sa_count[19].r.part1[9] );
tran (\sa_count[19][41] , \sa_count[19].f.upper[9] );
tran (\sa_count[19][42] , \sa_count[19].r.part1[10] );
tran (\sa_count[19][42] , \sa_count[19].f.upper[10] );
tran (\sa_count[19][43] , \sa_count[19].r.part1[11] );
tran (\sa_count[19][43] , \sa_count[19].f.upper[11] );
tran (\sa_count[19][44] , \sa_count[19].r.part1[12] );
tran (\sa_count[19][44] , \sa_count[19].f.upper[12] );
tran (\sa_count[19][45] , \sa_count[19].r.part1[13] );
tran (\sa_count[19][45] , \sa_count[19].f.upper[13] );
tran (\sa_count[19][46] , \sa_count[19].r.part1[14] );
tran (\sa_count[19][46] , \sa_count[19].f.upper[14] );
tran (\sa_count[19][47] , \sa_count[19].r.part1[15] );
tran (\sa_count[19][47] , \sa_count[19].f.upper[15] );
tran (\sa_count[19][48] , \sa_count[19].r.part1[16] );
tran (\sa_count[19][48] , \sa_count[19].f.upper[16] );
tran (\sa_count[19][49] , \sa_count[19].r.part1[17] );
tran (\sa_count[19][49] , \sa_count[19].f.upper[17] );
tran (\sa_count[19][50] , \sa_count[19].r.part1[18] );
tran (\sa_count[19][50] , \sa_count[19].f.unused[0] );
tran (\sa_count[19][51] , \sa_count[19].r.part1[19] );
tran (\sa_count[19][51] , \sa_count[19].f.unused[1] );
tran (\sa_count[19][52] , \sa_count[19].r.part1[20] );
tran (\sa_count[19][52] , \sa_count[19].f.unused[2] );
tran (\sa_count[19][53] , \sa_count[19].r.part1[21] );
tran (\sa_count[19][53] , \sa_count[19].f.unused[3] );
tran (\sa_count[19][54] , \sa_count[19].r.part1[22] );
tran (\sa_count[19][54] , \sa_count[19].f.unused[4] );
tran (\sa_count[19][55] , \sa_count[19].r.part1[23] );
tran (\sa_count[19][55] , \sa_count[19].f.unused[5] );
tran (\sa_count[19][56] , \sa_count[19].r.part1[24] );
tran (\sa_count[19][56] , \sa_count[19].f.unused[6] );
tran (\sa_count[19][57] , \sa_count[19].r.part1[25] );
tran (\sa_count[19][57] , \sa_count[19].f.unused[7] );
tran (\sa_count[19][58] , \sa_count[19].r.part1[26] );
tran (\sa_count[19][58] , \sa_count[19].f.unused[8] );
tran (\sa_count[19][59] , \sa_count[19].r.part1[27] );
tran (\sa_count[19][59] , \sa_count[19].f.unused[9] );
tran (\sa_count[19][60] , \sa_count[19].r.part1[28] );
tran (\sa_count[19][60] , \sa_count[19].f.unused[10] );
tran (\sa_count[19][61] , \sa_count[19].r.part1[29] );
tran (\sa_count[19][61] , \sa_count[19].f.unused[11] );
tran (\sa_count[19][62] , \sa_count[19].r.part1[30] );
tran (\sa_count[19][62] , \sa_count[19].f.unused[12] );
tran (\sa_count[19][63] , \sa_count[19].r.part1[31] );
tran (\sa_count[19][63] , \sa_count[19].f.unused[13] );
tran (\sa_count[20][0] , \sa_count[20].r.part0[0] );
tran (\sa_count[20][0] , \sa_count[20].f.lower[0] );
tran (\sa_count[20][1] , \sa_count[20].r.part0[1] );
tran (\sa_count[20][1] , \sa_count[20].f.lower[1] );
tran (\sa_count[20][2] , \sa_count[20].r.part0[2] );
tran (\sa_count[20][2] , \sa_count[20].f.lower[2] );
tran (\sa_count[20][3] , \sa_count[20].r.part0[3] );
tran (\sa_count[20][3] , \sa_count[20].f.lower[3] );
tran (\sa_count[20][4] , \sa_count[20].r.part0[4] );
tran (\sa_count[20][4] , \sa_count[20].f.lower[4] );
tran (\sa_count[20][5] , \sa_count[20].r.part0[5] );
tran (\sa_count[20][5] , \sa_count[20].f.lower[5] );
tran (\sa_count[20][6] , \sa_count[20].r.part0[6] );
tran (\sa_count[20][6] , \sa_count[20].f.lower[6] );
tran (\sa_count[20][7] , \sa_count[20].r.part0[7] );
tran (\sa_count[20][7] , \sa_count[20].f.lower[7] );
tran (\sa_count[20][8] , \sa_count[20].r.part0[8] );
tran (\sa_count[20][8] , \sa_count[20].f.lower[8] );
tran (\sa_count[20][9] , \sa_count[20].r.part0[9] );
tran (\sa_count[20][9] , \sa_count[20].f.lower[9] );
tran (\sa_count[20][10] , \sa_count[20].r.part0[10] );
tran (\sa_count[20][10] , \sa_count[20].f.lower[10] );
tran (\sa_count[20][11] , \sa_count[20].r.part0[11] );
tran (\sa_count[20][11] , \sa_count[20].f.lower[11] );
tran (\sa_count[20][12] , \sa_count[20].r.part0[12] );
tran (\sa_count[20][12] , \sa_count[20].f.lower[12] );
tran (\sa_count[20][13] , \sa_count[20].r.part0[13] );
tran (\sa_count[20][13] , \sa_count[20].f.lower[13] );
tran (\sa_count[20][14] , \sa_count[20].r.part0[14] );
tran (\sa_count[20][14] , \sa_count[20].f.lower[14] );
tran (\sa_count[20][15] , \sa_count[20].r.part0[15] );
tran (\sa_count[20][15] , \sa_count[20].f.lower[15] );
tran (\sa_count[20][16] , \sa_count[20].r.part0[16] );
tran (\sa_count[20][16] , \sa_count[20].f.lower[16] );
tran (\sa_count[20][17] , \sa_count[20].r.part0[17] );
tran (\sa_count[20][17] , \sa_count[20].f.lower[17] );
tran (\sa_count[20][18] , \sa_count[20].r.part0[18] );
tran (\sa_count[20][18] , \sa_count[20].f.lower[18] );
tran (\sa_count[20][19] , \sa_count[20].r.part0[19] );
tran (\sa_count[20][19] , \sa_count[20].f.lower[19] );
tran (\sa_count[20][20] , \sa_count[20].r.part0[20] );
tran (\sa_count[20][20] , \sa_count[20].f.lower[20] );
tran (\sa_count[20][21] , \sa_count[20].r.part0[21] );
tran (\sa_count[20][21] , \sa_count[20].f.lower[21] );
tran (\sa_count[20][22] , \sa_count[20].r.part0[22] );
tran (\sa_count[20][22] , \sa_count[20].f.lower[22] );
tran (\sa_count[20][23] , \sa_count[20].r.part0[23] );
tran (\sa_count[20][23] , \sa_count[20].f.lower[23] );
tran (\sa_count[20][24] , \sa_count[20].r.part0[24] );
tran (\sa_count[20][24] , \sa_count[20].f.lower[24] );
tran (\sa_count[20][25] , \sa_count[20].r.part0[25] );
tran (\sa_count[20][25] , \sa_count[20].f.lower[25] );
tran (\sa_count[20][26] , \sa_count[20].r.part0[26] );
tran (\sa_count[20][26] , \sa_count[20].f.lower[26] );
tran (\sa_count[20][27] , \sa_count[20].r.part0[27] );
tran (\sa_count[20][27] , \sa_count[20].f.lower[27] );
tran (\sa_count[20][28] , \sa_count[20].r.part0[28] );
tran (\sa_count[20][28] , \sa_count[20].f.lower[28] );
tran (\sa_count[20][29] , \sa_count[20].r.part0[29] );
tran (\sa_count[20][29] , \sa_count[20].f.lower[29] );
tran (\sa_count[20][30] , \sa_count[20].r.part0[30] );
tran (\sa_count[20][30] , \sa_count[20].f.lower[30] );
tran (\sa_count[20][31] , \sa_count[20].r.part0[31] );
tran (\sa_count[20][31] , \sa_count[20].f.lower[31] );
tran (\sa_count[20][32] , \sa_count[20].r.part1[0] );
tran (\sa_count[20][32] , \sa_count[20].f.upper[0] );
tran (\sa_count[20][33] , \sa_count[20].r.part1[1] );
tran (\sa_count[20][33] , \sa_count[20].f.upper[1] );
tran (\sa_count[20][34] , \sa_count[20].r.part1[2] );
tran (\sa_count[20][34] , \sa_count[20].f.upper[2] );
tran (\sa_count[20][35] , \sa_count[20].r.part1[3] );
tran (\sa_count[20][35] , \sa_count[20].f.upper[3] );
tran (\sa_count[20][36] , \sa_count[20].r.part1[4] );
tran (\sa_count[20][36] , \sa_count[20].f.upper[4] );
tran (\sa_count[20][37] , \sa_count[20].r.part1[5] );
tran (\sa_count[20][37] , \sa_count[20].f.upper[5] );
tran (\sa_count[20][38] , \sa_count[20].r.part1[6] );
tran (\sa_count[20][38] , \sa_count[20].f.upper[6] );
tran (\sa_count[20][39] , \sa_count[20].r.part1[7] );
tran (\sa_count[20][39] , \sa_count[20].f.upper[7] );
tran (\sa_count[20][40] , \sa_count[20].r.part1[8] );
tran (\sa_count[20][40] , \sa_count[20].f.upper[8] );
tran (\sa_count[20][41] , \sa_count[20].r.part1[9] );
tran (\sa_count[20][41] , \sa_count[20].f.upper[9] );
tran (\sa_count[20][42] , \sa_count[20].r.part1[10] );
tran (\sa_count[20][42] , \sa_count[20].f.upper[10] );
tran (\sa_count[20][43] , \sa_count[20].r.part1[11] );
tran (\sa_count[20][43] , \sa_count[20].f.upper[11] );
tran (\sa_count[20][44] , \sa_count[20].r.part1[12] );
tran (\sa_count[20][44] , \sa_count[20].f.upper[12] );
tran (\sa_count[20][45] , \sa_count[20].r.part1[13] );
tran (\sa_count[20][45] , \sa_count[20].f.upper[13] );
tran (\sa_count[20][46] , \sa_count[20].r.part1[14] );
tran (\sa_count[20][46] , \sa_count[20].f.upper[14] );
tran (\sa_count[20][47] , \sa_count[20].r.part1[15] );
tran (\sa_count[20][47] , \sa_count[20].f.upper[15] );
tran (\sa_count[20][48] , \sa_count[20].r.part1[16] );
tran (\sa_count[20][48] , \sa_count[20].f.upper[16] );
tran (\sa_count[20][49] , \sa_count[20].r.part1[17] );
tran (\sa_count[20][49] , \sa_count[20].f.upper[17] );
tran (\sa_count[20][50] , \sa_count[20].r.part1[18] );
tran (\sa_count[20][50] , \sa_count[20].f.unused[0] );
tran (\sa_count[20][51] , \sa_count[20].r.part1[19] );
tran (\sa_count[20][51] , \sa_count[20].f.unused[1] );
tran (\sa_count[20][52] , \sa_count[20].r.part1[20] );
tran (\sa_count[20][52] , \sa_count[20].f.unused[2] );
tran (\sa_count[20][53] , \sa_count[20].r.part1[21] );
tran (\sa_count[20][53] , \sa_count[20].f.unused[3] );
tran (\sa_count[20][54] , \sa_count[20].r.part1[22] );
tran (\sa_count[20][54] , \sa_count[20].f.unused[4] );
tran (\sa_count[20][55] , \sa_count[20].r.part1[23] );
tran (\sa_count[20][55] , \sa_count[20].f.unused[5] );
tran (\sa_count[20][56] , \sa_count[20].r.part1[24] );
tran (\sa_count[20][56] , \sa_count[20].f.unused[6] );
tran (\sa_count[20][57] , \sa_count[20].r.part1[25] );
tran (\sa_count[20][57] , \sa_count[20].f.unused[7] );
tran (\sa_count[20][58] , \sa_count[20].r.part1[26] );
tran (\sa_count[20][58] , \sa_count[20].f.unused[8] );
tran (\sa_count[20][59] , \sa_count[20].r.part1[27] );
tran (\sa_count[20][59] , \sa_count[20].f.unused[9] );
tran (\sa_count[20][60] , \sa_count[20].r.part1[28] );
tran (\sa_count[20][60] , \sa_count[20].f.unused[10] );
tran (\sa_count[20][61] , \sa_count[20].r.part1[29] );
tran (\sa_count[20][61] , \sa_count[20].f.unused[11] );
tran (\sa_count[20][62] , \sa_count[20].r.part1[30] );
tran (\sa_count[20][62] , \sa_count[20].f.unused[12] );
tran (\sa_count[20][63] , \sa_count[20].r.part1[31] );
tran (\sa_count[20][63] , \sa_count[20].f.unused[13] );
tran (\sa_count[21][0] , \sa_count[21].r.part0[0] );
tran (\sa_count[21][0] , \sa_count[21].f.lower[0] );
tran (\sa_count[21][1] , \sa_count[21].r.part0[1] );
tran (\sa_count[21][1] , \sa_count[21].f.lower[1] );
tran (\sa_count[21][2] , \sa_count[21].r.part0[2] );
tran (\sa_count[21][2] , \sa_count[21].f.lower[2] );
tran (\sa_count[21][3] , \sa_count[21].r.part0[3] );
tran (\sa_count[21][3] , \sa_count[21].f.lower[3] );
tran (\sa_count[21][4] , \sa_count[21].r.part0[4] );
tran (\sa_count[21][4] , \sa_count[21].f.lower[4] );
tran (\sa_count[21][5] , \sa_count[21].r.part0[5] );
tran (\sa_count[21][5] , \sa_count[21].f.lower[5] );
tran (\sa_count[21][6] , \sa_count[21].r.part0[6] );
tran (\sa_count[21][6] , \sa_count[21].f.lower[6] );
tran (\sa_count[21][7] , \sa_count[21].r.part0[7] );
tran (\sa_count[21][7] , \sa_count[21].f.lower[7] );
tran (\sa_count[21][8] , \sa_count[21].r.part0[8] );
tran (\sa_count[21][8] , \sa_count[21].f.lower[8] );
tran (\sa_count[21][9] , \sa_count[21].r.part0[9] );
tran (\sa_count[21][9] , \sa_count[21].f.lower[9] );
tran (\sa_count[21][10] , \sa_count[21].r.part0[10] );
tran (\sa_count[21][10] , \sa_count[21].f.lower[10] );
tran (\sa_count[21][11] , \sa_count[21].r.part0[11] );
tran (\sa_count[21][11] , \sa_count[21].f.lower[11] );
tran (\sa_count[21][12] , \sa_count[21].r.part0[12] );
tran (\sa_count[21][12] , \sa_count[21].f.lower[12] );
tran (\sa_count[21][13] , \sa_count[21].r.part0[13] );
tran (\sa_count[21][13] , \sa_count[21].f.lower[13] );
tran (\sa_count[21][14] , \sa_count[21].r.part0[14] );
tran (\sa_count[21][14] , \sa_count[21].f.lower[14] );
tran (\sa_count[21][15] , \sa_count[21].r.part0[15] );
tran (\sa_count[21][15] , \sa_count[21].f.lower[15] );
tran (\sa_count[21][16] , \sa_count[21].r.part0[16] );
tran (\sa_count[21][16] , \sa_count[21].f.lower[16] );
tran (\sa_count[21][17] , \sa_count[21].r.part0[17] );
tran (\sa_count[21][17] , \sa_count[21].f.lower[17] );
tran (\sa_count[21][18] , \sa_count[21].r.part0[18] );
tran (\sa_count[21][18] , \sa_count[21].f.lower[18] );
tran (\sa_count[21][19] , \sa_count[21].r.part0[19] );
tran (\sa_count[21][19] , \sa_count[21].f.lower[19] );
tran (\sa_count[21][20] , \sa_count[21].r.part0[20] );
tran (\sa_count[21][20] , \sa_count[21].f.lower[20] );
tran (\sa_count[21][21] , \sa_count[21].r.part0[21] );
tran (\sa_count[21][21] , \sa_count[21].f.lower[21] );
tran (\sa_count[21][22] , \sa_count[21].r.part0[22] );
tran (\sa_count[21][22] , \sa_count[21].f.lower[22] );
tran (\sa_count[21][23] , \sa_count[21].r.part0[23] );
tran (\sa_count[21][23] , \sa_count[21].f.lower[23] );
tran (\sa_count[21][24] , \sa_count[21].r.part0[24] );
tran (\sa_count[21][24] , \sa_count[21].f.lower[24] );
tran (\sa_count[21][25] , \sa_count[21].r.part0[25] );
tran (\sa_count[21][25] , \sa_count[21].f.lower[25] );
tran (\sa_count[21][26] , \sa_count[21].r.part0[26] );
tran (\sa_count[21][26] , \sa_count[21].f.lower[26] );
tran (\sa_count[21][27] , \sa_count[21].r.part0[27] );
tran (\sa_count[21][27] , \sa_count[21].f.lower[27] );
tran (\sa_count[21][28] , \sa_count[21].r.part0[28] );
tran (\sa_count[21][28] , \sa_count[21].f.lower[28] );
tran (\sa_count[21][29] , \sa_count[21].r.part0[29] );
tran (\sa_count[21][29] , \sa_count[21].f.lower[29] );
tran (\sa_count[21][30] , \sa_count[21].r.part0[30] );
tran (\sa_count[21][30] , \sa_count[21].f.lower[30] );
tran (\sa_count[21][31] , \sa_count[21].r.part0[31] );
tran (\sa_count[21][31] , \sa_count[21].f.lower[31] );
tran (\sa_count[21][32] , \sa_count[21].r.part1[0] );
tran (\sa_count[21][32] , \sa_count[21].f.upper[0] );
tran (\sa_count[21][33] , \sa_count[21].r.part1[1] );
tran (\sa_count[21][33] , \sa_count[21].f.upper[1] );
tran (\sa_count[21][34] , \sa_count[21].r.part1[2] );
tran (\sa_count[21][34] , \sa_count[21].f.upper[2] );
tran (\sa_count[21][35] , \sa_count[21].r.part1[3] );
tran (\sa_count[21][35] , \sa_count[21].f.upper[3] );
tran (\sa_count[21][36] , \sa_count[21].r.part1[4] );
tran (\sa_count[21][36] , \sa_count[21].f.upper[4] );
tran (\sa_count[21][37] , \sa_count[21].r.part1[5] );
tran (\sa_count[21][37] , \sa_count[21].f.upper[5] );
tran (\sa_count[21][38] , \sa_count[21].r.part1[6] );
tran (\sa_count[21][38] , \sa_count[21].f.upper[6] );
tran (\sa_count[21][39] , \sa_count[21].r.part1[7] );
tran (\sa_count[21][39] , \sa_count[21].f.upper[7] );
tran (\sa_count[21][40] , \sa_count[21].r.part1[8] );
tran (\sa_count[21][40] , \sa_count[21].f.upper[8] );
tran (\sa_count[21][41] , \sa_count[21].r.part1[9] );
tran (\sa_count[21][41] , \sa_count[21].f.upper[9] );
tran (\sa_count[21][42] , \sa_count[21].r.part1[10] );
tran (\sa_count[21][42] , \sa_count[21].f.upper[10] );
tran (\sa_count[21][43] , \sa_count[21].r.part1[11] );
tran (\sa_count[21][43] , \sa_count[21].f.upper[11] );
tran (\sa_count[21][44] , \sa_count[21].r.part1[12] );
tran (\sa_count[21][44] , \sa_count[21].f.upper[12] );
tran (\sa_count[21][45] , \sa_count[21].r.part1[13] );
tran (\sa_count[21][45] , \sa_count[21].f.upper[13] );
tran (\sa_count[21][46] , \sa_count[21].r.part1[14] );
tran (\sa_count[21][46] , \sa_count[21].f.upper[14] );
tran (\sa_count[21][47] , \sa_count[21].r.part1[15] );
tran (\sa_count[21][47] , \sa_count[21].f.upper[15] );
tran (\sa_count[21][48] , \sa_count[21].r.part1[16] );
tran (\sa_count[21][48] , \sa_count[21].f.upper[16] );
tran (\sa_count[21][49] , \sa_count[21].r.part1[17] );
tran (\sa_count[21][49] , \sa_count[21].f.upper[17] );
tran (\sa_count[21][50] , \sa_count[21].r.part1[18] );
tran (\sa_count[21][50] , \sa_count[21].f.unused[0] );
tran (\sa_count[21][51] , \sa_count[21].r.part1[19] );
tran (\sa_count[21][51] , \sa_count[21].f.unused[1] );
tran (\sa_count[21][52] , \sa_count[21].r.part1[20] );
tran (\sa_count[21][52] , \sa_count[21].f.unused[2] );
tran (\sa_count[21][53] , \sa_count[21].r.part1[21] );
tran (\sa_count[21][53] , \sa_count[21].f.unused[3] );
tran (\sa_count[21][54] , \sa_count[21].r.part1[22] );
tran (\sa_count[21][54] , \sa_count[21].f.unused[4] );
tran (\sa_count[21][55] , \sa_count[21].r.part1[23] );
tran (\sa_count[21][55] , \sa_count[21].f.unused[5] );
tran (\sa_count[21][56] , \sa_count[21].r.part1[24] );
tran (\sa_count[21][56] , \sa_count[21].f.unused[6] );
tran (\sa_count[21][57] , \sa_count[21].r.part1[25] );
tran (\sa_count[21][57] , \sa_count[21].f.unused[7] );
tran (\sa_count[21][58] , \sa_count[21].r.part1[26] );
tran (\sa_count[21][58] , \sa_count[21].f.unused[8] );
tran (\sa_count[21][59] , \sa_count[21].r.part1[27] );
tran (\sa_count[21][59] , \sa_count[21].f.unused[9] );
tran (\sa_count[21][60] , \sa_count[21].r.part1[28] );
tran (\sa_count[21][60] , \sa_count[21].f.unused[10] );
tran (\sa_count[21][61] , \sa_count[21].r.part1[29] );
tran (\sa_count[21][61] , \sa_count[21].f.unused[11] );
tran (\sa_count[21][62] , \sa_count[21].r.part1[30] );
tran (\sa_count[21][62] , \sa_count[21].f.unused[12] );
tran (\sa_count[21][63] , \sa_count[21].r.part1[31] );
tran (\sa_count[21][63] , \sa_count[21].f.unused[13] );
tran (\sa_count[22][0] , \sa_count[22].r.part0[0] );
tran (\sa_count[22][0] , \sa_count[22].f.lower[0] );
tran (\sa_count[22][1] , \sa_count[22].r.part0[1] );
tran (\sa_count[22][1] , \sa_count[22].f.lower[1] );
tran (\sa_count[22][2] , \sa_count[22].r.part0[2] );
tran (\sa_count[22][2] , \sa_count[22].f.lower[2] );
tran (\sa_count[22][3] , \sa_count[22].r.part0[3] );
tran (\sa_count[22][3] , \sa_count[22].f.lower[3] );
tran (\sa_count[22][4] , \sa_count[22].r.part0[4] );
tran (\sa_count[22][4] , \sa_count[22].f.lower[4] );
tran (\sa_count[22][5] , \sa_count[22].r.part0[5] );
tran (\sa_count[22][5] , \sa_count[22].f.lower[5] );
tran (\sa_count[22][6] , \sa_count[22].r.part0[6] );
tran (\sa_count[22][6] , \sa_count[22].f.lower[6] );
tran (\sa_count[22][7] , \sa_count[22].r.part0[7] );
tran (\sa_count[22][7] , \sa_count[22].f.lower[7] );
tran (\sa_count[22][8] , \sa_count[22].r.part0[8] );
tran (\sa_count[22][8] , \sa_count[22].f.lower[8] );
tran (\sa_count[22][9] , \sa_count[22].r.part0[9] );
tran (\sa_count[22][9] , \sa_count[22].f.lower[9] );
tran (\sa_count[22][10] , \sa_count[22].r.part0[10] );
tran (\sa_count[22][10] , \sa_count[22].f.lower[10] );
tran (\sa_count[22][11] , \sa_count[22].r.part0[11] );
tran (\sa_count[22][11] , \sa_count[22].f.lower[11] );
tran (\sa_count[22][12] , \sa_count[22].r.part0[12] );
tran (\sa_count[22][12] , \sa_count[22].f.lower[12] );
tran (\sa_count[22][13] , \sa_count[22].r.part0[13] );
tran (\sa_count[22][13] , \sa_count[22].f.lower[13] );
tran (\sa_count[22][14] , \sa_count[22].r.part0[14] );
tran (\sa_count[22][14] , \sa_count[22].f.lower[14] );
tran (\sa_count[22][15] , \sa_count[22].r.part0[15] );
tran (\sa_count[22][15] , \sa_count[22].f.lower[15] );
tran (\sa_count[22][16] , \sa_count[22].r.part0[16] );
tran (\sa_count[22][16] , \sa_count[22].f.lower[16] );
tran (\sa_count[22][17] , \sa_count[22].r.part0[17] );
tran (\sa_count[22][17] , \sa_count[22].f.lower[17] );
tran (\sa_count[22][18] , \sa_count[22].r.part0[18] );
tran (\sa_count[22][18] , \sa_count[22].f.lower[18] );
tran (\sa_count[22][19] , \sa_count[22].r.part0[19] );
tran (\sa_count[22][19] , \sa_count[22].f.lower[19] );
tran (\sa_count[22][20] , \sa_count[22].r.part0[20] );
tran (\sa_count[22][20] , \sa_count[22].f.lower[20] );
tran (\sa_count[22][21] , \sa_count[22].r.part0[21] );
tran (\sa_count[22][21] , \sa_count[22].f.lower[21] );
tran (\sa_count[22][22] , \sa_count[22].r.part0[22] );
tran (\sa_count[22][22] , \sa_count[22].f.lower[22] );
tran (\sa_count[22][23] , \sa_count[22].r.part0[23] );
tran (\sa_count[22][23] , \sa_count[22].f.lower[23] );
tran (\sa_count[22][24] , \sa_count[22].r.part0[24] );
tran (\sa_count[22][24] , \sa_count[22].f.lower[24] );
tran (\sa_count[22][25] , \sa_count[22].r.part0[25] );
tran (\sa_count[22][25] , \sa_count[22].f.lower[25] );
tran (\sa_count[22][26] , \sa_count[22].r.part0[26] );
tran (\sa_count[22][26] , \sa_count[22].f.lower[26] );
tran (\sa_count[22][27] , \sa_count[22].r.part0[27] );
tran (\sa_count[22][27] , \sa_count[22].f.lower[27] );
tran (\sa_count[22][28] , \sa_count[22].r.part0[28] );
tran (\sa_count[22][28] , \sa_count[22].f.lower[28] );
tran (\sa_count[22][29] , \sa_count[22].r.part0[29] );
tran (\sa_count[22][29] , \sa_count[22].f.lower[29] );
tran (\sa_count[22][30] , \sa_count[22].r.part0[30] );
tran (\sa_count[22][30] , \sa_count[22].f.lower[30] );
tran (\sa_count[22][31] , \sa_count[22].r.part0[31] );
tran (\sa_count[22][31] , \sa_count[22].f.lower[31] );
tran (\sa_count[22][32] , \sa_count[22].r.part1[0] );
tran (\sa_count[22][32] , \sa_count[22].f.upper[0] );
tran (\sa_count[22][33] , \sa_count[22].r.part1[1] );
tran (\sa_count[22][33] , \sa_count[22].f.upper[1] );
tran (\sa_count[22][34] , \sa_count[22].r.part1[2] );
tran (\sa_count[22][34] , \sa_count[22].f.upper[2] );
tran (\sa_count[22][35] , \sa_count[22].r.part1[3] );
tran (\sa_count[22][35] , \sa_count[22].f.upper[3] );
tran (\sa_count[22][36] , \sa_count[22].r.part1[4] );
tran (\sa_count[22][36] , \sa_count[22].f.upper[4] );
tran (\sa_count[22][37] , \sa_count[22].r.part1[5] );
tran (\sa_count[22][37] , \sa_count[22].f.upper[5] );
tran (\sa_count[22][38] , \sa_count[22].r.part1[6] );
tran (\sa_count[22][38] , \sa_count[22].f.upper[6] );
tran (\sa_count[22][39] , \sa_count[22].r.part1[7] );
tran (\sa_count[22][39] , \sa_count[22].f.upper[7] );
tran (\sa_count[22][40] , \sa_count[22].r.part1[8] );
tran (\sa_count[22][40] , \sa_count[22].f.upper[8] );
tran (\sa_count[22][41] , \sa_count[22].r.part1[9] );
tran (\sa_count[22][41] , \sa_count[22].f.upper[9] );
tran (\sa_count[22][42] , \sa_count[22].r.part1[10] );
tran (\sa_count[22][42] , \sa_count[22].f.upper[10] );
tran (\sa_count[22][43] , \sa_count[22].r.part1[11] );
tran (\sa_count[22][43] , \sa_count[22].f.upper[11] );
tran (\sa_count[22][44] , \sa_count[22].r.part1[12] );
tran (\sa_count[22][44] , \sa_count[22].f.upper[12] );
tran (\sa_count[22][45] , \sa_count[22].r.part1[13] );
tran (\sa_count[22][45] , \sa_count[22].f.upper[13] );
tran (\sa_count[22][46] , \sa_count[22].r.part1[14] );
tran (\sa_count[22][46] , \sa_count[22].f.upper[14] );
tran (\sa_count[22][47] , \sa_count[22].r.part1[15] );
tran (\sa_count[22][47] , \sa_count[22].f.upper[15] );
tran (\sa_count[22][48] , \sa_count[22].r.part1[16] );
tran (\sa_count[22][48] , \sa_count[22].f.upper[16] );
tran (\sa_count[22][49] , \sa_count[22].r.part1[17] );
tran (\sa_count[22][49] , \sa_count[22].f.upper[17] );
tran (\sa_count[22][50] , \sa_count[22].r.part1[18] );
tran (\sa_count[22][50] , \sa_count[22].f.unused[0] );
tran (\sa_count[22][51] , \sa_count[22].r.part1[19] );
tran (\sa_count[22][51] , \sa_count[22].f.unused[1] );
tran (\sa_count[22][52] , \sa_count[22].r.part1[20] );
tran (\sa_count[22][52] , \sa_count[22].f.unused[2] );
tran (\sa_count[22][53] , \sa_count[22].r.part1[21] );
tran (\sa_count[22][53] , \sa_count[22].f.unused[3] );
tran (\sa_count[22][54] , \sa_count[22].r.part1[22] );
tran (\sa_count[22][54] , \sa_count[22].f.unused[4] );
tran (\sa_count[22][55] , \sa_count[22].r.part1[23] );
tran (\sa_count[22][55] , \sa_count[22].f.unused[5] );
tran (\sa_count[22][56] , \sa_count[22].r.part1[24] );
tran (\sa_count[22][56] , \sa_count[22].f.unused[6] );
tran (\sa_count[22][57] , \sa_count[22].r.part1[25] );
tran (\sa_count[22][57] , \sa_count[22].f.unused[7] );
tran (\sa_count[22][58] , \sa_count[22].r.part1[26] );
tran (\sa_count[22][58] , \sa_count[22].f.unused[8] );
tran (\sa_count[22][59] , \sa_count[22].r.part1[27] );
tran (\sa_count[22][59] , \sa_count[22].f.unused[9] );
tran (\sa_count[22][60] , \sa_count[22].r.part1[28] );
tran (\sa_count[22][60] , \sa_count[22].f.unused[10] );
tran (\sa_count[22][61] , \sa_count[22].r.part1[29] );
tran (\sa_count[22][61] , \sa_count[22].f.unused[11] );
tran (\sa_count[22][62] , \sa_count[22].r.part1[30] );
tran (\sa_count[22][62] , \sa_count[22].f.unused[12] );
tran (\sa_count[22][63] , \sa_count[22].r.part1[31] );
tran (\sa_count[22][63] , \sa_count[22].f.unused[13] );
tran (\sa_count[23][0] , \sa_count[23].r.part0[0] );
tran (\sa_count[23][0] , \sa_count[23].f.lower[0] );
tran (\sa_count[23][1] , \sa_count[23].r.part0[1] );
tran (\sa_count[23][1] , \sa_count[23].f.lower[1] );
tran (\sa_count[23][2] , \sa_count[23].r.part0[2] );
tran (\sa_count[23][2] , \sa_count[23].f.lower[2] );
tran (\sa_count[23][3] , \sa_count[23].r.part0[3] );
tran (\sa_count[23][3] , \sa_count[23].f.lower[3] );
tran (\sa_count[23][4] , \sa_count[23].r.part0[4] );
tran (\sa_count[23][4] , \sa_count[23].f.lower[4] );
tran (\sa_count[23][5] , \sa_count[23].r.part0[5] );
tran (\sa_count[23][5] , \sa_count[23].f.lower[5] );
tran (\sa_count[23][6] , \sa_count[23].r.part0[6] );
tran (\sa_count[23][6] , \sa_count[23].f.lower[6] );
tran (\sa_count[23][7] , \sa_count[23].r.part0[7] );
tran (\sa_count[23][7] , \sa_count[23].f.lower[7] );
tran (\sa_count[23][8] , \sa_count[23].r.part0[8] );
tran (\sa_count[23][8] , \sa_count[23].f.lower[8] );
tran (\sa_count[23][9] , \sa_count[23].r.part0[9] );
tran (\sa_count[23][9] , \sa_count[23].f.lower[9] );
tran (\sa_count[23][10] , \sa_count[23].r.part0[10] );
tran (\sa_count[23][10] , \sa_count[23].f.lower[10] );
tran (\sa_count[23][11] , \sa_count[23].r.part0[11] );
tran (\sa_count[23][11] , \sa_count[23].f.lower[11] );
tran (\sa_count[23][12] , \sa_count[23].r.part0[12] );
tran (\sa_count[23][12] , \sa_count[23].f.lower[12] );
tran (\sa_count[23][13] , \sa_count[23].r.part0[13] );
tran (\sa_count[23][13] , \sa_count[23].f.lower[13] );
tran (\sa_count[23][14] , \sa_count[23].r.part0[14] );
tran (\sa_count[23][14] , \sa_count[23].f.lower[14] );
tran (\sa_count[23][15] , \sa_count[23].r.part0[15] );
tran (\sa_count[23][15] , \sa_count[23].f.lower[15] );
tran (\sa_count[23][16] , \sa_count[23].r.part0[16] );
tran (\sa_count[23][16] , \sa_count[23].f.lower[16] );
tran (\sa_count[23][17] , \sa_count[23].r.part0[17] );
tran (\sa_count[23][17] , \sa_count[23].f.lower[17] );
tran (\sa_count[23][18] , \sa_count[23].r.part0[18] );
tran (\sa_count[23][18] , \sa_count[23].f.lower[18] );
tran (\sa_count[23][19] , \sa_count[23].r.part0[19] );
tran (\sa_count[23][19] , \sa_count[23].f.lower[19] );
tran (\sa_count[23][20] , \sa_count[23].r.part0[20] );
tran (\sa_count[23][20] , \sa_count[23].f.lower[20] );
tran (\sa_count[23][21] , \sa_count[23].r.part0[21] );
tran (\sa_count[23][21] , \sa_count[23].f.lower[21] );
tran (\sa_count[23][22] , \sa_count[23].r.part0[22] );
tran (\sa_count[23][22] , \sa_count[23].f.lower[22] );
tran (\sa_count[23][23] , \sa_count[23].r.part0[23] );
tran (\sa_count[23][23] , \sa_count[23].f.lower[23] );
tran (\sa_count[23][24] , \sa_count[23].r.part0[24] );
tran (\sa_count[23][24] , \sa_count[23].f.lower[24] );
tran (\sa_count[23][25] , \sa_count[23].r.part0[25] );
tran (\sa_count[23][25] , \sa_count[23].f.lower[25] );
tran (\sa_count[23][26] , \sa_count[23].r.part0[26] );
tran (\sa_count[23][26] , \sa_count[23].f.lower[26] );
tran (\sa_count[23][27] , \sa_count[23].r.part0[27] );
tran (\sa_count[23][27] , \sa_count[23].f.lower[27] );
tran (\sa_count[23][28] , \sa_count[23].r.part0[28] );
tran (\sa_count[23][28] , \sa_count[23].f.lower[28] );
tran (\sa_count[23][29] , \sa_count[23].r.part0[29] );
tran (\sa_count[23][29] , \sa_count[23].f.lower[29] );
tran (\sa_count[23][30] , \sa_count[23].r.part0[30] );
tran (\sa_count[23][30] , \sa_count[23].f.lower[30] );
tran (\sa_count[23][31] , \sa_count[23].r.part0[31] );
tran (\sa_count[23][31] , \sa_count[23].f.lower[31] );
tran (\sa_count[23][32] , \sa_count[23].r.part1[0] );
tran (\sa_count[23][32] , \sa_count[23].f.upper[0] );
tran (\sa_count[23][33] , \sa_count[23].r.part1[1] );
tran (\sa_count[23][33] , \sa_count[23].f.upper[1] );
tran (\sa_count[23][34] , \sa_count[23].r.part1[2] );
tran (\sa_count[23][34] , \sa_count[23].f.upper[2] );
tran (\sa_count[23][35] , \sa_count[23].r.part1[3] );
tran (\sa_count[23][35] , \sa_count[23].f.upper[3] );
tran (\sa_count[23][36] , \sa_count[23].r.part1[4] );
tran (\sa_count[23][36] , \sa_count[23].f.upper[4] );
tran (\sa_count[23][37] , \sa_count[23].r.part1[5] );
tran (\sa_count[23][37] , \sa_count[23].f.upper[5] );
tran (\sa_count[23][38] , \sa_count[23].r.part1[6] );
tran (\sa_count[23][38] , \sa_count[23].f.upper[6] );
tran (\sa_count[23][39] , \sa_count[23].r.part1[7] );
tran (\sa_count[23][39] , \sa_count[23].f.upper[7] );
tran (\sa_count[23][40] , \sa_count[23].r.part1[8] );
tran (\sa_count[23][40] , \sa_count[23].f.upper[8] );
tran (\sa_count[23][41] , \sa_count[23].r.part1[9] );
tran (\sa_count[23][41] , \sa_count[23].f.upper[9] );
tran (\sa_count[23][42] , \sa_count[23].r.part1[10] );
tran (\sa_count[23][42] , \sa_count[23].f.upper[10] );
tran (\sa_count[23][43] , \sa_count[23].r.part1[11] );
tran (\sa_count[23][43] , \sa_count[23].f.upper[11] );
tran (\sa_count[23][44] , \sa_count[23].r.part1[12] );
tran (\sa_count[23][44] , \sa_count[23].f.upper[12] );
tran (\sa_count[23][45] , \sa_count[23].r.part1[13] );
tran (\sa_count[23][45] , \sa_count[23].f.upper[13] );
tran (\sa_count[23][46] , \sa_count[23].r.part1[14] );
tran (\sa_count[23][46] , \sa_count[23].f.upper[14] );
tran (\sa_count[23][47] , \sa_count[23].r.part1[15] );
tran (\sa_count[23][47] , \sa_count[23].f.upper[15] );
tran (\sa_count[23][48] , \sa_count[23].r.part1[16] );
tran (\sa_count[23][48] , \sa_count[23].f.upper[16] );
tran (\sa_count[23][49] , \sa_count[23].r.part1[17] );
tran (\sa_count[23][49] , \sa_count[23].f.upper[17] );
tran (\sa_count[23][50] , \sa_count[23].r.part1[18] );
tran (\sa_count[23][50] , \sa_count[23].f.unused[0] );
tran (\sa_count[23][51] , \sa_count[23].r.part1[19] );
tran (\sa_count[23][51] , \sa_count[23].f.unused[1] );
tran (\sa_count[23][52] , \sa_count[23].r.part1[20] );
tran (\sa_count[23][52] , \sa_count[23].f.unused[2] );
tran (\sa_count[23][53] , \sa_count[23].r.part1[21] );
tran (\sa_count[23][53] , \sa_count[23].f.unused[3] );
tran (\sa_count[23][54] , \sa_count[23].r.part1[22] );
tran (\sa_count[23][54] , \sa_count[23].f.unused[4] );
tran (\sa_count[23][55] , \sa_count[23].r.part1[23] );
tran (\sa_count[23][55] , \sa_count[23].f.unused[5] );
tran (\sa_count[23][56] , \sa_count[23].r.part1[24] );
tran (\sa_count[23][56] , \sa_count[23].f.unused[6] );
tran (\sa_count[23][57] , \sa_count[23].r.part1[25] );
tran (\sa_count[23][57] , \sa_count[23].f.unused[7] );
tran (\sa_count[23][58] , \sa_count[23].r.part1[26] );
tran (\sa_count[23][58] , \sa_count[23].f.unused[8] );
tran (\sa_count[23][59] , \sa_count[23].r.part1[27] );
tran (\sa_count[23][59] , \sa_count[23].f.unused[9] );
tran (\sa_count[23][60] , \sa_count[23].r.part1[28] );
tran (\sa_count[23][60] , \sa_count[23].f.unused[10] );
tran (\sa_count[23][61] , \sa_count[23].r.part1[29] );
tran (\sa_count[23][61] , \sa_count[23].f.unused[11] );
tran (\sa_count[23][62] , \sa_count[23].r.part1[30] );
tran (\sa_count[23][62] , \sa_count[23].f.unused[12] );
tran (\sa_count[23][63] , \sa_count[23].r.part1[31] );
tran (\sa_count[23][63] , \sa_count[23].f.unused[13] );
tran (\sa_count[24][0] , \sa_count[24].r.part0[0] );
tran (\sa_count[24][0] , \sa_count[24].f.lower[0] );
tran (\sa_count[24][1] , \sa_count[24].r.part0[1] );
tran (\sa_count[24][1] , \sa_count[24].f.lower[1] );
tran (\sa_count[24][2] , \sa_count[24].r.part0[2] );
tran (\sa_count[24][2] , \sa_count[24].f.lower[2] );
tran (\sa_count[24][3] , \sa_count[24].r.part0[3] );
tran (\sa_count[24][3] , \sa_count[24].f.lower[3] );
tran (\sa_count[24][4] , \sa_count[24].r.part0[4] );
tran (\sa_count[24][4] , \sa_count[24].f.lower[4] );
tran (\sa_count[24][5] , \sa_count[24].r.part0[5] );
tran (\sa_count[24][5] , \sa_count[24].f.lower[5] );
tran (\sa_count[24][6] , \sa_count[24].r.part0[6] );
tran (\sa_count[24][6] , \sa_count[24].f.lower[6] );
tran (\sa_count[24][7] , \sa_count[24].r.part0[7] );
tran (\sa_count[24][7] , \sa_count[24].f.lower[7] );
tran (\sa_count[24][8] , \sa_count[24].r.part0[8] );
tran (\sa_count[24][8] , \sa_count[24].f.lower[8] );
tran (\sa_count[24][9] , \sa_count[24].r.part0[9] );
tran (\sa_count[24][9] , \sa_count[24].f.lower[9] );
tran (\sa_count[24][10] , \sa_count[24].r.part0[10] );
tran (\sa_count[24][10] , \sa_count[24].f.lower[10] );
tran (\sa_count[24][11] , \sa_count[24].r.part0[11] );
tran (\sa_count[24][11] , \sa_count[24].f.lower[11] );
tran (\sa_count[24][12] , \sa_count[24].r.part0[12] );
tran (\sa_count[24][12] , \sa_count[24].f.lower[12] );
tran (\sa_count[24][13] , \sa_count[24].r.part0[13] );
tran (\sa_count[24][13] , \sa_count[24].f.lower[13] );
tran (\sa_count[24][14] , \sa_count[24].r.part0[14] );
tran (\sa_count[24][14] , \sa_count[24].f.lower[14] );
tran (\sa_count[24][15] , \sa_count[24].r.part0[15] );
tran (\sa_count[24][15] , \sa_count[24].f.lower[15] );
tran (\sa_count[24][16] , \sa_count[24].r.part0[16] );
tran (\sa_count[24][16] , \sa_count[24].f.lower[16] );
tran (\sa_count[24][17] , \sa_count[24].r.part0[17] );
tran (\sa_count[24][17] , \sa_count[24].f.lower[17] );
tran (\sa_count[24][18] , \sa_count[24].r.part0[18] );
tran (\sa_count[24][18] , \sa_count[24].f.lower[18] );
tran (\sa_count[24][19] , \sa_count[24].r.part0[19] );
tran (\sa_count[24][19] , \sa_count[24].f.lower[19] );
tran (\sa_count[24][20] , \sa_count[24].r.part0[20] );
tran (\sa_count[24][20] , \sa_count[24].f.lower[20] );
tran (\sa_count[24][21] , \sa_count[24].r.part0[21] );
tran (\sa_count[24][21] , \sa_count[24].f.lower[21] );
tran (\sa_count[24][22] , \sa_count[24].r.part0[22] );
tran (\sa_count[24][22] , \sa_count[24].f.lower[22] );
tran (\sa_count[24][23] , \sa_count[24].r.part0[23] );
tran (\sa_count[24][23] , \sa_count[24].f.lower[23] );
tran (\sa_count[24][24] , \sa_count[24].r.part0[24] );
tran (\sa_count[24][24] , \sa_count[24].f.lower[24] );
tran (\sa_count[24][25] , \sa_count[24].r.part0[25] );
tran (\sa_count[24][25] , \sa_count[24].f.lower[25] );
tran (\sa_count[24][26] , \sa_count[24].r.part0[26] );
tran (\sa_count[24][26] , \sa_count[24].f.lower[26] );
tran (\sa_count[24][27] , \sa_count[24].r.part0[27] );
tran (\sa_count[24][27] , \sa_count[24].f.lower[27] );
tran (\sa_count[24][28] , \sa_count[24].r.part0[28] );
tran (\sa_count[24][28] , \sa_count[24].f.lower[28] );
tran (\sa_count[24][29] , \sa_count[24].r.part0[29] );
tran (\sa_count[24][29] , \sa_count[24].f.lower[29] );
tran (\sa_count[24][30] , \sa_count[24].r.part0[30] );
tran (\sa_count[24][30] , \sa_count[24].f.lower[30] );
tran (\sa_count[24][31] , \sa_count[24].r.part0[31] );
tran (\sa_count[24][31] , \sa_count[24].f.lower[31] );
tran (\sa_count[24][32] , \sa_count[24].r.part1[0] );
tran (\sa_count[24][32] , \sa_count[24].f.upper[0] );
tran (\sa_count[24][33] , \sa_count[24].r.part1[1] );
tran (\sa_count[24][33] , \sa_count[24].f.upper[1] );
tran (\sa_count[24][34] , \sa_count[24].r.part1[2] );
tran (\sa_count[24][34] , \sa_count[24].f.upper[2] );
tran (\sa_count[24][35] , \sa_count[24].r.part1[3] );
tran (\sa_count[24][35] , \sa_count[24].f.upper[3] );
tran (\sa_count[24][36] , \sa_count[24].r.part1[4] );
tran (\sa_count[24][36] , \sa_count[24].f.upper[4] );
tran (\sa_count[24][37] , \sa_count[24].r.part1[5] );
tran (\sa_count[24][37] , \sa_count[24].f.upper[5] );
tran (\sa_count[24][38] , \sa_count[24].r.part1[6] );
tran (\sa_count[24][38] , \sa_count[24].f.upper[6] );
tran (\sa_count[24][39] , \sa_count[24].r.part1[7] );
tran (\sa_count[24][39] , \sa_count[24].f.upper[7] );
tran (\sa_count[24][40] , \sa_count[24].r.part1[8] );
tran (\sa_count[24][40] , \sa_count[24].f.upper[8] );
tran (\sa_count[24][41] , \sa_count[24].r.part1[9] );
tran (\sa_count[24][41] , \sa_count[24].f.upper[9] );
tran (\sa_count[24][42] , \sa_count[24].r.part1[10] );
tran (\sa_count[24][42] , \sa_count[24].f.upper[10] );
tran (\sa_count[24][43] , \sa_count[24].r.part1[11] );
tran (\sa_count[24][43] , \sa_count[24].f.upper[11] );
tran (\sa_count[24][44] , \sa_count[24].r.part1[12] );
tran (\sa_count[24][44] , \sa_count[24].f.upper[12] );
tran (\sa_count[24][45] , \sa_count[24].r.part1[13] );
tran (\sa_count[24][45] , \sa_count[24].f.upper[13] );
tran (\sa_count[24][46] , \sa_count[24].r.part1[14] );
tran (\sa_count[24][46] , \sa_count[24].f.upper[14] );
tran (\sa_count[24][47] , \sa_count[24].r.part1[15] );
tran (\sa_count[24][47] , \sa_count[24].f.upper[15] );
tran (\sa_count[24][48] , \sa_count[24].r.part1[16] );
tran (\sa_count[24][48] , \sa_count[24].f.upper[16] );
tran (\sa_count[24][49] , \sa_count[24].r.part1[17] );
tran (\sa_count[24][49] , \sa_count[24].f.upper[17] );
tran (\sa_count[24][50] , \sa_count[24].r.part1[18] );
tran (\sa_count[24][50] , \sa_count[24].f.unused[0] );
tran (\sa_count[24][51] , \sa_count[24].r.part1[19] );
tran (\sa_count[24][51] , \sa_count[24].f.unused[1] );
tran (\sa_count[24][52] , \sa_count[24].r.part1[20] );
tran (\sa_count[24][52] , \sa_count[24].f.unused[2] );
tran (\sa_count[24][53] , \sa_count[24].r.part1[21] );
tran (\sa_count[24][53] , \sa_count[24].f.unused[3] );
tran (\sa_count[24][54] , \sa_count[24].r.part1[22] );
tran (\sa_count[24][54] , \sa_count[24].f.unused[4] );
tran (\sa_count[24][55] , \sa_count[24].r.part1[23] );
tran (\sa_count[24][55] , \sa_count[24].f.unused[5] );
tran (\sa_count[24][56] , \sa_count[24].r.part1[24] );
tran (\sa_count[24][56] , \sa_count[24].f.unused[6] );
tran (\sa_count[24][57] , \sa_count[24].r.part1[25] );
tran (\sa_count[24][57] , \sa_count[24].f.unused[7] );
tran (\sa_count[24][58] , \sa_count[24].r.part1[26] );
tran (\sa_count[24][58] , \sa_count[24].f.unused[8] );
tran (\sa_count[24][59] , \sa_count[24].r.part1[27] );
tran (\sa_count[24][59] , \sa_count[24].f.unused[9] );
tran (\sa_count[24][60] , \sa_count[24].r.part1[28] );
tran (\sa_count[24][60] , \sa_count[24].f.unused[10] );
tran (\sa_count[24][61] , \sa_count[24].r.part1[29] );
tran (\sa_count[24][61] , \sa_count[24].f.unused[11] );
tran (\sa_count[24][62] , \sa_count[24].r.part1[30] );
tran (\sa_count[24][62] , \sa_count[24].f.unused[12] );
tran (\sa_count[24][63] , \sa_count[24].r.part1[31] );
tran (\sa_count[24][63] , \sa_count[24].f.unused[13] );
tran (\sa_count[25][0] , \sa_count[25].r.part0[0] );
tran (\sa_count[25][0] , \sa_count[25].f.lower[0] );
tran (\sa_count[25][1] , \sa_count[25].r.part0[1] );
tran (\sa_count[25][1] , \sa_count[25].f.lower[1] );
tran (\sa_count[25][2] , \sa_count[25].r.part0[2] );
tran (\sa_count[25][2] , \sa_count[25].f.lower[2] );
tran (\sa_count[25][3] , \sa_count[25].r.part0[3] );
tran (\sa_count[25][3] , \sa_count[25].f.lower[3] );
tran (\sa_count[25][4] , \sa_count[25].r.part0[4] );
tran (\sa_count[25][4] , \sa_count[25].f.lower[4] );
tran (\sa_count[25][5] , \sa_count[25].r.part0[5] );
tran (\sa_count[25][5] , \sa_count[25].f.lower[5] );
tran (\sa_count[25][6] , \sa_count[25].r.part0[6] );
tran (\sa_count[25][6] , \sa_count[25].f.lower[6] );
tran (\sa_count[25][7] , \sa_count[25].r.part0[7] );
tran (\sa_count[25][7] , \sa_count[25].f.lower[7] );
tran (\sa_count[25][8] , \sa_count[25].r.part0[8] );
tran (\sa_count[25][8] , \sa_count[25].f.lower[8] );
tran (\sa_count[25][9] , \sa_count[25].r.part0[9] );
tran (\sa_count[25][9] , \sa_count[25].f.lower[9] );
tran (\sa_count[25][10] , \sa_count[25].r.part0[10] );
tran (\sa_count[25][10] , \sa_count[25].f.lower[10] );
tran (\sa_count[25][11] , \sa_count[25].r.part0[11] );
tran (\sa_count[25][11] , \sa_count[25].f.lower[11] );
tran (\sa_count[25][12] , \sa_count[25].r.part0[12] );
tran (\sa_count[25][12] , \sa_count[25].f.lower[12] );
tran (\sa_count[25][13] , \sa_count[25].r.part0[13] );
tran (\sa_count[25][13] , \sa_count[25].f.lower[13] );
tran (\sa_count[25][14] , \sa_count[25].r.part0[14] );
tran (\sa_count[25][14] , \sa_count[25].f.lower[14] );
tran (\sa_count[25][15] , \sa_count[25].r.part0[15] );
tran (\sa_count[25][15] , \sa_count[25].f.lower[15] );
tran (\sa_count[25][16] , \sa_count[25].r.part0[16] );
tran (\sa_count[25][16] , \sa_count[25].f.lower[16] );
tran (\sa_count[25][17] , \sa_count[25].r.part0[17] );
tran (\sa_count[25][17] , \sa_count[25].f.lower[17] );
tran (\sa_count[25][18] , \sa_count[25].r.part0[18] );
tran (\sa_count[25][18] , \sa_count[25].f.lower[18] );
tran (\sa_count[25][19] , \sa_count[25].r.part0[19] );
tran (\sa_count[25][19] , \sa_count[25].f.lower[19] );
tran (\sa_count[25][20] , \sa_count[25].r.part0[20] );
tran (\sa_count[25][20] , \sa_count[25].f.lower[20] );
tran (\sa_count[25][21] , \sa_count[25].r.part0[21] );
tran (\sa_count[25][21] , \sa_count[25].f.lower[21] );
tran (\sa_count[25][22] , \sa_count[25].r.part0[22] );
tran (\sa_count[25][22] , \sa_count[25].f.lower[22] );
tran (\sa_count[25][23] , \sa_count[25].r.part0[23] );
tran (\sa_count[25][23] , \sa_count[25].f.lower[23] );
tran (\sa_count[25][24] , \sa_count[25].r.part0[24] );
tran (\sa_count[25][24] , \sa_count[25].f.lower[24] );
tran (\sa_count[25][25] , \sa_count[25].r.part0[25] );
tran (\sa_count[25][25] , \sa_count[25].f.lower[25] );
tran (\sa_count[25][26] , \sa_count[25].r.part0[26] );
tran (\sa_count[25][26] , \sa_count[25].f.lower[26] );
tran (\sa_count[25][27] , \sa_count[25].r.part0[27] );
tran (\sa_count[25][27] , \sa_count[25].f.lower[27] );
tran (\sa_count[25][28] , \sa_count[25].r.part0[28] );
tran (\sa_count[25][28] , \sa_count[25].f.lower[28] );
tran (\sa_count[25][29] , \sa_count[25].r.part0[29] );
tran (\sa_count[25][29] , \sa_count[25].f.lower[29] );
tran (\sa_count[25][30] , \sa_count[25].r.part0[30] );
tran (\sa_count[25][30] , \sa_count[25].f.lower[30] );
tran (\sa_count[25][31] , \sa_count[25].r.part0[31] );
tran (\sa_count[25][31] , \sa_count[25].f.lower[31] );
tran (\sa_count[25][32] , \sa_count[25].r.part1[0] );
tran (\sa_count[25][32] , \sa_count[25].f.upper[0] );
tran (\sa_count[25][33] , \sa_count[25].r.part1[1] );
tran (\sa_count[25][33] , \sa_count[25].f.upper[1] );
tran (\sa_count[25][34] , \sa_count[25].r.part1[2] );
tran (\sa_count[25][34] , \sa_count[25].f.upper[2] );
tran (\sa_count[25][35] , \sa_count[25].r.part1[3] );
tran (\sa_count[25][35] , \sa_count[25].f.upper[3] );
tran (\sa_count[25][36] , \sa_count[25].r.part1[4] );
tran (\sa_count[25][36] , \sa_count[25].f.upper[4] );
tran (\sa_count[25][37] , \sa_count[25].r.part1[5] );
tran (\sa_count[25][37] , \sa_count[25].f.upper[5] );
tran (\sa_count[25][38] , \sa_count[25].r.part1[6] );
tran (\sa_count[25][38] , \sa_count[25].f.upper[6] );
tran (\sa_count[25][39] , \sa_count[25].r.part1[7] );
tran (\sa_count[25][39] , \sa_count[25].f.upper[7] );
tran (\sa_count[25][40] , \sa_count[25].r.part1[8] );
tran (\sa_count[25][40] , \sa_count[25].f.upper[8] );
tran (\sa_count[25][41] , \sa_count[25].r.part1[9] );
tran (\sa_count[25][41] , \sa_count[25].f.upper[9] );
tran (\sa_count[25][42] , \sa_count[25].r.part1[10] );
tran (\sa_count[25][42] , \sa_count[25].f.upper[10] );
tran (\sa_count[25][43] , \sa_count[25].r.part1[11] );
tran (\sa_count[25][43] , \sa_count[25].f.upper[11] );
tran (\sa_count[25][44] , \sa_count[25].r.part1[12] );
tran (\sa_count[25][44] , \sa_count[25].f.upper[12] );
tran (\sa_count[25][45] , \sa_count[25].r.part1[13] );
tran (\sa_count[25][45] , \sa_count[25].f.upper[13] );
tran (\sa_count[25][46] , \sa_count[25].r.part1[14] );
tran (\sa_count[25][46] , \sa_count[25].f.upper[14] );
tran (\sa_count[25][47] , \sa_count[25].r.part1[15] );
tran (\sa_count[25][47] , \sa_count[25].f.upper[15] );
tran (\sa_count[25][48] , \sa_count[25].r.part1[16] );
tran (\sa_count[25][48] , \sa_count[25].f.upper[16] );
tran (\sa_count[25][49] , \sa_count[25].r.part1[17] );
tran (\sa_count[25][49] , \sa_count[25].f.upper[17] );
tran (\sa_count[25][50] , \sa_count[25].r.part1[18] );
tran (\sa_count[25][50] , \sa_count[25].f.unused[0] );
tran (\sa_count[25][51] , \sa_count[25].r.part1[19] );
tran (\sa_count[25][51] , \sa_count[25].f.unused[1] );
tran (\sa_count[25][52] , \sa_count[25].r.part1[20] );
tran (\sa_count[25][52] , \sa_count[25].f.unused[2] );
tran (\sa_count[25][53] , \sa_count[25].r.part1[21] );
tran (\sa_count[25][53] , \sa_count[25].f.unused[3] );
tran (\sa_count[25][54] , \sa_count[25].r.part1[22] );
tran (\sa_count[25][54] , \sa_count[25].f.unused[4] );
tran (\sa_count[25][55] , \sa_count[25].r.part1[23] );
tran (\sa_count[25][55] , \sa_count[25].f.unused[5] );
tran (\sa_count[25][56] , \sa_count[25].r.part1[24] );
tran (\sa_count[25][56] , \sa_count[25].f.unused[6] );
tran (\sa_count[25][57] , \sa_count[25].r.part1[25] );
tran (\sa_count[25][57] , \sa_count[25].f.unused[7] );
tran (\sa_count[25][58] , \sa_count[25].r.part1[26] );
tran (\sa_count[25][58] , \sa_count[25].f.unused[8] );
tran (\sa_count[25][59] , \sa_count[25].r.part1[27] );
tran (\sa_count[25][59] , \sa_count[25].f.unused[9] );
tran (\sa_count[25][60] , \sa_count[25].r.part1[28] );
tran (\sa_count[25][60] , \sa_count[25].f.unused[10] );
tran (\sa_count[25][61] , \sa_count[25].r.part1[29] );
tran (\sa_count[25][61] , \sa_count[25].f.unused[11] );
tran (\sa_count[25][62] , \sa_count[25].r.part1[30] );
tran (\sa_count[25][62] , \sa_count[25].f.unused[12] );
tran (\sa_count[25][63] , \sa_count[25].r.part1[31] );
tran (\sa_count[25][63] , \sa_count[25].f.unused[13] );
tran (\sa_count[26][0] , \sa_count[26].r.part0[0] );
tran (\sa_count[26][0] , \sa_count[26].f.lower[0] );
tran (\sa_count[26][1] , \sa_count[26].r.part0[1] );
tran (\sa_count[26][1] , \sa_count[26].f.lower[1] );
tran (\sa_count[26][2] , \sa_count[26].r.part0[2] );
tran (\sa_count[26][2] , \sa_count[26].f.lower[2] );
tran (\sa_count[26][3] , \sa_count[26].r.part0[3] );
tran (\sa_count[26][3] , \sa_count[26].f.lower[3] );
tran (\sa_count[26][4] , \sa_count[26].r.part0[4] );
tran (\sa_count[26][4] , \sa_count[26].f.lower[4] );
tran (\sa_count[26][5] , \sa_count[26].r.part0[5] );
tran (\sa_count[26][5] , \sa_count[26].f.lower[5] );
tran (\sa_count[26][6] , \sa_count[26].r.part0[6] );
tran (\sa_count[26][6] , \sa_count[26].f.lower[6] );
tran (\sa_count[26][7] , \sa_count[26].r.part0[7] );
tran (\sa_count[26][7] , \sa_count[26].f.lower[7] );
tran (\sa_count[26][8] , \sa_count[26].r.part0[8] );
tran (\sa_count[26][8] , \sa_count[26].f.lower[8] );
tran (\sa_count[26][9] , \sa_count[26].r.part0[9] );
tran (\sa_count[26][9] , \sa_count[26].f.lower[9] );
tran (\sa_count[26][10] , \sa_count[26].r.part0[10] );
tran (\sa_count[26][10] , \sa_count[26].f.lower[10] );
tran (\sa_count[26][11] , \sa_count[26].r.part0[11] );
tran (\sa_count[26][11] , \sa_count[26].f.lower[11] );
tran (\sa_count[26][12] , \sa_count[26].r.part0[12] );
tran (\sa_count[26][12] , \sa_count[26].f.lower[12] );
tran (\sa_count[26][13] , \sa_count[26].r.part0[13] );
tran (\sa_count[26][13] , \sa_count[26].f.lower[13] );
tran (\sa_count[26][14] , \sa_count[26].r.part0[14] );
tran (\sa_count[26][14] , \sa_count[26].f.lower[14] );
tran (\sa_count[26][15] , \sa_count[26].r.part0[15] );
tran (\sa_count[26][15] , \sa_count[26].f.lower[15] );
tran (\sa_count[26][16] , \sa_count[26].r.part0[16] );
tran (\sa_count[26][16] , \sa_count[26].f.lower[16] );
tran (\sa_count[26][17] , \sa_count[26].r.part0[17] );
tran (\sa_count[26][17] , \sa_count[26].f.lower[17] );
tran (\sa_count[26][18] , \sa_count[26].r.part0[18] );
tran (\sa_count[26][18] , \sa_count[26].f.lower[18] );
tran (\sa_count[26][19] , \sa_count[26].r.part0[19] );
tran (\sa_count[26][19] , \sa_count[26].f.lower[19] );
tran (\sa_count[26][20] , \sa_count[26].r.part0[20] );
tran (\sa_count[26][20] , \sa_count[26].f.lower[20] );
tran (\sa_count[26][21] , \sa_count[26].r.part0[21] );
tran (\sa_count[26][21] , \sa_count[26].f.lower[21] );
tran (\sa_count[26][22] , \sa_count[26].r.part0[22] );
tran (\sa_count[26][22] , \sa_count[26].f.lower[22] );
tran (\sa_count[26][23] , \sa_count[26].r.part0[23] );
tran (\sa_count[26][23] , \sa_count[26].f.lower[23] );
tran (\sa_count[26][24] , \sa_count[26].r.part0[24] );
tran (\sa_count[26][24] , \sa_count[26].f.lower[24] );
tran (\sa_count[26][25] , \sa_count[26].r.part0[25] );
tran (\sa_count[26][25] , \sa_count[26].f.lower[25] );
tran (\sa_count[26][26] , \sa_count[26].r.part0[26] );
tran (\sa_count[26][26] , \sa_count[26].f.lower[26] );
tran (\sa_count[26][27] , \sa_count[26].r.part0[27] );
tran (\sa_count[26][27] , \sa_count[26].f.lower[27] );
tran (\sa_count[26][28] , \sa_count[26].r.part0[28] );
tran (\sa_count[26][28] , \sa_count[26].f.lower[28] );
tran (\sa_count[26][29] , \sa_count[26].r.part0[29] );
tran (\sa_count[26][29] , \sa_count[26].f.lower[29] );
tran (\sa_count[26][30] , \sa_count[26].r.part0[30] );
tran (\sa_count[26][30] , \sa_count[26].f.lower[30] );
tran (\sa_count[26][31] , \sa_count[26].r.part0[31] );
tran (\sa_count[26][31] , \sa_count[26].f.lower[31] );
tran (\sa_count[26][32] , \sa_count[26].r.part1[0] );
tran (\sa_count[26][32] , \sa_count[26].f.upper[0] );
tran (\sa_count[26][33] , \sa_count[26].r.part1[1] );
tran (\sa_count[26][33] , \sa_count[26].f.upper[1] );
tran (\sa_count[26][34] , \sa_count[26].r.part1[2] );
tran (\sa_count[26][34] , \sa_count[26].f.upper[2] );
tran (\sa_count[26][35] , \sa_count[26].r.part1[3] );
tran (\sa_count[26][35] , \sa_count[26].f.upper[3] );
tran (\sa_count[26][36] , \sa_count[26].r.part1[4] );
tran (\sa_count[26][36] , \sa_count[26].f.upper[4] );
tran (\sa_count[26][37] , \sa_count[26].r.part1[5] );
tran (\sa_count[26][37] , \sa_count[26].f.upper[5] );
tran (\sa_count[26][38] , \sa_count[26].r.part1[6] );
tran (\sa_count[26][38] , \sa_count[26].f.upper[6] );
tran (\sa_count[26][39] , \sa_count[26].r.part1[7] );
tran (\sa_count[26][39] , \sa_count[26].f.upper[7] );
tran (\sa_count[26][40] , \sa_count[26].r.part1[8] );
tran (\sa_count[26][40] , \sa_count[26].f.upper[8] );
tran (\sa_count[26][41] , \sa_count[26].r.part1[9] );
tran (\sa_count[26][41] , \sa_count[26].f.upper[9] );
tran (\sa_count[26][42] , \sa_count[26].r.part1[10] );
tran (\sa_count[26][42] , \sa_count[26].f.upper[10] );
tran (\sa_count[26][43] , \sa_count[26].r.part1[11] );
tran (\sa_count[26][43] , \sa_count[26].f.upper[11] );
tran (\sa_count[26][44] , \sa_count[26].r.part1[12] );
tran (\sa_count[26][44] , \sa_count[26].f.upper[12] );
tran (\sa_count[26][45] , \sa_count[26].r.part1[13] );
tran (\sa_count[26][45] , \sa_count[26].f.upper[13] );
tran (\sa_count[26][46] , \sa_count[26].r.part1[14] );
tran (\sa_count[26][46] , \sa_count[26].f.upper[14] );
tran (\sa_count[26][47] , \sa_count[26].r.part1[15] );
tran (\sa_count[26][47] , \sa_count[26].f.upper[15] );
tran (\sa_count[26][48] , \sa_count[26].r.part1[16] );
tran (\sa_count[26][48] , \sa_count[26].f.upper[16] );
tran (\sa_count[26][49] , \sa_count[26].r.part1[17] );
tran (\sa_count[26][49] , \sa_count[26].f.upper[17] );
tran (\sa_count[26][50] , \sa_count[26].r.part1[18] );
tran (\sa_count[26][50] , \sa_count[26].f.unused[0] );
tran (\sa_count[26][51] , \sa_count[26].r.part1[19] );
tran (\sa_count[26][51] , \sa_count[26].f.unused[1] );
tran (\sa_count[26][52] , \sa_count[26].r.part1[20] );
tran (\sa_count[26][52] , \sa_count[26].f.unused[2] );
tran (\sa_count[26][53] , \sa_count[26].r.part1[21] );
tran (\sa_count[26][53] , \sa_count[26].f.unused[3] );
tran (\sa_count[26][54] , \sa_count[26].r.part1[22] );
tran (\sa_count[26][54] , \sa_count[26].f.unused[4] );
tran (\sa_count[26][55] , \sa_count[26].r.part1[23] );
tran (\sa_count[26][55] , \sa_count[26].f.unused[5] );
tran (\sa_count[26][56] , \sa_count[26].r.part1[24] );
tran (\sa_count[26][56] , \sa_count[26].f.unused[6] );
tran (\sa_count[26][57] , \sa_count[26].r.part1[25] );
tran (\sa_count[26][57] , \sa_count[26].f.unused[7] );
tran (\sa_count[26][58] , \sa_count[26].r.part1[26] );
tran (\sa_count[26][58] , \sa_count[26].f.unused[8] );
tran (\sa_count[26][59] , \sa_count[26].r.part1[27] );
tran (\sa_count[26][59] , \sa_count[26].f.unused[9] );
tran (\sa_count[26][60] , \sa_count[26].r.part1[28] );
tran (\sa_count[26][60] , \sa_count[26].f.unused[10] );
tran (\sa_count[26][61] , \sa_count[26].r.part1[29] );
tran (\sa_count[26][61] , \sa_count[26].f.unused[11] );
tran (\sa_count[26][62] , \sa_count[26].r.part1[30] );
tran (\sa_count[26][62] , \sa_count[26].f.unused[12] );
tran (\sa_count[26][63] , \sa_count[26].r.part1[31] );
tran (\sa_count[26][63] , \sa_count[26].f.unused[13] );
tran (\sa_count[27][0] , \sa_count[27].r.part0[0] );
tran (\sa_count[27][0] , \sa_count[27].f.lower[0] );
tran (\sa_count[27][1] , \sa_count[27].r.part0[1] );
tran (\sa_count[27][1] , \sa_count[27].f.lower[1] );
tran (\sa_count[27][2] , \sa_count[27].r.part0[2] );
tran (\sa_count[27][2] , \sa_count[27].f.lower[2] );
tran (\sa_count[27][3] , \sa_count[27].r.part0[3] );
tran (\sa_count[27][3] , \sa_count[27].f.lower[3] );
tran (\sa_count[27][4] , \sa_count[27].r.part0[4] );
tran (\sa_count[27][4] , \sa_count[27].f.lower[4] );
tran (\sa_count[27][5] , \sa_count[27].r.part0[5] );
tran (\sa_count[27][5] , \sa_count[27].f.lower[5] );
tran (\sa_count[27][6] , \sa_count[27].r.part0[6] );
tran (\sa_count[27][6] , \sa_count[27].f.lower[6] );
tran (\sa_count[27][7] , \sa_count[27].r.part0[7] );
tran (\sa_count[27][7] , \sa_count[27].f.lower[7] );
tran (\sa_count[27][8] , \sa_count[27].r.part0[8] );
tran (\sa_count[27][8] , \sa_count[27].f.lower[8] );
tran (\sa_count[27][9] , \sa_count[27].r.part0[9] );
tran (\sa_count[27][9] , \sa_count[27].f.lower[9] );
tran (\sa_count[27][10] , \sa_count[27].r.part0[10] );
tran (\sa_count[27][10] , \sa_count[27].f.lower[10] );
tran (\sa_count[27][11] , \sa_count[27].r.part0[11] );
tran (\sa_count[27][11] , \sa_count[27].f.lower[11] );
tran (\sa_count[27][12] , \sa_count[27].r.part0[12] );
tran (\sa_count[27][12] , \sa_count[27].f.lower[12] );
tran (\sa_count[27][13] , \sa_count[27].r.part0[13] );
tran (\sa_count[27][13] , \sa_count[27].f.lower[13] );
tran (\sa_count[27][14] , \sa_count[27].r.part0[14] );
tran (\sa_count[27][14] , \sa_count[27].f.lower[14] );
tran (\sa_count[27][15] , \sa_count[27].r.part0[15] );
tran (\sa_count[27][15] , \sa_count[27].f.lower[15] );
tran (\sa_count[27][16] , \sa_count[27].r.part0[16] );
tran (\sa_count[27][16] , \sa_count[27].f.lower[16] );
tran (\sa_count[27][17] , \sa_count[27].r.part0[17] );
tran (\sa_count[27][17] , \sa_count[27].f.lower[17] );
tran (\sa_count[27][18] , \sa_count[27].r.part0[18] );
tran (\sa_count[27][18] , \sa_count[27].f.lower[18] );
tran (\sa_count[27][19] , \sa_count[27].r.part0[19] );
tran (\sa_count[27][19] , \sa_count[27].f.lower[19] );
tran (\sa_count[27][20] , \sa_count[27].r.part0[20] );
tran (\sa_count[27][20] , \sa_count[27].f.lower[20] );
tran (\sa_count[27][21] , \sa_count[27].r.part0[21] );
tran (\sa_count[27][21] , \sa_count[27].f.lower[21] );
tran (\sa_count[27][22] , \sa_count[27].r.part0[22] );
tran (\sa_count[27][22] , \sa_count[27].f.lower[22] );
tran (\sa_count[27][23] , \sa_count[27].r.part0[23] );
tran (\sa_count[27][23] , \sa_count[27].f.lower[23] );
tran (\sa_count[27][24] , \sa_count[27].r.part0[24] );
tran (\sa_count[27][24] , \sa_count[27].f.lower[24] );
tran (\sa_count[27][25] , \sa_count[27].r.part0[25] );
tran (\sa_count[27][25] , \sa_count[27].f.lower[25] );
tran (\sa_count[27][26] , \sa_count[27].r.part0[26] );
tran (\sa_count[27][26] , \sa_count[27].f.lower[26] );
tran (\sa_count[27][27] , \sa_count[27].r.part0[27] );
tran (\sa_count[27][27] , \sa_count[27].f.lower[27] );
tran (\sa_count[27][28] , \sa_count[27].r.part0[28] );
tran (\sa_count[27][28] , \sa_count[27].f.lower[28] );
tran (\sa_count[27][29] , \sa_count[27].r.part0[29] );
tran (\sa_count[27][29] , \sa_count[27].f.lower[29] );
tran (\sa_count[27][30] , \sa_count[27].r.part0[30] );
tran (\sa_count[27][30] , \sa_count[27].f.lower[30] );
tran (\sa_count[27][31] , \sa_count[27].r.part0[31] );
tran (\sa_count[27][31] , \sa_count[27].f.lower[31] );
tran (\sa_count[27][32] , \sa_count[27].r.part1[0] );
tran (\sa_count[27][32] , \sa_count[27].f.upper[0] );
tran (\sa_count[27][33] , \sa_count[27].r.part1[1] );
tran (\sa_count[27][33] , \sa_count[27].f.upper[1] );
tran (\sa_count[27][34] , \sa_count[27].r.part1[2] );
tran (\sa_count[27][34] , \sa_count[27].f.upper[2] );
tran (\sa_count[27][35] , \sa_count[27].r.part1[3] );
tran (\sa_count[27][35] , \sa_count[27].f.upper[3] );
tran (\sa_count[27][36] , \sa_count[27].r.part1[4] );
tran (\sa_count[27][36] , \sa_count[27].f.upper[4] );
tran (\sa_count[27][37] , \sa_count[27].r.part1[5] );
tran (\sa_count[27][37] , \sa_count[27].f.upper[5] );
tran (\sa_count[27][38] , \sa_count[27].r.part1[6] );
tran (\sa_count[27][38] , \sa_count[27].f.upper[6] );
tran (\sa_count[27][39] , \sa_count[27].r.part1[7] );
tran (\sa_count[27][39] , \sa_count[27].f.upper[7] );
tran (\sa_count[27][40] , \sa_count[27].r.part1[8] );
tran (\sa_count[27][40] , \sa_count[27].f.upper[8] );
tran (\sa_count[27][41] , \sa_count[27].r.part1[9] );
tran (\sa_count[27][41] , \sa_count[27].f.upper[9] );
tran (\sa_count[27][42] , \sa_count[27].r.part1[10] );
tran (\sa_count[27][42] , \sa_count[27].f.upper[10] );
tran (\sa_count[27][43] , \sa_count[27].r.part1[11] );
tran (\sa_count[27][43] , \sa_count[27].f.upper[11] );
tran (\sa_count[27][44] , \sa_count[27].r.part1[12] );
tran (\sa_count[27][44] , \sa_count[27].f.upper[12] );
tran (\sa_count[27][45] , \sa_count[27].r.part1[13] );
tran (\sa_count[27][45] , \sa_count[27].f.upper[13] );
tran (\sa_count[27][46] , \sa_count[27].r.part1[14] );
tran (\sa_count[27][46] , \sa_count[27].f.upper[14] );
tran (\sa_count[27][47] , \sa_count[27].r.part1[15] );
tran (\sa_count[27][47] , \sa_count[27].f.upper[15] );
tran (\sa_count[27][48] , \sa_count[27].r.part1[16] );
tran (\sa_count[27][48] , \sa_count[27].f.upper[16] );
tran (\sa_count[27][49] , \sa_count[27].r.part1[17] );
tran (\sa_count[27][49] , \sa_count[27].f.upper[17] );
tran (\sa_count[27][50] , \sa_count[27].r.part1[18] );
tran (\sa_count[27][50] , \sa_count[27].f.unused[0] );
tran (\sa_count[27][51] , \sa_count[27].r.part1[19] );
tran (\sa_count[27][51] , \sa_count[27].f.unused[1] );
tran (\sa_count[27][52] , \sa_count[27].r.part1[20] );
tran (\sa_count[27][52] , \sa_count[27].f.unused[2] );
tran (\sa_count[27][53] , \sa_count[27].r.part1[21] );
tran (\sa_count[27][53] , \sa_count[27].f.unused[3] );
tran (\sa_count[27][54] , \sa_count[27].r.part1[22] );
tran (\sa_count[27][54] , \sa_count[27].f.unused[4] );
tran (\sa_count[27][55] , \sa_count[27].r.part1[23] );
tran (\sa_count[27][55] , \sa_count[27].f.unused[5] );
tran (\sa_count[27][56] , \sa_count[27].r.part1[24] );
tran (\sa_count[27][56] , \sa_count[27].f.unused[6] );
tran (\sa_count[27][57] , \sa_count[27].r.part1[25] );
tran (\sa_count[27][57] , \sa_count[27].f.unused[7] );
tran (\sa_count[27][58] , \sa_count[27].r.part1[26] );
tran (\sa_count[27][58] , \sa_count[27].f.unused[8] );
tran (\sa_count[27][59] , \sa_count[27].r.part1[27] );
tran (\sa_count[27][59] , \sa_count[27].f.unused[9] );
tran (\sa_count[27][60] , \sa_count[27].r.part1[28] );
tran (\sa_count[27][60] , \sa_count[27].f.unused[10] );
tran (\sa_count[27][61] , \sa_count[27].r.part1[29] );
tran (\sa_count[27][61] , \sa_count[27].f.unused[11] );
tran (\sa_count[27][62] , \sa_count[27].r.part1[30] );
tran (\sa_count[27][62] , \sa_count[27].f.unused[12] );
tran (\sa_count[27][63] , \sa_count[27].r.part1[31] );
tran (\sa_count[27][63] , \sa_count[27].f.unused[13] );
tran (\sa_count[28][0] , \sa_count[28].r.part0[0] );
tran (\sa_count[28][0] , \sa_count[28].f.lower[0] );
tran (\sa_count[28][1] , \sa_count[28].r.part0[1] );
tran (\sa_count[28][1] , \sa_count[28].f.lower[1] );
tran (\sa_count[28][2] , \sa_count[28].r.part0[2] );
tran (\sa_count[28][2] , \sa_count[28].f.lower[2] );
tran (\sa_count[28][3] , \sa_count[28].r.part0[3] );
tran (\sa_count[28][3] , \sa_count[28].f.lower[3] );
tran (\sa_count[28][4] , \sa_count[28].r.part0[4] );
tran (\sa_count[28][4] , \sa_count[28].f.lower[4] );
tran (\sa_count[28][5] , \sa_count[28].r.part0[5] );
tran (\sa_count[28][5] , \sa_count[28].f.lower[5] );
tran (\sa_count[28][6] , \sa_count[28].r.part0[6] );
tran (\sa_count[28][6] , \sa_count[28].f.lower[6] );
tran (\sa_count[28][7] , \sa_count[28].r.part0[7] );
tran (\sa_count[28][7] , \sa_count[28].f.lower[7] );
tran (\sa_count[28][8] , \sa_count[28].r.part0[8] );
tran (\sa_count[28][8] , \sa_count[28].f.lower[8] );
tran (\sa_count[28][9] , \sa_count[28].r.part0[9] );
tran (\sa_count[28][9] , \sa_count[28].f.lower[9] );
tran (\sa_count[28][10] , \sa_count[28].r.part0[10] );
tran (\sa_count[28][10] , \sa_count[28].f.lower[10] );
tran (\sa_count[28][11] , \sa_count[28].r.part0[11] );
tran (\sa_count[28][11] , \sa_count[28].f.lower[11] );
tran (\sa_count[28][12] , \sa_count[28].r.part0[12] );
tran (\sa_count[28][12] , \sa_count[28].f.lower[12] );
tran (\sa_count[28][13] , \sa_count[28].r.part0[13] );
tran (\sa_count[28][13] , \sa_count[28].f.lower[13] );
tran (\sa_count[28][14] , \sa_count[28].r.part0[14] );
tran (\sa_count[28][14] , \sa_count[28].f.lower[14] );
tran (\sa_count[28][15] , \sa_count[28].r.part0[15] );
tran (\sa_count[28][15] , \sa_count[28].f.lower[15] );
tran (\sa_count[28][16] , \sa_count[28].r.part0[16] );
tran (\sa_count[28][16] , \sa_count[28].f.lower[16] );
tran (\sa_count[28][17] , \sa_count[28].r.part0[17] );
tran (\sa_count[28][17] , \sa_count[28].f.lower[17] );
tran (\sa_count[28][18] , \sa_count[28].r.part0[18] );
tran (\sa_count[28][18] , \sa_count[28].f.lower[18] );
tran (\sa_count[28][19] , \sa_count[28].r.part0[19] );
tran (\sa_count[28][19] , \sa_count[28].f.lower[19] );
tran (\sa_count[28][20] , \sa_count[28].r.part0[20] );
tran (\sa_count[28][20] , \sa_count[28].f.lower[20] );
tran (\sa_count[28][21] , \sa_count[28].r.part0[21] );
tran (\sa_count[28][21] , \sa_count[28].f.lower[21] );
tran (\sa_count[28][22] , \sa_count[28].r.part0[22] );
tran (\sa_count[28][22] , \sa_count[28].f.lower[22] );
tran (\sa_count[28][23] , \sa_count[28].r.part0[23] );
tran (\sa_count[28][23] , \sa_count[28].f.lower[23] );
tran (\sa_count[28][24] , \sa_count[28].r.part0[24] );
tran (\sa_count[28][24] , \sa_count[28].f.lower[24] );
tran (\sa_count[28][25] , \sa_count[28].r.part0[25] );
tran (\sa_count[28][25] , \sa_count[28].f.lower[25] );
tran (\sa_count[28][26] , \sa_count[28].r.part0[26] );
tran (\sa_count[28][26] , \sa_count[28].f.lower[26] );
tran (\sa_count[28][27] , \sa_count[28].r.part0[27] );
tran (\sa_count[28][27] , \sa_count[28].f.lower[27] );
tran (\sa_count[28][28] , \sa_count[28].r.part0[28] );
tran (\sa_count[28][28] , \sa_count[28].f.lower[28] );
tran (\sa_count[28][29] , \sa_count[28].r.part0[29] );
tran (\sa_count[28][29] , \sa_count[28].f.lower[29] );
tran (\sa_count[28][30] , \sa_count[28].r.part0[30] );
tran (\sa_count[28][30] , \sa_count[28].f.lower[30] );
tran (\sa_count[28][31] , \sa_count[28].r.part0[31] );
tran (\sa_count[28][31] , \sa_count[28].f.lower[31] );
tran (\sa_count[28][32] , \sa_count[28].r.part1[0] );
tran (\sa_count[28][32] , \sa_count[28].f.upper[0] );
tran (\sa_count[28][33] , \sa_count[28].r.part1[1] );
tran (\sa_count[28][33] , \sa_count[28].f.upper[1] );
tran (\sa_count[28][34] , \sa_count[28].r.part1[2] );
tran (\sa_count[28][34] , \sa_count[28].f.upper[2] );
tran (\sa_count[28][35] , \sa_count[28].r.part1[3] );
tran (\sa_count[28][35] , \sa_count[28].f.upper[3] );
tran (\sa_count[28][36] , \sa_count[28].r.part1[4] );
tran (\sa_count[28][36] , \sa_count[28].f.upper[4] );
tran (\sa_count[28][37] , \sa_count[28].r.part1[5] );
tran (\sa_count[28][37] , \sa_count[28].f.upper[5] );
tran (\sa_count[28][38] , \sa_count[28].r.part1[6] );
tran (\sa_count[28][38] , \sa_count[28].f.upper[6] );
tran (\sa_count[28][39] , \sa_count[28].r.part1[7] );
tran (\sa_count[28][39] , \sa_count[28].f.upper[7] );
tran (\sa_count[28][40] , \sa_count[28].r.part1[8] );
tran (\sa_count[28][40] , \sa_count[28].f.upper[8] );
tran (\sa_count[28][41] , \sa_count[28].r.part1[9] );
tran (\sa_count[28][41] , \sa_count[28].f.upper[9] );
tran (\sa_count[28][42] , \sa_count[28].r.part1[10] );
tran (\sa_count[28][42] , \sa_count[28].f.upper[10] );
tran (\sa_count[28][43] , \sa_count[28].r.part1[11] );
tran (\sa_count[28][43] , \sa_count[28].f.upper[11] );
tran (\sa_count[28][44] , \sa_count[28].r.part1[12] );
tran (\sa_count[28][44] , \sa_count[28].f.upper[12] );
tran (\sa_count[28][45] , \sa_count[28].r.part1[13] );
tran (\sa_count[28][45] , \sa_count[28].f.upper[13] );
tran (\sa_count[28][46] , \sa_count[28].r.part1[14] );
tran (\sa_count[28][46] , \sa_count[28].f.upper[14] );
tran (\sa_count[28][47] , \sa_count[28].r.part1[15] );
tran (\sa_count[28][47] , \sa_count[28].f.upper[15] );
tran (\sa_count[28][48] , \sa_count[28].r.part1[16] );
tran (\sa_count[28][48] , \sa_count[28].f.upper[16] );
tran (\sa_count[28][49] , \sa_count[28].r.part1[17] );
tran (\sa_count[28][49] , \sa_count[28].f.upper[17] );
tran (\sa_count[28][50] , \sa_count[28].r.part1[18] );
tran (\sa_count[28][50] , \sa_count[28].f.unused[0] );
tran (\sa_count[28][51] , \sa_count[28].r.part1[19] );
tran (\sa_count[28][51] , \sa_count[28].f.unused[1] );
tran (\sa_count[28][52] , \sa_count[28].r.part1[20] );
tran (\sa_count[28][52] , \sa_count[28].f.unused[2] );
tran (\sa_count[28][53] , \sa_count[28].r.part1[21] );
tran (\sa_count[28][53] , \sa_count[28].f.unused[3] );
tran (\sa_count[28][54] , \sa_count[28].r.part1[22] );
tran (\sa_count[28][54] , \sa_count[28].f.unused[4] );
tran (\sa_count[28][55] , \sa_count[28].r.part1[23] );
tran (\sa_count[28][55] , \sa_count[28].f.unused[5] );
tran (\sa_count[28][56] , \sa_count[28].r.part1[24] );
tran (\sa_count[28][56] , \sa_count[28].f.unused[6] );
tran (\sa_count[28][57] , \sa_count[28].r.part1[25] );
tran (\sa_count[28][57] , \sa_count[28].f.unused[7] );
tran (\sa_count[28][58] , \sa_count[28].r.part1[26] );
tran (\sa_count[28][58] , \sa_count[28].f.unused[8] );
tran (\sa_count[28][59] , \sa_count[28].r.part1[27] );
tran (\sa_count[28][59] , \sa_count[28].f.unused[9] );
tran (\sa_count[28][60] , \sa_count[28].r.part1[28] );
tran (\sa_count[28][60] , \sa_count[28].f.unused[10] );
tran (\sa_count[28][61] , \sa_count[28].r.part1[29] );
tran (\sa_count[28][61] , \sa_count[28].f.unused[11] );
tran (\sa_count[28][62] , \sa_count[28].r.part1[30] );
tran (\sa_count[28][62] , \sa_count[28].f.unused[12] );
tran (\sa_count[28][63] , \sa_count[28].r.part1[31] );
tran (\sa_count[28][63] , \sa_count[28].f.unused[13] );
tran (\sa_count[29][0] , \sa_count[29].r.part0[0] );
tran (\sa_count[29][0] , \sa_count[29].f.lower[0] );
tran (\sa_count[29][1] , \sa_count[29].r.part0[1] );
tran (\sa_count[29][1] , \sa_count[29].f.lower[1] );
tran (\sa_count[29][2] , \sa_count[29].r.part0[2] );
tran (\sa_count[29][2] , \sa_count[29].f.lower[2] );
tran (\sa_count[29][3] , \sa_count[29].r.part0[3] );
tran (\sa_count[29][3] , \sa_count[29].f.lower[3] );
tran (\sa_count[29][4] , \sa_count[29].r.part0[4] );
tran (\sa_count[29][4] , \sa_count[29].f.lower[4] );
tran (\sa_count[29][5] , \sa_count[29].r.part0[5] );
tran (\sa_count[29][5] , \sa_count[29].f.lower[5] );
tran (\sa_count[29][6] , \sa_count[29].r.part0[6] );
tran (\sa_count[29][6] , \sa_count[29].f.lower[6] );
tran (\sa_count[29][7] , \sa_count[29].r.part0[7] );
tran (\sa_count[29][7] , \sa_count[29].f.lower[7] );
tran (\sa_count[29][8] , \sa_count[29].r.part0[8] );
tran (\sa_count[29][8] , \sa_count[29].f.lower[8] );
tran (\sa_count[29][9] , \sa_count[29].r.part0[9] );
tran (\sa_count[29][9] , \sa_count[29].f.lower[9] );
tran (\sa_count[29][10] , \sa_count[29].r.part0[10] );
tran (\sa_count[29][10] , \sa_count[29].f.lower[10] );
tran (\sa_count[29][11] , \sa_count[29].r.part0[11] );
tran (\sa_count[29][11] , \sa_count[29].f.lower[11] );
tran (\sa_count[29][12] , \sa_count[29].r.part0[12] );
tran (\sa_count[29][12] , \sa_count[29].f.lower[12] );
tran (\sa_count[29][13] , \sa_count[29].r.part0[13] );
tran (\sa_count[29][13] , \sa_count[29].f.lower[13] );
tran (\sa_count[29][14] , \sa_count[29].r.part0[14] );
tran (\sa_count[29][14] , \sa_count[29].f.lower[14] );
tran (\sa_count[29][15] , \sa_count[29].r.part0[15] );
tran (\sa_count[29][15] , \sa_count[29].f.lower[15] );
tran (\sa_count[29][16] , \sa_count[29].r.part0[16] );
tran (\sa_count[29][16] , \sa_count[29].f.lower[16] );
tran (\sa_count[29][17] , \sa_count[29].r.part0[17] );
tran (\sa_count[29][17] , \sa_count[29].f.lower[17] );
tran (\sa_count[29][18] , \sa_count[29].r.part0[18] );
tran (\sa_count[29][18] , \sa_count[29].f.lower[18] );
tran (\sa_count[29][19] , \sa_count[29].r.part0[19] );
tran (\sa_count[29][19] , \sa_count[29].f.lower[19] );
tran (\sa_count[29][20] , \sa_count[29].r.part0[20] );
tran (\sa_count[29][20] , \sa_count[29].f.lower[20] );
tran (\sa_count[29][21] , \sa_count[29].r.part0[21] );
tran (\sa_count[29][21] , \sa_count[29].f.lower[21] );
tran (\sa_count[29][22] , \sa_count[29].r.part0[22] );
tran (\sa_count[29][22] , \sa_count[29].f.lower[22] );
tran (\sa_count[29][23] , \sa_count[29].r.part0[23] );
tran (\sa_count[29][23] , \sa_count[29].f.lower[23] );
tran (\sa_count[29][24] , \sa_count[29].r.part0[24] );
tran (\sa_count[29][24] , \sa_count[29].f.lower[24] );
tran (\sa_count[29][25] , \sa_count[29].r.part0[25] );
tran (\sa_count[29][25] , \sa_count[29].f.lower[25] );
tran (\sa_count[29][26] , \sa_count[29].r.part0[26] );
tran (\sa_count[29][26] , \sa_count[29].f.lower[26] );
tran (\sa_count[29][27] , \sa_count[29].r.part0[27] );
tran (\sa_count[29][27] , \sa_count[29].f.lower[27] );
tran (\sa_count[29][28] , \sa_count[29].r.part0[28] );
tran (\sa_count[29][28] , \sa_count[29].f.lower[28] );
tran (\sa_count[29][29] , \sa_count[29].r.part0[29] );
tran (\sa_count[29][29] , \sa_count[29].f.lower[29] );
tran (\sa_count[29][30] , \sa_count[29].r.part0[30] );
tran (\sa_count[29][30] , \sa_count[29].f.lower[30] );
tran (\sa_count[29][31] , \sa_count[29].r.part0[31] );
tran (\sa_count[29][31] , \sa_count[29].f.lower[31] );
tran (\sa_count[29][32] , \sa_count[29].r.part1[0] );
tran (\sa_count[29][32] , \sa_count[29].f.upper[0] );
tran (\sa_count[29][33] , \sa_count[29].r.part1[1] );
tran (\sa_count[29][33] , \sa_count[29].f.upper[1] );
tran (\sa_count[29][34] , \sa_count[29].r.part1[2] );
tran (\sa_count[29][34] , \sa_count[29].f.upper[2] );
tran (\sa_count[29][35] , \sa_count[29].r.part1[3] );
tran (\sa_count[29][35] , \sa_count[29].f.upper[3] );
tran (\sa_count[29][36] , \sa_count[29].r.part1[4] );
tran (\sa_count[29][36] , \sa_count[29].f.upper[4] );
tran (\sa_count[29][37] , \sa_count[29].r.part1[5] );
tran (\sa_count[29][37] , \sa_count[29].f.upper[5] );
tran (\sa_count[29][38] , \sa_count[29].r.part1[6] );
tran (\sa_count[29][38] , \sa_count[29].f.upper[6] );
tran (\sa_count[29][39] , \sa_count[29].r.part1[7] );
tran (\sa_count[29][39] , \sa_count[29].f.upper[7] );
tran (\sa_count[29][40] , \sa_count[29].r.part1[8] );
tran (\sa_count[29][40] , \sa_count[29].f.upper[8] );
tran (\sa_count[29][41] , \sa_count[29].r.part1[9] );
tran (\sa_count[29][41] , \sa_count[29].f.upper[9] );
tran (\sa_count[29][42] , \sa_count[29].r.part1[10] );
tran (\sa_count[29][42] , \sa_count[29].f.upper[10] );
tran (\sa_count[29][43] , \sa_count[29].r.part1[11] );
tran (\sa_count[29][43] , \sa_count[29].f.upper[11] );
tran (\sa_count[29][44] , \sa_count[29].r.part1[12] );
tran (\sa_count[29][44] , \sa_count[29].f.upper[12] );
tran (\sa_count[29][45] , \sa_count[29].r.part1[13] );
tran (\sa_count[29][45] , \sa_count[29].f.upper[13] );
tran (\sa_count[29][46] , \sa_count[29].r.part1[14] );
tran (\sa_count[29][46] , \sa_count[29].f.upper[14] );
tran (\sa_count[29][47] , \sa_count[29].r.part1[15] );
tran (\sa_count[29][47] , \sa_count[29].f.upper[15] );
tran (\sa_count[29][48] , \sa_count[29].r.part1[16] );
tran (\sa_count[29][48] , \sa_count[29].f.upper[16] );
tran (\sa_count[29][49] , \sa_count[29].r.part1[17] );
tran (\sa_count[29][49] , \sa_count[29].f.upper[17] );
tran (\sa_count[29][50] , \sa_count[29].r.part1[18] );
tran (\sa_count[29][50] , \sa_count[29].f.unused[0] );
tran (\sa_count[29][51] , \sa_count[29].r.part1[19] );
tran (\sa_count[29][51] , \sa_count[29].f.unused[1] );
tran (\sa_count[29][52] , \sa_count[29].r.part1[20] );
tran (\sa_count[29][52] , \sa_count[29].f.unused[2] );
tran (\sa_count[29][53] , \sa_count[29].r.part1[21] );
tran (\sa_count[29][53] , \sa_count[29].f.unused[3] );
tran (\sa_count[29][54] , \sa_count[29].r.part1[22] );
tran (\sa_count[29][54] , \sa_count[29].f.unused[4] );
tran (\sa_count[29][55] , \sa_count[29].r.part1[23] );
tran (\sa_count[29][55] , \sa_count[29].f.unused[5] );
tran (\sa_count[29][56] , \sa_count[29].r.part1[24] );
tran (\sa_count[29][56] , \sa_count[29].f.unused[6] );
tran (\sa_count[29][57] , \sa_count[29].r.part1[25] );
tran (\sa_count[29][57] , \sa_count[29].f.unused[7] );
tran (\sa_count[29][58] , \sa_count[29].r.part1[26] );
tran (\sa_count[29][58] , \sa_count[29].f.unused[8] );
tran (\sa_count[29][59] , \sa_count[29].r.part1[27] );
tran (\sa_count[29][59] , \sa_count[29].f.unused[9] );
tran (\sa_count[29][60] , \sa_count[29].r.part1[28] );
tran (\sa_count[29][60] , \sa_count[29].f.unused[10] );
tran (\sa_count[29][61] , \sa_count[29].r.part1[29] );
tran (\sa_count[29][61] , \sa_count[29].f.unused[11] );
tran (\sa_count[29][62] , \sa_count[29].r.part1[30] );
tran (\sa_count[29][62] , \sa_count[29].f.unused[12] );
tran (\sa_count[29][63] , \sa_count[29].r.part1[31] );
tran (\sa_count[29][63] , \sa_count[29].f.unused[13] );
tran (\sa_count[30][0] , \sa_count[30].r.part0[0] );
tran (\sa_count[30][0] , \sa_count[30].f.lower[0] );
tran (\sa_count[30][1] , \sa_count[30].r.part0[1] );
tran (\sa_count[30][1] , \sa_count[30].f.lower[1] );
tran (\sa_count[30][2] , \sa_count[30].r.part0[2] );
tran (\sa_count[30][2] , \sa_count[30].f.lower[2] );
tran (\sa_count[30][3] , \sa_count[30].r.part0[3] );
tran (\sa_count[30][3] , \sa_count[30].f.lower[3] );
tran (\sa_count[30][4] , \sa_count[30].r.part0[4] );
tran (\sa_count[30][4] , \sa_count[30].f.lower[4] );
tran (\sa_count[30][5] , \sa_count[30].r.part0[5] );
tran (\sa_count[30][5] , \sa_count[30].f.lower[5] );
tran (\sa_count[30][6] , \sa_count[30].r.part0[6] );
tran (\sa_count[30][6] , \sa_count[30].f.lower[6] );
tran (\sa_count[30][7] , \sa_count[30].r.part0[7] );
tran (\sa_count[30][7] , \sa_count[30].f.lower[7] );
tran (\sa_count[30][8] , \sa_count[30].r.part0[8] );
tran (\sa_count[30][8] , \sa_count[30].f.lower[8] );
tran (\sa_count[30][9] , \sa_count[30].r.part0[9] );
tran (\sa_count[30][9] , \sa_count[30].f.lower[9] );
tran (\sa_count[30][10] , \sa_count[30].r.part0[10] );
tran (\sa_count[30][10] , \sa_count[30].f.lower[10] );
tran (\sa_count[30][11] , \sa_count[30].r.part0[11] );
tran (\sa_count[30][11] , \sa_count[30].f.lower[11] );
tran (\sa_count[30][12] , \sa_count[30].r.part0[12] );
tran (\sa_count[30][12] , \sa_count[30].f.lower[12] );
tran (\sa_count[30][13] , \sa_count[30].r.part0[13] );
tran (\sa_count[30][13] , \sa_count[30].f.lower[13] );
tran (\sa_count[30][14] , \sa_count[30].r.part0[14] );
tran (\sa_count[30][14] , \sa_count[30].f.lower[14] );
tran (\sa_count[30][15] , \sa_count[30].r.part0[15] );
tran (\sa_count[30][15] , \sa_count[30].f.lower[15] );
tran (\sa_count[30][16] , \sa_count[30].r.part0[16] );
tran (\sa_count[30][16] , \sa_count[30].f.lower[16] );
tran (\sa_count[30][17] , \sa_count[30].r.part0[17] );
tran (\sa_count[30][17] , \sa_count[30].f.lower[17] );
tran (\sa_count[30][18] , \sa_count[30].r.part0[18] );
tran (\sa_count[30][18] , \sa_count[30].f.lower[18] );
tran (\sa_count[30][19] , \sa_count[30].r.part0[19] );
tran (\sa_count[30][19] , \sa_count[30].f.lower[19] );
tran (\sa_count[30][20] , \sa_count[30].r.part0[20] );
tran (\sa_count[30][20] , \sa_count[30].f.lower[20] );
tran (\sa_count[30][21] , \sa_count[30].r.part0[21] );
tran (\sa_count[30][21] , \sa_count[30].f.lower[21] );
tran (\sa_count[30][22] , \sa_count[30].r.part0[22] );
tran (\sa_count[30][22] , \sa_count[30].f.lower[22] );
tran (\sa_count[30][23] , \sa_count[30].r.part0[23] );
tran (\sa_count[30][23] , \sa_count[30].f.lower[23] );
tran (\sa_count[30][24] , \sa_count[30].r.part0[24] );
tran (\sa_count[30][24] , \sa_count[30].f.lower[24] );
tran (\sa_count[30][25] , \sa_count[30].r.part0[25] );
tran (\sa_count[30][25] , \sa_count[30].f.lower[25] );
tran (\sa_count[30][26] , \sa_count[30].r.part0[26] );
tran (\sa_count[30][26] , \sa_count[30].f.lower[26] );
tran (\sa_count[30][27] , \sa_count[30].r.part0[27] );
tran (\sa_count[30][27] , \sa_count[30].f.lower[27] );
tran (\sa_count[30][28] , \sa_count[30].r.part0[28] );
tran (\sa_count[30][28] , \sa_count[30].f.lower[28] );
tran (\sa_count[30][29] , \sa_count[30].r.part0[29] );
tran (\sa_count[30][29] , \sa_count[30].f.lower[29] );
tran (\sa_count[30][30] , \sa_count[30].r.part0[30] );
tran (\sa_count[30][30] , \sa_count[30].f.lower[30] );
tran (\sa_count[30][31] , \sa_count[30].r.part0[31] );
tran (\sa_count[30][31] , \sa_count[30].f.lower[31] );
tran (\sa_count[30][32] , \sa_count[30].r.part1[0] );
tran (\sa_count[30][32] , \sa_count[30].f.upper[0] );
tran (\sa_count[30][33] , \sa_count[30].r.part1[1] );
tran (\sa_count[30][33] , \sa_count[30].f.upper[1] );
tran (\sa_count[30][34] , \sa_count[30].r.part1[2] );
tran (\sa_count[30][34] , \sa_count[30].f.upper[2] );
tran (\sa_count[30][35] , \sa_count[30].r.part1[3] );
tran (\sa_count[30][35] , \sa_count[30].f.upper[3] );
tran (\sa_count[30][36] , \sa_count[30].r.part1[4] );
tran (\sa_count[30][36] , \sa_count[30].f.upper[4] );
tran (\sa_count[30][37] , \sa_count[30].r.part1[5] );
tran (\sa_count[30][37] , \sa_count[30].f.upper[5] );
tran (\sa_count[30][38] , \sa_count[30].r.part1[6] );
tran (\sa_count[30][38] , \sa_count[30].f.upper[6] );
tran (\sa_count[30][39] , \sa_count[30].r.part1[7] );
tran (\sa_count[30][39] , \sa_count[30].f.upper[7] );
tran (\sa_count[30][40] , \sa_count[30].r.part1[8] );
tran (\sa_count[30][40] , \sa_count[30].f.upper[8] );
tran (\sa_count[30][41] , \sa_count[30].r.part1[9] );
tran (\sa_count[30][41] , \sa_count[30].f.upper[9] );
tran (\sa_count[30][42] , \sa_count[30].r.part1[10] );
tran (\sa_count[30][42] , \sa_count[30].f.upper[10] );
tran (\sa_count[30][43] , \sa_count[30].r.part1[11] );
tran (\sa_count[30][43] , \sa_count[30].f.upper[11] );
tran (\sa_count[30][44] , \sa_count[30].r.part1[12] );
tran (\sa_count[30][44] , \sa_count[30].f.upper[12] );
tran (\sa_count[30][45] , \sa_count[30].r.part1[13] );
tran (\sa_count[30][45] , \sa_count[30].f.upper[13] );
tran (\sa_count[30][46] , \sa_count[30].r.part1[14] );
tran (\sa_count[30][46] , \sa_count[30].f.upper[14] );
tran (\sa_count[30][47] , \sa_count[30].r.part1[15] );
tran (\sa_count[30][47] , \sa_count[30].f.upper[15] );
tran (\sa_count[30][48] , \sa_count[30].r.part1[16] );
tran (\sa_count[30][48] , \sa_count[30].f.upper[16] );
tran (\sa_count[30][49] , \sa_count[30].r.part1[17] );
tran (\sa_count[30][49] , \sa_count[30].f.upper[17] );
tran (\sa_count[30][50] , \sa_count[30].r.part1[18] );
tran (\sa_count[30][50] , \sa_count[30].f.unused[0] );
tran (\sa_count[30][51] , \sa_count[30].r.part1[19] );
tran (\sa_count[30][51] , \sa_count[30].f.unused[1] );
tran (\sa_count[30][52] , \sa_count[30].r.part1[20] );
tran (\sa_count[30][52] , \sa_count[30].f.unused[2] );
tran (\sa_count[30][53] , \sa_count[30].r.part1[21] );
tran (\sa_count[30][53] , \sa_count[30].f.unused[3] );
tran (\sa_count[30][54] , \sa_count[30].r.part1[22] );
tran (\sa_count[30][54] , \sa_count[30].f.unused[4] );
tran (\sa_count[30][55] , \sa_count[30].r.part1[23] );
tran (\sa_count[30][55] , \sa_count[30].f.unused[5] );
tran (\sa_count[30][56] , \sa_count[30].r.part1[24] );
tran (\sa_count[30][56] , \sa_count[30].f.unused[6] );
tran (\sa_count[30][57] , \sa_count[30].r.part1[25] );
tran (\sa_count[30][57] , \sa_count[30].f.unused[7] );
tran (\sa_count[30][58] , \sa_count[30].r.part1[26] );
tran (\sa_count[30][58] , \sa_count[30].f.unused[8] );
tran (\sa_count[30][59] , \sa_count[30].r.part1[27] );
tran (\sa_count[30][59] , \sa_count[30].f.unused[9] );
tran (\sa_count[30][60] , \sa_count[30].r.part1[28] );
tran (\sa_count[30][60] , \sa_count[30].f.unused[10] );
tran (\sa_count[30][61] , \sa_count[30].r.part1[29] );
tran (\sa_count[30][61] , \sa_count[30].f.unused[11] );
tran (\sa_count[30][62] , \sa_count[30].r.part1[30] );
tran (\sa_count[30][62] , \sa_count[30].f.unused[12] );
tran (\sa_count[30][63] , \sa_count[30].r.part1[31] );
tran (\sa_count[30][63] , \sa_count[30].f.unused[13] );
tran (\sa_count[31][0] , \sa_count[31].r.part0[0] );
tran (\sa_count[31][0] , \sa_count[31].f.lower[0] );
tran (\sa_count[31][1] , \sa_count[31].r.part0[1] );
tran (\sa_count[31][1] , \sa_count[31].f.lower[1] );
tran (\sa_count[31][2] , \sa_count[31].r.part0[2] );
tran (\sa_count[31][2] , \sa_count[31].f.lower[2] );
tran (\sa_count[31][3] , \sa_count[31].r.part0[3] );
tran (\sa_count[31][3] , \sa_count[31].f.lower[3] );
tran (\sa_count[31][4] , \sa_count[31].r.part0[4] );
tran (\sa_count[31][4] , \sa_count[31].f.lower[4] );
tran (\sa_count[31][5] , \sa_count[31].r.part0[5] );
tran (\sa_count[31][5] , \sa_count[31].f.lower[5] );
tran (\sa_count[31][6] , \sa_count[31].r.part0[6] );
tran (\sa_count[31][6] , \sa_count[31].f.lower[6] );
tran (\sa_count[31][7] , \sa_count[31].r.part0[7] );
tran (\sa_count[31][7] , \sa_count[31].f.lower[7] );
tran (\sa_count[31][8] , \sa_count[31].r.part0[8] );
tran (\sa_count[31][8] , \sa_count[31].f.lower[8] );
tran (\sa_count[31][9] , \sa_count[31].r.part0[9] );
tran (\sa_count[31][9] , \sa_count[31].f.lower[9] );
tran (\sa_count[31][10] , \sa_count[31].r.part0[10] );
tran (\sa_count[31][10] , \sa_count[31].f.lower[10] );
tran (\sa_count[31][11] , \sa_count[31].r.part0[11] );
tran (\sa_count[31][11] , \sa_count[31].f.lower[11] );
tran (\sa_count[31][12] , \sa_count[31].r.part0[12] );
tran (\sa_count[31][12] , \sa_count[31].f.lower[12] );
tran (\sa_count[31][13] , \sa_count[31].r.part0[13] );
tran (\sa_count[31][13] , \sa_count[31].f.lower[13] );
tran (\sa_count[31][14] , \sa_count[31].r.part0[14] );
tran (\sa_count[31][14] , \sa_count[31].f.lower[14] );
tran (\sa_count[31][15] , \sa_count[31].r.part0[15] );
tran (\sa_count[31][15] , \sa_count[31].f.lower[15] );
tran (\sa_count[31][16] , \sa_count[31].r.part0[16] );
tran (\sa_count[31][16] , \sa_count[31].f.lower[16] );
tran (\sa_count[31][17] , \sa_count[31].r.part0[17] );
tran (\sa_count[31][17] , \sa_count[31].f.lower[17] );
tran (\sa_count[31][18] , \sa_count[31].r.part0[18] );
tran (\sa_count[31][18] , \sa_count[31].f.lower[18] );
tran (\sa_count[31][19] , \sa_count[31].r.part0[19] );
tran (\sa_count[31][19] , \sa_count[31].f.lower[19] );
tran (\sa_count[31][20] , \sa_count[31].r.part0[20] );
tran (\sa_count[31][20] , \sa_count[31].f.lower[20] );
tran (\sa_count[31][21] , \sa_count[31].r.part0[21] );
tran (\sa_count[31][21] , \sa_count[31].f.lower[21] );
tran (\sa_count[31][22] , \sa_count[31].r.part0[22] );
tran (\sa_count[31][22] , \sa_count[31].f.lower[22] );
tran (\sa_count[31][23] , \sa_count[31].r.part0[23] );
tran (\sa_count[31][23] , \sa_count[31].f.lower[23] );
tran (\sa_count[31][24] , \sa_count[31].r.part0[24] );
tran (\sa_count[31][24] , \sa_count[31].f.lower[24] );
tran (\sa_count[31][25] , \sa_count[31].r.part0[25] );
tran (\sa_count[31][25] , \sa_count[31].f.lower[25] );
tran (\sa_count[31][26] , \sa_count[31].r.part0[26] );
tran (\sa_count[31][26] , \sa_count[31].f.lower[26] );
tran (\sa_count[31][27] , \sa_count[31].r.part0[27] );
tran (\sa_count[31][27] , \sa_count[31].f.lower[27] );
tran (\sa_count[31][28] , \sa_count[31].r.part0[28] );
tran (\sa_count[31][28] , \sa_count[31].f.lower[28] );
tran (\sa_count[31][29] , \sa_count[31].r.part0[29] );
tran (\sa_count[31][29] , \sa_count[31].f.lower[29] );
tran (\sa_count[31][30] , \sa_count[31].r.part0[30] );
tran (\sa_count[31][30] , \sa_count[31].f.lower[30] );
tran (\sa_count[31][31] , \sa_count[31].r.part0[31] );
tran (\sa_count[31][31] , \sa_count[31].f.lower[31] );
tran (\sa_count[31][32] , \sa_count[31].r.part1[0] );
tran (\sa_count[31][32] , \sa_count[31].f.upper[0] );
tran (\sa_count[31][33] , \sa_count[31].r.part1[1] );
tran (\sa_count[31][33] , \sa_count[31].f.upper[1] );
tran (\sa_count[31][34] , \sa_count[31].r.part1[2] );
tran (\sa_count[31][34] , \sa_count[31].f.upper[2] );
tran (\sa_count[31][35] , \sa_count[31].r.part1[3] );
tran (\sa_count[31][35] , \sa_count[31].f.upper[3] );
tran (\sa_count[31][36] , \sa_count[31].r.part1[4] );
tran (\sa_count[31][36] , \sa_count[31].f.upper[4] );
tran (\sa_count[31][37] , \sa_count[31].r.part1[5] );
tran (\sa_count[31][37] , \sa_count[31].f.upper[5] );
tran (\sa_count[31][38] , \sa_count[31].r.part1[6] );
tran (\sa_count[31][38] , \sa_count[31].f.upper[6] );
tran (\sa_count[31][39] , \sa_count[31].r.part1[7] );
tran (\sa_count[31][39] , \sa_count[31].f.upper[7] );
tran (\sa_count[31][40] , \sa_count[31].r.part1[8] );
tran (\sa_count[31][40] , \sa_count[31].f.upper[8] );
tran (\sa_count[31][41] , \sa_count[31].r.part1[9] );
tran (\sa_count[31][41] , \sa_count[31].f.upper[9] );
tran (\sa_count[31][42] , \sa_count[31].r.part1[10] );
tran (\sa_count[31][42] , \sa_count[31].f.upper[10] );
tran (\sa_count[31][43] , \sa_count[31].r.part1[11] );
tran (\sa_count[31][43] , \sa_count[31].f.upper[11] );
tran (\sa_count[31][44] , \sa_count[31].r.part1[12] );
tran (\sa_count[31][44] , \sa_count[31].f.upper[12] );
tran (\sa_count[31][45] , \sa_count[31].r.part1[13] );
tran (\sa_count[31][45] , \sa_count[31].f.upper[13] );
tran (\sa_count[31][46] , \sa_count[31].r.part1[14] );
tran (\sa_count[31][46] , \sa_count[31].f.upper[14] );
tran (\sa_count[31][47] , \sa_count[31].r.part1[15] );
tran (\sa_count[31][47] , \sa_count[31].f.upper[15] );
tran (\sa_count[31][48] , \sa_count[31].r.part1[16] );
tran (\sa_count[31][48] , \sa_count[31].f.upper[16] );
tran (\sa_count[31][49] , \sa_count[31].r.part1[17] );
tran (\sa_count[31][49] , \sa_count[31].f.upper[17] );
tran (\sa_count[31][50] , \sa_count[31].r.part1[18] );
tran (\sa_count[31][50] , \sa_count[31].f.unused[0] );
tran (\sa_count[31][51] , \sa_count[31].r.part1[19] );
tran (\sa_count[31][51] , \sa_count[31].f.unused[1] );
tran (\sa_count[31][52] , \sa_count[31].r.part1[20] );
tran (\sa_count[31][52] , \sa_count[31].f.unused[2] );
tran (\sa_count[31][53] , \sa_count[31].r.part1[21] );
tran (\sa_count[31][53] , \sa_count[31].f.unused[3] );
tran (\sa_count[31][54] , \sa_count[31].r.part1[22] );
tran (\sa_count[31][54] , \sa_count[31].f.unused[4] );
tran (\sa_count[31][55] , \sa_count[31].r.part1[23] );
tran (\sa_count[31][55] , \sa_count[31].f.unused[5] );
tran (\sa_count[31][56] , \sa_count[31].r.part1[24] );
tran (\sa_count[31][56] , \sa_count[31].f.unused[6] );
tran (\sa_count[31][57] , \sa_count[31].r.part1[25] );
tran (\sa_count[31][57] , \sa_count[31].f.unused[7] );
tran (\sa_count[31][58] , \sa_count[31].r.part1[26] );
tran (\sa_count[31][58] , \sa_count[31].f.unused[8] );
tran (\sa_count[31][59] , \sa_count[31].r.part1[27] );
tran (\sa_count[31][59] , \sa_count[31].f.unused[9] );
tran (\sa_count[31][60] , \sa_count[31].r.part1[28] );
tran (\sa_count[31][60] , \sa_count[31].f.unused[10] );
tran (\sa_count[31][61] , \sa_count[31].r.part1[29] );
tran (\sa_count[31][61] , \sa_count[31].f.unused[11] );
tran (\sa_count[31][62] , \sa_count[31].r.part1[30] );
tran (\sa_count[31][62] , \sa_count[31].f.unused[12] );
tran (\sa_count[31][63] , \sa_count[31].r.part1[31] );
tran (\sa_count[31][63] , \sa_count[31].f.unused[13] );
tran (cddip3_im_din[6], \cddip3_im_din.desc.im_meta [6]);
tran (cddip3_im_din[8], \cddip3_im_din.desc.im_meta [8]);
tran (cddip3_im_din[9], \cddip3_im_din.desc.im_meta [9]);
tran (cddip3_im_din[10], \cddip3_im_din.desc.im_meta [10]);
tran (cddip3_im_din[11], \cddip3_im_din.desc.im_meta [11]);
tran (cddip3_im_din[12], \cddip3_im_din.desc.im_meta [12]);
tran (cddip3_im_din[13], \cddip3_im_din.desc.im_meta [13]);
tran (cddip3_im_din[14], \cddip3_im_din.desc.im_meta [14]);
tran (cddip3_im_din[23], \cddip3_im_din.desc.bytes_vld [0]);
tran (cddip3_im_din[24], \cddip3_im_din.desc.bytes_vld [1]);
tran (cddip3_im_din[25], \cddip3_im_din.desc.bytes_vld [2]);
tran (cddip3_im_din[26], \cddip3_im_din.desc.bytes_vld [3]);
tran (cddip3_im_din[27], \cddip3_im_din.desc.bytes_vld [4]);
tran (cddip3_im_din[28], \cddip3_im_din.desc.bytes_vld [5]);
tran (cddip3_im_din[29], \cddip3_im_din.desc.bytes_vld [6]);
tran (cddip3_im_din[30], \cddip3_im_din.desc.bytes_vld [7]);
tran (cddip3_im_din[31], \cddip3_im_din.desc.eob );
tran (cddip3_im_din[7], \cddip3_im_din.desc.im_meta [7]);
tran (cddip3_im_din[32], \cddip3_im_din.data.data [0]);
tran (cddip3_im_din[33], \cddip3_im_din.data.data [1]);
tran (cddip3_im_din[34], \cddip3_im_din.data.data [2]);
tran (cddip3_im_din[35], \cddip3_im_din.data.data [3]);
tran (cddip3_im_din[36], \cddip3_im_din.data.data [4]);
tran (cddip3_im_din[37], \cddip3_im_din.data.data [5]);
tran (cddip3_im_din[38], \cddip3_im_din.data.data [6]);
tran (cddip3_im_din[39], \cddip3_im_din.data.data [7]);
tran (cddip3_im_din[40], \cddip3_im_din.data.data [8]);
tran (cddip3_im_din[41], \cddip3_im_din.data.data [9]);
tran (cddip3_im_din[42], \cddip3_im_din.data.data [10]);
tran (cddip3_im_din[43], \cddip3_im_din.data.data [11]);
tran (cddip3_im_din[44], \cddip3_im_din.data.data [12]);
tran (cddip3_im_din[45], \cddip3_im_din.data.data [13]);
tran (cddip3_im_din[46], \cddip3_im_din.data.data [14]);
tran (cddip3_im_din[47], \cddip3_im_din.data.data [15]);
tran (cddip3_im_din[48], \cddip3_im_din.data.data [16]);
tran (cddip3_im_din[49], \cddip3_im_din.data.data [17]);
tran (cddip3_im_din[50], \cddip3_im_din.data.data [18]);
tran (cddip3_im_din[51], \cddip3_im_din.data.data [19]);
tran (cddip3_im_din[52], \cddip3_im_din.data.data [20]);
tran (cddip3_im_din[53], \cddip3_im_din.data.data [21]);
tran (cddip3_im_din[54], \cddip3_im_din.data.data [22]);
tran (cddip3_im_din[55], \cddip3_im_din.data.data [23]);
tran (cddip3_im_din[56], \cddip3_im_din.data.data [24]);
tran (cddip3_im_din[57], \cddip3_im_din.data.data [25]);
tran (cddip3_im_din[58], \cddip3_im_din.data.data [26]);
tran (cddip3_im_din[59], \cddip3_im_din.data.data [27]);
tran (cddip3_im_din[60], \cddip3_im_din.data.data [28]);
tran (cddip3_im_din[61], \cddip3_im_din.data.data [29]);
tran (cddip3_im_din[62], \cddip3_im_din.data.data [30]);
tran (cddip3_im_din[63], \cddip3_im_din.data.data [31]);
tran (cddip3_im_din[64], \cddip3_im_din.data.data [32]);
tran (cddip3_im_din[65], \cddip3_im_din.data.data [33]);
tran (cddip3_im_din[66], \cddip3_im_din.data.data [34]);
tran (cddip3_im_din[67], \cddip3_im_din.data.data [35]);
tran (cddip3_im_din[68], \cddip3_im_din.data.data [36]);
tran (cddip3_im_din[69], \cddip3_im_din.data.data [37]);
tran (cddip3_im_din[70], \cddip3_im_din.data.data [38]);
tran (cddip3_im_din[71], \cddip3_im_din.data.data [39]);
tran (cddip3_im_din[72], \cddip3_im_din.data.data [40]);
tran (cddip3_im_din[73], \cddip3_im_din.data.data [41]);
tran (cddip3_im_din[74], \cddip3_im_din.data.data [42]);
tran (cddip3_im_din[75], \cddip3_im_din.data.data [43]);
tran (cddip3_im_din[76], \cddip3_im_din.data.data [44]);
tran (cddip3_im_din[77], \cddip3_im_din.data.data [45]);
tran (cddip3_im_din[78], \cddip3_im_din.data.data [46]);
tran (cddip3_im_din[79], \cddip3_im_din.data.data [47]);
tran (cddip3_im_din[80], \cddip3_im_din.data.data [48]);
tran (cddip3_im_din[81], \cddip3_im_din.data.data [49]);
tran (cddip3_im_din[82], \cddip3_im_din.data.data [50]);
tran (cddip3_im_din[83], \cddip3_im_din.data.data [51]);
tran (cddip3_im_din[84], \cddip3_im_din.data.data [52]);
tran (cddip3_im_din[85], \cddip3_im_din.data.data [53]);
tran (cddip3_im_din[86], \cddip3_im_din.data.data [54]);
tran (cddip3_im_din[87], \cddip3_im_din.data.data [55]);
tran (cddip3_im_din[88], \cddip3_im_din.data.data [56]);
tran (cddip3_im_din[89], \cddip3_im_din.data.data [57]);
tran (cddip3_im_din[90], \cddip3_im_din.data.data [58]);
tran (cddip3_im_din[91], \cddip3_im_din.data.data [59]);
tran (cddip3_im_din[92], \cddip3_im_din.data.data [60]);
tran (cddip3_im_din[93], \cddip3_im_din.data.data [61]);
tran (cddip3_im_din[94], \cddip3_im_din.data.data [62]);
tran (cddip3_im_din[95], \cddip3_im_din.data.data [63]);
tran (cceip3_im_din[6], \cceip3_im_din.desc.im_meta [6]);
tran (cceip3_im_din[8], \cceip3_im_din.desc.im_meta [8]);
tran (cceip3_im_din[9], \cceip3_im_din.desc.im_meta [9]);
tran (cceip3_im_din[10], \cceip3_im_din.desc.im_meta [10]);
tran (cceip3_im_din[11], \cceip3_im_din.desc.im_meta [11]);
tran (cceip3_im_din[12], \cceip3_im_din.desc.im_meta [12]);
tran (cceip3_im_din[13], \cceip3_im_din.desc.im_meta [13]);
tran (cceip3_im_din[14], \cceip3_im_din.desc.im_meta [14]);
tran (cceip3_im_din[23], \cceip3_im_din.desc.bytes_vld [0]);
tran (cceip3_im_din[24], \cceip3_im_din.desc.bytes_vld [1]);
tran (cceip3_im_din[25], \cceip3_im_din.desc.bytes_vld [2]);
tran (cceip3_im_din[26], \cceip3_im_din.desc.bytes_vld [3]);
tran (cceip3_im_din[27], \cceip3_im_din.desc.bytes_vld [4]);
tran (cceip3_im_din[28], \cceip3_im_din.desc.bytes_vld [5]);
tran (cceip3_im_din[29], \cceip3_im_din.desc.bytes_vld [6]);
tran (cceip3_im_din[30], \cceip3_im_din.desc.bytes_vld [7]);
tran (cceip3_im_din[31], \cceip3_im_din.desc.eob );
tran (cceip3_im_din[7], \cceip3_im_din.desc.im_meta [7]);
tran (cceip3_im_din[32], \cceip3_im_din.data.data [0]);
tran (cceip3_im_din[33], \cceip3_im_din.data.data [1]);
tran (cceip3_im_din[34], \cceip3_im_din.data.data [2]);
tran (cceip3_im_din[35], \cceip3_im_din.data.data [3]);
tran (cceip3_im_din[36], \cceip3_im_din.data.data [4]);
tran (cceip3_im_din[37], \cceip3_im_din.data.data [5]);
tran (cceip3_im_din[38], \cceip3_im_din.data.data [6]);
tran (cceip3_im_din[39], \cceip3_im_din.data.data [7]);
tran (cceip3_im_din[40], \cceip3_im_din.data.data [8]);
tran (cceip3_im_din[41], \cceip3_im_din.data.data [9]);
tran (cceip3_im_din[42], \cceip3_im_din.data.data [10]);
tran (cceip3_im_din[43], \cceip3_im_din.data.data [11]);
tran (cceip3_im_din[44], \cceip3_im_din.data.data [12]);
tran (cceip3_im_din[45], \cceip3_im_din.data.data [13]);
tran (cceip3_im_din[46], \cceip3_im_din.data.data [14]);
tran (cceip3_im_din[47], \cceip3_im_din.data.data [15]);
tran (cceip3_im_din[48], \cceip3_im_din.data.data [16]);
tran (cceip3_im_din[49], \cceip3_im_din.data.data [17]);
tran (cceip3_im_din[50], \cceip3_im_din.data.data [18]);
tran (cceip3_im_din[51], \cceip3_im_din.data.data [19]);
tran (cceip3_im_din[52], \cceip3_im_din.data.data [20]);
tran (cceip3_im_din[53], \cceip3_im_din.data.data [21]);
tran (cceip3_im_din[54], \cceip3_im_din.data.data [22]);
tran (cceip3_im_din[55], \cceip3_im_din.data.data [23]);
tran (cceip3_im_din[56], \cceip3_im_din.data.data [24]);
tran (cceip3_im_din[57], \cceip3_im_din.data.data [25]);
tran (cceip3_im_din[58], \cceip3_im_din.data.data [26]);
tran (cceip3_im_din[59], \cceip3_im_din.data.data [27]);
tran (cceip3_im_din[60], \cceip3_im_din.data.data [28]);
tran (cceip3_im_din[61], \cceip3_im_din.data.data [29]);
tran (cceip3_im_din[62], \cceip3_im_din.data.data [30]);
tran (cceip3_im_din[63], \cceip3_im_din.data.data [31]);
tran (cceip3_im_din[64], \cceip3_im_din.data.data [32]);
tran (cceip3_im_din[65], \cceip3_im_din.data.data [33]);
tran (cceip3_im_din[66], \cceip3_im_din.data.data [34]);
tran (cceip3_im_din[67], \cceip3_im_din.data.data [35]);
tran (cceip3_im_din[68], \cceip3_im_din.data.data [36]);
tran (cceip3_im_din[69], \cceip3_im_din.data.data [37]);
tran (cceip3_im_din[70], \cceip3_im_din.data.data [38]);
tran (cceip3_im_din[71], \cceip3_im_din.data.data [39]);
tran (cceip3_im_din[72], \cceip3_im_din.data.data [40]);
tran (cceip3_im_din[73], \cceip3_im_din.data.data [41]);
tran (cceip3_im_din[74], \cceip3_im_din.data.data [42]);
tran (cceip3_im_din[75], \cceip3_im_din.data.data [43]);
tran (cceip3_im_din[76], \cceip3_im_din.data.data [44]);
tran (cceip3_im_din[77], \cceip3_im_din.data.data [45]);
tran (cceip3_im_din[78], \cceip3_im_din.data.data [46]);
tran (cceip3_im_din[79], \cceip3_im_din.data.data [47]);
tran (cceip3_im_din[80], \cceip3_im_din.data.data [48]);
tran (cceip3_im_din[81], \cceip3_im_din.data.data [49]);
tran (cceip3_im_din[82], \cceip3_im_din.data.data [50]);
tran (cceip3_im_din[83], \cceip3_im_din.data.data [51]);
tran (cceip3_im_din[84], \cceip3_im_din.data.data [52]);
tran (cceip3_im_din[85], \cceip3_im_din.data.data [53]);
tran (cceip3_im_din[86], \cceip3_im_din.data.data [54]);
tran (cceip3_im_din[87], \cceip3_im_din.data.data [55]);
tran (cceip3_im_din[88], \cceip3_im_din.data.data [56]);
tran (cceip3_im_din[89], \cceip3_im_din.data.data [57]);
tran (cceip3_im_din[90], \cceip3_im_din.data.data [58]);
tran (cceip3_im_din[91], \cceip3_im_din.data.data [59]);
tran (cceip3_im_din[92], \cceip3_im_din.data.data [60]);
tran (cceip3_im_din[93], \cceip3_im_din.data.data [61]);
tran (cceip3_im_din[94], \cceip3_im_din.data.data [62]);
tran (cceip3_im_din[95], \cceip3_im_din.data.data [63]);
tran (cddip2_im_din[6], \cddip2_im_din.desc.im_meta [6]);
tran (cddip2_im_din[8], \cddip2_im_din.desc.im_meta [8]);
tran (cddip2_im_din[9], \cddip2_im_din.desc.im_meta [9]);
tran (cddip2_im_din[10], \cddip2_im_din.desc.im_meta [10]);
tran (cddip2_im_din[11], \cddip2_im_din.desc.im_meta [11]);
tran (cddip2_im_din[12], \cddip2_im_din.desc.im_meta [12]);
tran (cddip2_im_din[13], \cddip2_im_din.desc.im_meta [13]);
tran (cddip2_im_din[14], \cddip2_im_din.desc.im_meta [14]);
tran (cddip2_im_din[23], \cddip2_im_din.desc.bytes_vld [0]);
tran (cddip2_im_din[24], \cddip2_im_din.desc.bytes_vld [1]);
tran (cddip2_im_din[25], \cddip2_im_din.desc.bytes_vld [2]);
tran (cddip2_im_din[26], \cddip2_im_din.desc.bytes_vld [3]);
tran (cddip2_im_din[27], \cddip2_im_din.desc.bytes_vld [4]);
tran (cddip2_im_din[28], \cddip2_im_din.desc.bytes_vld [5]);
tran (cddip2_im_din[29], \cddip2_im_din.desc.bytes_vld [6]);
tran (cddip2_im_din[30], \cddip2_im_din.desc.bytes_vld [7]);
tran (cddip2_im_din[31], \cddip2_im_din.desc.eob );
tran (cddip2_im_din[7], \cddip2_im_din.desc.im_meta [7]);
tran (cddip2_im_din[32], \cddip2_im_din.data.data [0]);
tran (cddip2_im_din[33], \cddip2_im_din.data.data [1]);
tran (cddip2_im_din[34], \cddip2_im_din.data.data [2]);
tran (cddip2_im_din[35], \cddip2_im_din.data.data [3]);
tran (cddip2_im_din[36], \cddip2_im_din.data.data [4]);
tran (cddip2_im_din[37], \cddip2_im_din.data.data [5]);
tran (cddip2_im_din[38], \cddip2_im_din.data.data [6]);
tran (cddip2_im_din[39], \cddip2_im_din.data.data [7]);
tran (cddip2_im_din[40], \cddip2_im_din.data.data [8]);
tran (cddip2_im_din[41], \cddip2_im_din.data.data [9]);
tran (cddip2_im_din[42], \cddip2_im_din.data.data [10]);
tran (cddip2_im_din[43], \cddip2_im_din.data.data [11]);
tran (cddip2_im_din[44], \cddip2_im_din.data.data [12]);
tran (cddip2_im_din[45], \cddip2_im_din.data.data [13]);
tran (cddip2_im_din[46], \cddip2_im_din.data.data [14]);
tran (cddip2_im_din[47], \cddip2_im_din.data.data [15]);
tran (cddip2_im_din[48], \cddip2_im_din.data.data [16]);
tran (cddip2_im_din[49], \cddip2_im_din.data.data [17]);
tran (cddip2_im_din[50], \cddip2_im_din.data.data [18]);
tran (cddip2_im_din[51], \cddip2_im_din.data.data [19]);
tran (cddip2_im_din[52], \cddip2_im_din.data.data [20]);
tran (cddip2_im_din[53], \cddip2_im_din.data.data [21]);
tran (cddip2_im_din[54], \cddip2_im_din.data.data [22]);
tran (cddip2_im_din[55], \cddip2_im_din.data.data [23]);
tran (cddip2_im_din[56], \cddip2_im_din.data.data [24]);
tran (cddip2_im_din[57], \cddip2_im_din.data.data [25]);
tran (cddip2_im_din[58], \cddip2_im_din.data.data [26]);
tran (cddip2_im_din[59], \cddip2_im_din.data.data [27]);
tran (cddip2_im_din[60], \cddip2_im_din.data.data [28]);
tran (cddip2_im_din[61], \cddip2_im_din.data.data [29]);
tran (cddip2_im_din[62], \cddip2_im_din.data.data [30]);
tran (cddip2_im_din[63], \cddip2_im_din.data.data [31]);
tran (cddip2_im_din[64], \cddip2_im_din.data.data [32]);
tran (cddip2_im_din[65], \cddip2_im_din.data.data [33]);
tran (cddip2_im_din[66], \cddip2_im_din.data.data [34]);
tran (cddip2_im_din[67], \cddip2_im_din.data.data [35]);
tran (cddip2_im_din[68], \cddip2_im_din.data.data [36]);
tran (cddip2_im_din[69], \cddip2_im_din.data.data [37]);
tran (cddip2_im_din[70], \cddip2_im_din.data.data [38]);
tran (cddip2_im_din[71], \cddip2_im_din.data.data [39]);
tran (cddip2_im_din[72], \cddip2_im_din.data.data [40]);
tran (cddip2_im_din[73], \cddip2_im_din.data.data [41]);
tran (cddip2_im_din[74], \cddip2_im_din.data.data [42]);
tran (cddip2_im_din[75], \cddip2_im_din.data.data [43]);
tran (cddip2_im_din[76], \cddip2_im_din.data.data [44]);
tran (cddip2_im_din[77], \cddip2_im_din.data.data [45]);
tran (cddip2_im_din[78], \cddip2_im_din.data.data [46]);
tran (cddip2_im_din[79], \cddip2_im_din.data.data [47]);
tran (cddip2_im_din[80], \cddip2_im_din.data.data [48]);
tran (cddip2_im_din[81], \cddip2_im_din.data.data [49]);
tran (cddip2_im_din[82], \cddip2_im_din.data.data [50]);
tran (cddip2_im_din[83], \cddip2_im_din.data.data [51]);
tran (cddip2_im_din[84], \cddip2_im_din.data.data [52]);
tran (cddip2_im_din[85], \cddip2_im_din.data.data [53]);
tran (cddip2_im_din[86], \cddip2_im_din.data.data [54]);
tran (cddip2_im_din[87], \cddip2_im_din.data.data [55]);
tran (cddip2_im_din[88], \cddip2_im_din.data.data [56]);
tran (cddip2_im_din[89], \cddip2_im_din.data.data [57]);
tran (cddip2_im_din[90], \cddip2_im_din.data.data [58]);
tran (cddip2_im_din[91], \cddip2_im_din.data.data [59]);
tran (cddip2_im_din[92], \cddip2_im_din.data.data [60]);
tran (cddip2_im_din[93], \cddip2_im_din.data.data [61]);
tran (cddip2_im_din[94], \cddip2_im_din.data.data [62]);
tran (cddip2_im_din[95], \cddip2_im_din.data.data [63]);
tran (cceip2_im_din[6], \cceip2_im_din.desc.im_meta [6]);
tran (cceip2_im_din[8], \cceip2_im_din.desc.im_meta [8]);
tran (cceip2_im_din[9], \cceip2_im_din.desc.im_meta [9]);
tran (cceip2_im_din[10], \cceip2_im_din.desc.im_meta [10]);
tran (cceip2_im_din[11], \cceip2_im_din.desc.im_meta [11]);
tran (cceip2_im_din[12], \cceip2_im_din.desc.im_meta [12]);
tran (cceip2_im_din[13], \cceip2_im_din.desc.im_meta [13]);
tran (cceip2_im_din[14], \cceip2_im_din.desc.im_meta [14]);
tran (cceip2_im_din[23], \cceip2_im_din.desc.bytes_vld [0]);
tran (cceip2_im_din[24], \cceip2_im_din.desc.bytes_vld [1]);
tran (cceip2_im_din[25], \cceip2_im_din.desc.bytes_vld [2]);
tran (cceip2_im_din[26], \cceip2_im_din.desc.bytes_vld [3]);
tran (cceip2_im_din[27], \cceip2_im_din.desc.bytes_vld [4]);
tran (cceip2_im_din[28], \cceip2_im_din.desc.bytes_vld [5]);
tran (cceip2_im_din[29], \cceip2_im_din.desc.bytes_vld [6]);
tran (cceip2_im_din[30], \cceip2_im_din.desc.bytes_vld [7]);
tran (cceip2_im_din[31], \cceip2_im_din.desc.eob );
tran (cceip2_im_din[7], \cceip2_im_din.desc.im_meta [7]);
tran (cceip2_im_din[32], \cceip2_im_din.data.data [0]);
tran (cceip2_im_din[33], \cceip2_im_din.data.data [1]);
tran (cceip2_im_din[34], \cceip2_im_din.data.data [2]);
tran (cceip2_im_din[35], \cceip2_im_din.data.data [3]);
tran (cceip2_im_din[36], \cceip2_im_din.data.data [4]);
tran (cceip2_im_din[37], \cceip2_im_din.data.data [5]);
tran (cceip2_im_din[38], \cceip2_im_din.data.data [6]);
tran (cceip2_im_din[39], \cceip2_im_din.data.data [7]);
tran (cceip2_im_din[40], \cceip2_im_din.data.data [8]);
tran (cceip2_im_din[41], \cceip2_im_din.data.data [9]);
tran (cceip2_im_din[42], \cceip2_im_din.data.data [10]);
tran (cceip2_im_din[43], \cceip2_im_din.data.data [11]);
tran (cceip2_im_din[44], \cceip2_im_din.data.data [12]);
tran (cceip2_im_din[45], \cceip2_im_din.data.data [13]);
tran (cceip2_im_din[46], \cceip2_im_din.data.data [14]);
tran (cceip2_im_din[47], \cceip2_im_din.data.data [15]);
tran (cceip2_im_din[48], \cceip2_im_din.data.data [16]);
tran (cceip2_im_din[49], \cceip2_im_din.data.data [17]);
tran (cceip2_im_din[50], \cceip2_im_din.data.data [18]);
tran (cceip2_im_din[51], \cceip2_im_din.data.data [19]);
tran (cceip2_im_din[52], \cceip2_im_din.data.data [20]);
tran (cceip2_im_din[53], \cceip2_im_din.data.data [21]);
tran (cceip2_im_din[54], \cceip2_im_din.data.data [22]);
tran (cceip2_im_din[55], \cceip2_im_din.data.data [23]);
tran (cceip2_im_din[56], \cceip2_im_din.data.data [24]);
tran (cceip2_im_din[57], \cceip2_im_din.data.data [25]);
tran (cceip2_im_din[58], \cceip2_im_din.data.data [26]);
tran (cceip2_im_din[59], \cceip2_im_din.data.data [27]);
tran (cceip2_im_din[60], \cceip2_im_din.data.data [28]);
tran (cceip2_im_din[61], \cceip2_im_din.data.data [29]);
tran (cceip2_im_din[62], \cceip2_im_din.data.data [30]);
tran (cceip2_im_din[63], \cceip2_im_din.data.data [31]);
tran (cceip2_im_din[64], \cceip2_im_din.data.data [32]);
tran (cceip2_im_din[65], \cceip2_im_din.data.data [33]);
tran (cceip2_im_din[66], \cceip2_im_din.data.data [34]);
tran (cceip2_im_din[67], \cceip2_im_din.data.data [35]);
tran (cceip2_im_din[68], \cceip2_im_din.data.data [36]);
tran (cceip2_im_din[69], \cceip2_im_din.data.data [37]);
tran (cceip2_im_din[70], \cceip2_im_din.data.data [38]);
tran (cceip2_im_din[71], \cceip2_im_din.data.data [39]);
tran (cceip2_im_din[72], \cceip2_im_din.data.data [40]);
tran (cceip2_im_din[73], \cceip2_im_din.data.data [41]);
tran (cceip2_im_din[74], \cceip2_im_din.data.data [42]);
tran (cceip2_im_din[75], \cceip2_im_din.data.data [43]);
tran (cceip2_im_din[76], \cceip2_im_din.data.data [44]);
tran (cceip2_im_din[77], \cceip2_im_din.data.data [45]);
tran (cceip2_im_din[78], \cceip2_im_din.data.data [46]);
tran (cceip2_im_din[79], \cceip2_im_din.data.data [47]);
tran (cceip2_im_din[80], \cceip2_im_din.data.data [48]);
tran (cceip2_im_din[81], \cceip2_im_din.data.data [49]);
tran (cceip2_im_din[82], \cceip2_im_din.data.data [50]);
tran (cceip2_im_din[83], \cceip2_im_din.data.data [51]);
tran (cceip2_im_din[84], \cceip2_im_din.data.data [52]);
tran (cceip2_im_din[85], \cceip2_im_din.data.data [53]);
tran (cceip2_im_din[86], \cceip2_im_din.data.data [54]);
tran (cceip2_im_din[87], \cceip2_im_din.data.data [55]);
tran (cceip2_im_din[88], \cceip2_im_din.data.data [56]);
tran (cceip2_im_din[89], \cceip2_im_din.data.data [57]);
tran (cceip2_im_din[90], \cceip2_im_din.data.data [58]);
tran (cceip2_im_din[91], \cceip2_im_din.data.data [59]);
tran (cceip2_im_din[92], \cceip2_im_din.data.data [60]);
tran (cceip2_im_din[93], \cceip2_im_din.data.data [61]);
tran (cceip2_im_din[94], \cceip2_im_din.data.data [62]);
tran (cceip2_im_din[95], \cceip2_im_din.data.data [63]);
tran (cddip1_im_din[6], \cddip1_im_din.desc.im_meta [6]);
tran (cddip1_im_din[8], \cddip1_im_din.desc.im_meta [8]);
tran (cddip1_im_din[9], \cddip1_im_din.desc.im_meta [9]);
tran (cddip1_im_din[10], \cddip1_im_din.desc.im_meta [10]);
tran (cddip1_im_din[11], \cddip1_im_din.desc.im_meta [11]);
tran (cddip1_im_din[12], \cddip1_im_din.desc.im_meta [12]);
tran (cddip1_im_din[13], \cddip1_im_din.desc.im_meta [13]);
tran (cddip1_im_din[14], \cddip1_im_din.desc.im_meta [14]);
tran (cddip1_im_din[23], \cddip1_im_din.desc.bytes_vld [0]);
tran (cddip1_im_din[24], \cddip1_im_din.desc.bytes_vld [1]);
tran (cddip1_im_din[25], \cddip1_im_din.desc.bytes_vld [2]);
tran (cddip1_im_din[26], \cddip1_im_din.desc.bytes_vld [3]);
tran (cddip1_im_din[27], \cddip1_im_din.desc.bytes_vld [4]);
tran (cddip1_im_din[28], \cddip1_im_din.desc.bytes_vld [5]);
tran (cddip1_im_din[29], \cddip1_im_din.desc.bytes_vld [6]);
tran (cddip1_im_din[30], \cddip1_im_din.desc.bytes_vld [7]);
tran (cddip1_im_din[31], \cddip1_im_din.desc.eob );
tran (cddip1_im_din[7], \cddip1_im_din.desc.im_meta [7]);
tran (cddip1_im_din[32], \cddip1_im_din.data.data [0]);
tran (cddip1_im_din[33], \cddip1_im_din.data.data [1]);
tran (cddip1_im_din[34], \cddip1_im_din.data.data [2]);
tran (cddip1_im_din[35], \cddip1_im_din.data.data [3]);
tran (cddip1_im_din[36], \cddip1_im_din.data.data [4]);
tran (cddip1_im_din[37], \cddip1_im_din.data.data [5]);
tran (cddip1_im_din[38], \cddip1_im_din.data.data [6]);
tran (cddip1_im_din[39], \cddip1_im_din.data.data [7]);
tran (cddip1_im_din[40], \cddip1_im_din.data.data [8]);
tran (cddip1_im_din[41], \cddip1_im_din.data.data [9]);
tran (cddip1_im_din[42], \cddip1_im_din.data.data [10]);
tran (cddip1_im_din[43], \cddip1_im_din.data.data [11]);
tran (cddip1_im_din[44], \cddip1_im_din.data.data [12]);
tran (cddip1_im_din[45], \cddip1_im_din.data.data [13]);
tran (cddip1_im_din[46], \cddip1_im_din.data.data [14]);
tran (cddip1_im_din[47], \cddip1_im_din.data.data [15]);
tran (cddip1_im_din[48], \cddip1_im_din.data.data [16]);
tran (cddip1_im_din[49], \cddip1_im_din.data.data [17]);
tran (cddip1_im_din[50], \cddip1_im_din.data.data [18]);
tran (cddip1_im_din[51], \cddip1_im_din.data.data [19]);
tran (cddip1_im_din[52], \cddip1_im_din.data.data [20]);
tran (cddip1_im_din[53], \cddip1_im_din.data.data [21]);
tran (cddip1_im_din[54], \cddip1_im_din.data.data [22]);
tran (cddip1_im_din[55], \cddip1_im_din.data.data [23]);
tran (cddip1_im_din[56], \cddip1_im_din.data.data [24]);
tran (cddip1_im_din[57], \cddip1_im_din.data.data [25]);
tran (cddip1_im_din[58], \cddip1_im_din.data.data [26]);
tran (cddip1_im_din[59], \cddip1_im_din.data.data [27]);
tran (cddip1_im_din[60], \cddip1_im_din.data.data [28]);
tran (cddip1_im_din[61], \cddip1_im_din.data.data [29]);
tran (cddip1_im_din[62], \cddip1_im_din.data.data [30]);
tran (cddip1_im_din[63], \cddip1_im_din.data.data [31]);
tran (cddip1_im_din[64], \cddip1_im_din.data.data [32]);
tran (cddip1_im_din[65], \cddip1_im_din.data.data [33]);
tran (cddip1_im_din[66], \cddip1_im_din.data.data [34]);
tran (cddip1_im_din[67], \cddip1_im_din.data.data [35]);
tran (cddip1_im_din[68], \cddip1_im_din.data.data [36]);
tran (cddip1_im_din[69], \cddip1_im_din.data.data [37]);
tran (cddip1_im_din[70], \cddip1_im_din.data.data [38]);
tran (cddip1_im_din[71], \cddip1_im_din.data.data [39]);
tran (cddip1_im_din[72], \cddip1_im_din.data.data [40]);
tran (cddip1_im_din[73], \cddip1_im_din.data.data [41]);
tran (cddip1_im_din[74], \cddip1_im_din.data.data [42]);
tran (cddip1_im_din[75], \cddip1_im_din.data.data [43]);
tran (cddip1_im_din[76], \cddip1_im_din.data.data [44]);
tran (cddip1_im_din[77], \cddip1_im_din.data.data [45]);
tran (cddip1_im_din[78], \cddip1_im_din.data.data [46]);
tran (cddip1_im_din[79], \cddip1_im_din.data.data [47]);
tran (cddip1_im_din[80], \cddip1_im_din.data.data [48]);
tran (cddip1_im_din[81], \cddip1_im_din.data.data [49]);
tran (cddip1_im_din[82], \cddip1_im_din.data.data [50]);
tran (cddip1_im_din[83], \cddip1_im_din.data.data [51]);
tran (cddip1_im_din[84], \cddip1_im_din.data.data [52]);
tran (cddip1_im_din[85], \cddip1_im_din.data.data [53]);
tran (cddip1_im_din[86], \cddip1_im_din.data.data [54]);
tran (cddip1_im_din[87], \cddip1_im_din.data.data [55]);
tran (cddip1_im_din[88], \cddip1_im_din.data.data [56]);
tran (cddip1_im_din[89], \cddip1_im_din.data.data [57]);
tran (cddip1_im_din[90], \cddip1_im_din.data.data [58]);
tran (cddip1_im_din[91], \cddip1_im_din.data.data [59]);
tran (cddip1_im_din[92], \cddip1_im_din.data.data [60]);
tran (cddip1_im_din[93], \cddip1_im_din.data.data [61]);
tran (cddip1_im_din[94], \cddip1_im_din.data.data [62]);
tran (cddip1_im_din[95], \cddip1_im_din.data.data [63]);
tran (cceip1_im_din[6], \cceip1_im_din.desc.im_meta [6]);
tran (cceip1_im_din[8], \cceip1_im_din.desc.im_meta [8]);
tran (cceip1_im_din[9], \cceip1_im_din.desc.im_meta [9]);
tran (cceip1_im_din[10], \cceip1_im_din.desc.im_meta [10]);
tran (cceip1_im_din[11], \cceip1_im_din.desc.im_meta [11]);
tran (cceip1_im_din[12], \cceip1_im_din.desc.im_meta [12]);
tran (cceip1_im_din[13], \cceip1_im_din.desc.im_meta [13]);
tran (cceip1_im_din[14], \cceip1_im_din.desc.im_meta [14]);
tran (cceip1_im_din[23], \cceip1_im_din.desc.bytes_vld [0]);
tran (cceip1_im_din[24], \cceip1_im_din.desc.bytes_vld [1]);
tran (cceip1_im_din[25], \cceip1_im_din.desc.bytes_vld [2]);
tran (cceip1_im_din[26], \cceip1_im_din.desc.bytes_vld [3]);
tran (cceip1_im_din[27], \cceip1_im_din.desc.bytes_vld [4]);
tran (cceip1_im_din[28], \cceip1_im_din.desc.bytes_vld [5]);
tran (cceip1_im_din[29], \cceip1_im_din.desc.bytes_vld [6]);
tran (cceip1_im_din[30], \cceip1_im_din.desc.bytes_vld [7]);
tran (cceip1_im_din[31], \cceip1_im_din.desc.eob );
tran (cceip1_im_din[7], \cceip1_im_din.desc.im_meta [7]);
tran (cceip1_im_din[32], \cceip1_im_din.data.data [0]);
tran (cceip1_im_din[33], \cceip1_im_din.data.data [1]);
tran (cceip1_im_din[34], \cceip1_im_din.data.data [2]);
tran (cceip1_im_din[35], \cceip1_im_din.data.data [3]);
tran (cceip1_im_din[36], \cceip1_im_din.data.data [4]);
tran (cceip1_im_din[37], \cceip1_im_din.data.data [5]);
tran (cceip1_im_din[38], \cceip1_im_din.data.data [6]);
tran (cceip1_im_din[39], \cceip1_im_din.data.data [7]);
tran (cceip1_im_din[40], \cceip1_im_din.data.data [8]);
tran (cceip1_im_din[41], \cceip1_im_din.data.data [9]);
tran (cceip1_im_din[42], \cceip1_im_din.data.data [10]);
tran (cceip1_im_din[43], \cceip1_im_din.data.data [11]);
tran (cceip1_im_din[44], \cceip1_im_din.data.data [12]);
tran (cceip1_im_din[45], \cceip1_im_din.data.data [13]);
tran (cceip1_im_din[46], \cceip1_im_din.data.data [14]);
tran (cceip1_im_din[47], \cceip1_im_din.data.data [15]);
tran (cceip1_im_din[48], \cceip1_im_din.data.data [16]);
tran (cceip1_im_din[49], \cceip1_im_din.data.data [17]);
tran (cceip1_im_din[50], \cceip1_im_din.data.data [18]);
tran (cceip1_im_din[51], \cceip1_im_din.data.data [19]);
tran (cceip1_im_din[52], \cceip1_im_din.data.data [20]);
tran (cceip1_im_din[53], \cceip1_im_din.data.data [21]);
tran (cceip1_im_din[54], \cceip1_im_din.data.data [22]);
tran (cceip1_im_din[55], \cceip1_im_din.data.data [23]);
tran (cceip1_im_din[56], \cceip1_im_din.data.data [24]);
tran (cceip1_im_din[57], \cceip1_im_din.data.data [25]);
tran (cceip1_im_din[58], \cceip1_im_din.data.data [26]);
tran (cceip1_im_din[59], \cceip1_im_din.data.data [27]);
tran (cceip1_im_din[60], \cceip1_im_din.data.data [28]);
tran (cceip1_im_din[61], \cceip1_im_din.data.data [29]);
tran (cceip1_im_din[62], \cceip1_im_din.data.data [30]);
tran (cceip1_im_din[63], \cceip1_im_din.data.data [31]);
tran (cceip1_im_din[64], \cceip1_im_din.data.data [32]);
tran (cceip1_im_din[65], \cceip1_im_din.data.data [33]);
tran (cceip1_im_din[66], \cceip1_im_din.data.data [34]);
tran (cceip1_im_din[67], \cceip1_im_din.data.data [35]);
tran (cceip1_im_din[68], \cceip1_im_din.data.data [36]);
tran (cceip1_im_din[69], \cceip1_im_din.data.data [37]);
tran (cceip1_im_din[70], \cceip1_im_din.data.data [38]);
tran (cceip1_im_din[71], \cceip1_im_din.data.data [39]);
tran (cceip1_im_din[72], \cceip1_im_din.data.data [40]);
tran (cceip1_im_din[73], \cceip1_im_din.data.data [41]);
tran (cceip1_im_din[74], \cceip1_im_din.data.data [42]);
tran (cceip1_im_din[75], \cceip1_im_din.data.data [43]);
tran (cceip1_im_din[76], \cceip1_im_din.data.data [44]);
tran (cceip1_im_din[77], \cceip1_im_din.data.data [45]);
tran (cceip1_im_din[78], \cceip1_im_din.data.data [46]);
tran (cceip1_im_din[79], \cceip1_im_din.data.data [47]);
tran (cceip1_im_din[80], \cceip1_im_din.data.data [48]);
tran (cceip1_im_din[81], \cceip1_im_din.data.data [49]);
tran (cceip1_im_din[82], \cceip1_im_din.data.data [50]);
tran (cceip1_im_din[83], \cceip1_im_din.data.data [51]);
tran (cceip1_im_din[84], \cceip1_im_din.data.data [52]);
tran (cceip1_im_din[85], \cceip1_im_din.data.data [53]);
tran (cceip1_im_din[86], \cceip1_im_din.data.data [54]);
tran (cceip1_im_din[87], \cceip1_im_din.data.data [55]);
tran (cceip1_im_din[88], \cceip1_im_din.data.data [56]);
tran (cceip1_im_din[89], \cceip1_im_din.data.data [57]);
tran (cceip1_im_din[90], \cceip1_im_din.data.data [58]);
tran (cceip1_im_din[91], \cceip1_im_din.data.data [59]);
tran (cceip1_im_din[92], \cceip1_im_din.data.data [60]);
tran (cceip1_im_din[93], \cceip1_im_din.data.data [61]);
tran (cceip1_im_din[94], \cceip1_im_din.data.data [62]);
tran (cceip1_im_din[95], \cceip1_im_din.data.data [63]);
tran (cddip0_im_din[6], \cddip0_im_din.desc.im_meta [6]);
tran (cddip0_im_din[8], \cddip0_im_din.desc.im_meta [8]);
tran (cddip0_im_din[9], \cddip0_im_din.desc.im_meta [9]);
tran (cddip0_im_din[10], \cddip0_im_din.desc.im_meta [10]);
tran (cddip0_im_din[11], \cddip0_im_din.desc.im_meta [11]);
tran (cddip0_im_din[12], \cddip0_im_din.desc.im_meta [12]);
tran (cddip0_im_din[13], \cddip0_im_din.desc.im_meta [13]);
tran (cddip0_im_din[14], \cddip0_im_din.desc.im_meta [14]);
tran (cddip0_im_din[23], \cddip0_im_din.desc.bytes_vld [0]);
tran (cddip0_im_din[24], \cddip0_im_din.desc.bytes_vld [1]);
tran (cddip0_im_din[25], \cddip0_im_din.desc.bytes_vld [2]);
tran (cddip0_im_din[26], \cddip0_im_din.desc.bytes_vld [3]);
tran (cddip0_im_din[27], \cddip0_im_din.desc.bytes_vld [4]);
tran (cddip0_im_din[28], \cddip0_im_din.desc.bytes_vld [5]);
tran (cddip0_im_din[29], \cddip0_im_din.desc.bytes_vld [6]);
tran (cddip0_im_din[30], \cddip0_im_din.desc.bytes_vld [7]);
tran (cddip0_im_din[31], \cddip0_im_din.desc.eob );
tran (cddip0_im_din[7], \cddip0_im_din.desc.im_meta [7]);
tran (cddip0_im_din[32], \cddip0_im_din.data.data [0]);
tran (cddip0_im_din[33], \cddip0_im_din.data.data [1]);
tran (cddip0_im_din[34], \cddip0_im_din.data.data [2]);
tran (cddip0_im_din[35], \cddip0_im_din.data.data [3]);
tran (cddip0_im_din[36], \cddip0_im_din.data.data [4]);
tran (cddip0_im_din[37], \cddip0_im_din.data.data [5]);
tran (cddip0_im_din[38], \cddip0_im_din.data.data [6]);
tran (cddip0_im_din[39], \cddip0_im_din.data.data [7]);
tran (cddip0_im_din[40], \cddip0_im_din.data.data [8]);
tran (cddip0_im_din[41], \cddip0_im_din.data.data [9]);
tran (cddip0_im_din[42], \cddip0_im_din.data.data [10]);
tran (cddip0_im_din[43], \cddip0_im_din.data.data [11]);
tran (cddip0_im_din[44], \cddip0_im_din.data.data [12]);
tran (cddip0_im_din[45], \cddip0_im_din.data.data [13]);
tran (cddip0_im_din[46], \cddip0_im_din.data.data [14]);
tran (cddip0_im_din[47], \cddip0_im_din.data.data [15]);
tran (cddip0_im_din[48], \cddip0_im_din.data.data [16]);
tran (cddip0_im_din[49], \cddip0_im_din.data.data [17]);
tran (cddip0_im_din[50], \cddip0_im_din.data.data [18]);
tran (cddip0_im_din[51], \cddip0_im_din.data.data [19]);
tran (cddip0_im_din[52], \cddip0_im_din.data.data [20]);
tran (cddip0_im_din[53], \cddip0_im_din.data.data [21]);
tran (cddip0_im_din[54], \cddip0_im_din.data.data [22]);
tran (cddip0_im_din[55], \cddip0_im_din.data.data [23]);
tran (cddip0_im_din[56], \cddip0_im_din.data.data [24]);
tran (cddip0_im_din[57], \cddip0_im_din.data.data [25]);
tran (cddip0_im_din[58], \cddip0_im_din.data.data [26]);
tran (cddip0_im_din[59], \cddip0_im_din.data.data [27]);
tran (cddip0_im_din[60], \cddip0_im_din.data.data [28]);
tran (cddip0_im_din[61], \cddip0_im_din.data.data [29]);
tran (cddip0_im_din[62], \cddip0_im_din.data.data [30]);
tran (cddip0_im_din[63], \cddip0_im_din.data.data [31]);
tran (cddip0_im_din[64], \cddip0_im_din.data.data [32]);
tran (cddip0_im_din[65], \cddip0_im_din.data.data [33]);
tran (cddip0_im_din[66], \cddip0_im_din.data.data [34]);
tran (cddip0_im_din[67], \cddip0_im_din.data.data [35]);
tran (cddip0_im_din[68], \cddip0_im_din.data.data [36]);
tran (cddip0_im_din[69], \cddip0_im_din.data.data [37]);
tran (cddip0_im_din[70], \cddip0_im_din.data.data [38]);
tran (cddip0_im_din[71], \cddip0_im_din.data.data [39]);
tran (cddip0_im_din[72], \cddip0_im_din.data.data [40]);
tran (cddip0_im_din[73], \cddip0_im_din.data.data [41]);
tran (cddip0_im_din[74], \cddip0_im_din.data.data [42]);
tran (cddip0_im_din[75], \cddip0_im_din.data.data [43]);
tran (cddip0_im_din[76], \cddip0_im_din.data.data [44]);
tran (cddip0_im_din[77], \cddip0_im_din.data.data [45]);
tran (cddip0_im_din[78], \cddip0_im_din.data.data [46]);
tran (cddip0_im_din[79], \cddip0_im_din.data.data [47]);
tran (cddip0_im_din[80], \cddip0_im_din.data.data [48]);
tran (cddip0_im_din[81], \cddip0_im_din.data.data [49]);
tran (cddip0_im_din[82], \cddip0_im_din.data.data [50]);
tran (cddip0_im_din[83], \cddip0_im_din.data.data [51]);
tran (cddip0_im_din[84], \cddip0_im_din.data.data [52]);
tran (cddip0_im_din[85], \cddip0_im_din.data.data [53]);
tran (cddip0_im_din[86], \cddip0_im_din.data.data [54]);
tran (cddip0_im_din[87], \cddip0_im_din.data.data [55]);
tran (cddip0_im_din[88], \cddip0_im_din.data.data [56]);
tran (cddip0_im_din[89], \cddip0_im_din.data.data [57]);
tran (cddip0_im_din[90], \cddip0_im_din.data.data [58]);
tran (cddip0_im_din[91], \cddip0_im_din.data.data [59]);
tran (cddip0_im_din[92], \cddip0_im_din.data.data [60]);
tran (cddip0_im_din[93], \cddip0_im_din.data.data [61]);
tran (cddip0_im_din[94], \cddip0_im_din.data.data [62]);
tran (cddip0_im_din[95], \cddip0_im_din.data.data [63]);
tran (cceip0_im_din[6], \cceip0_im_din.desc.im_meta [6]);
tran (cceip0_im_din[8], \cceip0_im_din.desc.im_meta [8]);
tran (cceip0_im_din[9], \cceip0_im_din.desc.im_meta [9]);
tran (cceip0_im_din[10], \cceip0_im_din.desc.im_meta [10]);
tran (cceip0_im_din[11], \cceip0_im_din.desc.im_meta [11]);
tran (cceip0_im_din[12], \cceip0_im_din.desc.im_meta [12]);
tran (cceip0_im_din[13], \cceip0_im_din.desc.im_meta [13]);
tran (cceip0_im_din[14], \cceip0_im_din.desc.im_meta [14]);
tran (cceip0_im_din[23], \cceip0_im_din.desc.bytes_vld [0]);
tran (cceip0_im_din[24], \cceip0_im_din.desc.bytes_vld [1]);
tran (cceip0_im_din[25], \cceip0_im_din.desc.bytes_vld [2]);
tran (cceip0_im_din[26], \cceip0_im_din.desc.bytes_vld [3]);
tran (cceip0_im_din[27], \cceip0_im_din.desc.bytes_vld [4]);
tran (cceip0_im_din[28], \cceip0_im_din.desc.bytes_vld [5]);
tran (cceip0_im_din[29], \cceip0_im_din.desc.bytes_vld [6]);
tran (cceip0_im_din[30], \cceip0_im_din.desc.bytes_vld [7]);
tran (cceip0_im_din[31], \cceip0_im_din.desc.eob );
tran (cceip0_im_din[7], \cceip0_im_din.desc.im_meta [7]);
tran (cceip0_im_din[32], \cceip0_im_din.data.data [0]);
tran (cceip0_im_din[33], \cceip0_im_din.data.data [1]);
tran (cceip0_im_din[34], \cceip0_im_din.data.data [2]);
tran (cceip0_im_din[35], \cceip0_im_din.data.data [3]);
tran (cceip0_im_din[36], \cceip0_im_din.data.data [4]);
tran (cceip0_im_din[37], \cceip0_im_din.data.data [5]);
tran (cceip0_im_din[38], \cceip0_im_din.data.data [6]);
tran (cceip0_im_din[39], \cceip0_im_din.data.data [7]);
tran (cceip0_im_din[40], \cceip0_im_din.data.data [8]);
tran (cceip0_im_din[41], \cceip0_im_din.data.data [9]);
tran (cceip0_im_din[42], \cceip0_im_din.data.data [10]);
tran (cceip0_im_din[43], \cceip0_im_din.data.data [11]);
tran (cceip0_im_din[44], \cceip0_im_din.data.data [12]);
tran (cceip0_im_din[45], \cceip0_im_din.data.data [13]);
tran (cceip0_im_din[46], \cceip0_im_din.data.data [14]);
tran (cceip0_im_din[47], \cceip0_im_din.data.data [15]);
tran (cceip0_im_din[48], \cceip0_im_din.data.data [16]);
tran (cceip0_im_din[49], \cceip0_im_din.data.data [17]);
tran (cceip0_im_din[50], \cceip0_im_din.data.data [18]);
tran (cceip0_im_din[51], \cceip0_im_din.data.data [19]);
tran (cceip0_im_din[52], \cceip0_im_din.data.data [20]);
tran (cceip0_im_din[53], \cceip0_im_din.data.data [21]);
tran (cceip0_im_din[54], \cceip0_im_din.data.data [22]);
tran (cceip0_im_din[55], \cceip0_im_din.data.data [23]);
tran (cceip0_im_din[56], \cceip0_im_din.data.data [24]);
tran (cceip0_im_din[57], \cceip0_im_din.data.data [25]);
tran (cceip0_im_din[58], \cceip0_im_din.data.data [26]);
tran (cceip0_im_din[59], \cceip0_im_din.data.data [27]);
tran (cceip0_im_din[60], \cceip0_im_din.data.data [28]);
tran (cceip0_im_din[61], \cceip0_im_din.data.data [29]);
tran (cceip0_im_din[62], \cceip0_im_din.data.data [30]);
tran (cceip0_im_din[63], \cceip0_im_din.data.data [31]);
tran (cceip0_im_din[64], \cceip0_im_din.data.data [32]);
tran (cceip0_im_din[65], \cceip0_im_din.data.data [33]);
tran (cceip0_im_din[66], \cceip0_im_din.data.data [34]);
tran (cceip0_im_din[67], \cceip0_im_din.data.data [35]);
tran (cceip0_im_din[68], \cceip0_im_din.data.data [36]);
tran (cceip0_im_din[69], \cceip0_im_din.data.data [37]);
tran (cceip0_im_din[70], \cceip0_im_din.data.data [38]);
tran (cceip0_im_din[71], \cceip0_im_din.data.data [39]);
tran (cceip0_im_din[72], \cceip0_im_din.data.data [40]);
tran (cceip0_im_din[73], \cceip0_im_din.data.data [41]);
tran (cceip0_im_din[74], \cceip0_im_din.data.data [42]);
tran (cceip0_im_din[75], \cceip0_im_din.data.data [43]);
tran (cceip0_im_din[76], \cceip0_im_din.data.data [44]);
tran (cceip0_im_din[77], \cceip0_im_din.data.data [45]);
tran (cceip0_im_din[78], \cceip0_im_din.data.data [46]);
tran (cceip0_im_din[79], \cceip0_im_din.data.data [47]);
tran (cceip0_im_din[80], \cceip0_im_din.data.data [48]);
tran (cceip0_im_din[81], \cceip0_im_din.data.data [49]);
tran (cceip0_im_din[82], \cceip0_im_din.data.data [50]);
tran (cceip0_im_din[83], \cceip0_im_din.data.data [51]);
tran (cceip0_im_din[84], \cceip0_im_din.data.data [52]);
tran (cceip0_im_din[85], \cceip0_im_din.data.data [53]);
tran (cceip0_im_din[86], \cceip0_im_din.data.data [54]);
tran (cceip0_im_din[87], \cceip0_im_din.data.data [55]);
tran (cceip0_im_din[88], \cceip0_im_din.data.data [56]);
tran (cceip0_im_din[89], \cceip0_im_din.data.data [57]);
tran (cceip0_im_din[90], \cceip0_im_din.data.data [58]);
tran (cceip0_im_din[91], \cceip0_im_din.data.data [59]);
tran (cceip0_im_din[92], \cceip0_im_din.data.data [60]);
tran (cceip0_im_din[93], \cceip0_im_din.data.data [61]);
tran (cceip0_im_din[94], \cceip0_im_din.data.data [62]);
tran (cceip0_im_din[95], \cceip0_im_din.data.data [63]);
tran (spare[31], \spare.r.part0 [31]);
tran (spare[31], \spare.f.spare [31]);
tran (spare[30], \spare.r.part0 [30]);
tran (spare[30], \spare.f.spare [30]);
tran (spare[29], \spare.r.part0 [29]);
tran (spare[29], \spare.f.spare [29]);
tran (spare[28], \spare.r.part0 [28]);
tran (spare[28], \spare.f.spare [28]);
tran (spare[27], \spare.r.part0 [27]);
tran (spare[27], \spare.f.spare [27]);
tran (spare[26], \spare.r.part0 [26]);
tran (spare[26], \spare.f.spare [26]);
tran (spare[25], \spare.r.part0 [25]);
tran (spare[25], \spare.f.spare [25]);
tran (spare[24], \spare.r.part0 [24]);
tran (spare[24], \spare.f.spare [24]);
tran (spare[23], \spare.r.part0 [23]);
tran (spare[23], \spare.f.spare [23]);
tran (spare[22], \spare.r.part0 [22]);
tran (spare[22], \spare.f.spare [22]);
tran (spare[21], \spare.r.part0 [21]);
tran (spare[21], \spare.f.spare [21]);
tran (spare[20], \spare.r.part0 [20]);
tran (spare[20], \spare.f.spare [20]);
tran (spare[19], \spare.r.part0 [19]);
tran (spare[19], \spare.f.spare [19]);
tran (spare[18], \spare.r.part0 [18]);
tran (spare[18], \spare.f.spare [18]);
tran (spare[17], \spare.r.part0 [17]);
tran (spare[17], \spare.f.spare [17]);
tran (spare[16], \spare.r.part0 [16]);
tran (spare[16], \spare.f.spare [16]);
tran (spare[15], \spare.r.part0 [15]);
tran (spare[15], \spare.f.spare [15]);
tran (spare[14], \spare.r.part0 [14]);
tran (spare[14], \spare.f.spare [14]);
tran (spare[13], \spare.r.part0 [13]);
tran (spare[13], \spare.f.spare [13]);
tran (spare[12], \spare.r.part0 [12]);
tran (spare[12], \spare.f.spare [12]);
tran (spare[11], \spare.r.part0 [11]);
tran (spare[11], \spare.f.spare [11]);
tran (spare[10], \spare.r.part0 [10]);
tran (spare[10], \spare.f.spare [10]);
tran (spare[9], \spare.r.part0 [9]);
tran (spare[9], \spare.f.spare [9]);
tran (spare[8], \spare.r.part0 [8]);
tran (spare[8], \spare.f.spare [8]);
tran (spare[7], \spare.r.part0 [7]);
tran (spare[7], \spare.f.spare [7]);
tran (spare[3], \spare.r.part0 [3]);
tran (spare[3], \spare.f.spare [3]);
tran (cceip0_out_ia_wdata[31], \cceip0_out_ia_wdata.r.part0 [31]);
tran (cceip0_out_ia_wdata[31], \cceip0_out_ia_wdata.f.eob );
tran (cceip0_out_ia_wdata[30], \cceip0_out_ia_wdata.r.part0 [30]);
tran (cceip0_out_ia_wdata[30], \cceip0_out_ia_wdata.f.bytes_vld [7]);
tran (cceip0_out_ia_wdata[29], \cceip0_out_ia_wdata.r.part0 [29]);
tran (cceip0_out_ia_wdata[29], \cceip0_out_ia_wdata.f.bytes_vld [6]);
tran (cceip0_out_ia_wdata[28], \cceip0_out_ia_wdata.r.part0 [28]);
tran (cceip0_out_ia_wdata[28], \cceip0_out_ia_wdata.f.bytes_vld [5]);
tran (cceip0_out_ia_wdata[27], \cceip0_out_ia_wdata.r.part0 [27]);
tran (cceip0_out_ia_wdata[27], \cceip0_out_ia_wdata.f.bytes_vld [4]);
tran (cceip0_out_ia_wdata[26], \cceip0_out_ia_wdata.r.part0 [26]);
tran (cceip0_out_ia_wdata[26], \cceip0_out_ia_wdata.f.bytes_vld [3]);
tran (cceip0_out_ia_wdata[25], \cceip0_out_ia_wdata.r.part0 [25]);
tran (cceip0_out_ia_wdata[25], \cceip0_out_ia_wdata.f.bytes_vld [2]);
tran (cceip0_out_ia_wdata[24], \cceip0_out_ia_wdata.r.part0 [24]);
tran (cceip0_out_ia_wdata[24], \cceip0_out_ia_wdata.f.bytes_vld [1]);
tran (cceip0_out_ia_wdata[23], \cceip0_out_ia_wdata.r.part0 [23]);
tran (cceip0_out_ia_wdata[23], \cceip0_out_ia_wdata.f.bytes_vld [0]);
tran (cceip0_out_ia_wdata[22], \cceip0_out_ia_wdata.r.part0 [22]);
tran (cceip0_out_ia_wdata[22], \cceip0_out_ia_wdata.f.unused1 [7]);
tran (cceip0_out_ia_wdata[21], \cceip0_out_ia_wdata.r.part0 [21]);
tran (cceip0_out_ia_wdata[21], \cceip0_out_ia_wdata.f.unused1 [6]);
tran (cceip0_out_ia_wdata[20], \cceip0_out_ia_wdata.r.part0 [20]);
tran (cceip0_out_ia_wdata[20], \cceip0_out_ia_wdata.f.unused1 [5]);
tran (cceip0_out_ia_wdata[19], \cceip0_out_ia_wdata.r.part0 [19]);
tran (cceip0_out_ia_wdata[19], \cceip0_out_ia_wdata.f.unused1 [4]);
tran (cceip0_out_ia_wdata[18], \cceip0_out_ia_wdata.r.part0 [18]);
tran (cceip0_out_ia_wdata[18], \cceip0_out_ia_wdata.f.unused1 [3]);
tran (cceip0_out_ia_wdata[17], \cceip0_out_ia_wdata.r.part0 [17]);
tran (cceip0_out_ia_wdata[17], \cceip0_out_ia_wdata.f.unused1 [2]);
tran (cceip0_out_ia_wdata[16], \cceip0_out_ia_wdata.r.part0 [16]);
tran (cceip0_out_ia_wdata[16], \cceip0_out_ia_wdata.f.unused1 [1]);
tran (cceip0_out_ia_wdata[15], \cceip0_out_ia_wdata.r.part0 [15]);
tran (cceip0_out_ia_wdata[15], \cceip0_out_ia_wdata.f.unused1 [0]);
tran (cceip0_out_ia_wdata[14], \cceip0_out_ia_wdata.r.part0 [14]);
tran (cceip0_out_ia_wdata[14], \cceip0_out_ia_wdata.f.tid );
tran (cceip0_out_ia_wdata[13], \cceip0_out_ia_wdata.r.part0 [13]);
tran (cceip0_out_ia_wdata[13], \cceip0_out_ia_wdata.f.tuser [7]);
tran (cceip0_out_ia_wdata[12], \cceip0_out_ia_wdata.r.part0 [12]);
tran (cceip0_out_ia_wdata[12], \cceip0_out_ia_wdata.f.tuser [6]);
tran (cceip0_out_ia_wdata[11], \cceip0_out_ia_wdata.r.part0 [11]);
tran (cceip0_out_ia_wdata[11], \cceip0_out_ia_wdata.f.tuser [5]);
tran (cceip0_out_ia_wdata[10], \cceip0_out_ia_wdata.r.part0 [10]);
tran (cceip0_out_ia_wdata[10], \cceip0_out_ia_wdata.f.tuser [4]);
tran (cceip0_out_ia_wdata[9], \cceip0_out_ia_wdata.r.part0 [9]);
tran (cceip0_out_ia_wdata[9], \cceip0_out_ia_wdata.f.tuser [3]);
tran (cceip0_out_ia_wdata[8], \cceip0_out_ia_wdata.r.part0 [8]);
tran (cceip0_out_ia_wdata[8], \cceip0_out_ia_wdata.f.tuser [2]);
tran (cceip0_out_ia_wdata[7], \cceip0_out_ia_wdata.r.part0 [7]);
tran (cceip0_out_ia_wdata[7], \cceip0_out_ia_wdata.f.tuser [1]);
tran (cceip0_out_ia_wdata[6], \cceip0_out_ia_wdata.r.part0 [6]);
tran (cceip0_out_ia_wdata[6], \cceip0_out_ia_wdata.f.tuser [0]);
tran (cceip0_out_ia_wdata[5], \cceip0_out_ia_wdata.r.part0 [5]);
tran (cceip0_out_ia_wdata[5], \cceip0_out_ia_wdata.f.unused0 [5]);
tran (cceip0_out_ia_wdata[4], \cceip0_out_ia_wdata.r.part0 [4]);
tran (cceip0_out_ia_wdata[4], \cceip0_out_ia_wdata.f.unused0 [4]);
tran (cceip0_out_ia_wdata[3], \cceip0_out_ia_wdata.r.part0 [3]);
tran (cceip0_out_ia_wdata[3], \cceip0_out_ia_wdata.f.unused0 [3]);
tran (cceip0_out_ia_wdata[2], \cceip0_out_ia_wdata.r.part0 [2]);
tran (cceip0_out_ia_wdata[2], \cceip0_out_ia_wdata.f.unused0 [2]);
tran (cceip0_out_ia_wdata[1], \cceip0_out_ia_wdata.r.part0 [1]);
tran (cceip0_out_ia_wdata[1], \cceip0_out_ia_wdata.f.unused0 [1]);
tran (cceip0_out_ia_wdata[0], \cceip0_out_ia_wdata.r.part0 [0]);
tran (cceip0_out_ia_wdata[0], \cceip0_out_ia_wdata.f.unused0 [0]);
tran (cceip0_out_ia_wdata[63], \cceip0_out_ia_wdata.r.part1 [31]);
tran (cceip0_out_ia_wdata[63], \cceip0_out_ia_wdata.f.tdata_lo [31]);
tran (cceip0_out_ia_wdata[62], \cceip0_out_ia_wdata.r.part1 [30]);
tran (cceip0_out_ia_wdata[62], \cceip0_out_ia_wdata.f.tdata_lo [30]);
tran (cceip0_out_ia_wdata[61], \cceip0_out_ia_wdata.r.part1 [29]);
tran (cceip0_out_ia_wdata[61], \cceip0_out_ia_wdata.f.tdata_lo [29]);
tran (cceip0_out_ia_wdata[60], \cceip0_out_ia_wdata.r.part1 [28]);
tran (cceip0_out_ia_wdata[60], \cceip0_out_ia_wdata.f.tdata_lo [28]);
tran (cceip0_out_ia_wdata[59], \cceip0_out_ia_wdata.r.part1 [27]);
tran (cceip0_out_ia_wdata[59], \cceip0_out_ia_wdata.f.tdata_lo [27]);
tran (cceip0_out_ia_wdata[58], \cceip0_out_ia_wdata.r.part1 [26]);
tran (cceip0_out_ia_wdata[58], \cceip0_out_ia_wdata.f.tdata_lo [26]);
tran (cceip0_out_ia_wdata[57], \cceip0_out_ia_wdata.r.part1 [25]);
tran (cceip0_out_ia_wdata[57], \cceip0_out_ia_wdata.f.tdata_lo [25]);
tran (cceip0_out_ia_wdata[56], \cceip0_out_ia_wdata.r.part1 [24]);
tran (cceip0_out_ia_wdata[56], \cceip0_out_ia_wdata.f.tdata_lo [24]);
tran (cceip0_out_ia_wdata[55], \cceip0_out_ia_wdata.r.part1 [23]);
tran (cceip0_out_ia_wdata[55], \cceip0_out_ia_wdata.f.tdata_lo [23]);
tran (cceip0_out_ia_wdata[54], \cceip0_out_ia_wdata.r.part1 [22]);
tran (cceip0_out_ia_wdata[54], \cceip0_out_ia_wdata.f.tdata_lo [22]);
tran (cceip0_out_ia_wdata[53], \cceip0_out_ia_wdata.r.part1 [21]);
tran (cceip0_out_ia_wdata[53], \cceip0_out_ia_wdata.f.tdata_lo [21]);
tran (cceip0_out_ia_wdata[52], \cceip0_out_ia_wdata.r.part1 [20]);
tran (cceip0_out_ia_wdata[52], \cceip0_out_ia_wdata.f.tdata_lo [20]);
tran (cceip0_out_ia_wdata[51], \cceip0_out_ia_wdata.r.part1 [19]);
tran (cceip0_out_ia_wdata[51], \cceip0_out_ia_wdata.f.tdata_lo [19]);
tran (cceip0_out_ia_wdata[50], \cceip0_out_ia_wdata.r.part1 [18]);
tran (cceip0_out_ia_wdata[50], \cceip0_out_ia_wdata.f.tdata_lo [18]);
tran (cceip0_out_ia_wdata[49], \cceip0_out_ia_wdata.r.part1 [17]);
tran (cceip0_out_ia_wdata[49], \cceip0_out_ia_wdata.f.tdata_lo [17]);
tran (cceip0_out_ia_wdata[48], \cceip0_out_ia_wdata.r.part1 [16]);
tran (cceip0_out_ia_wdata[48], \cceip0_out_ia_wdata.f.tdata_lo [16]);
tran (cceip0_out_ia_wdata[47], \cceip0_out_ia_wdata.r.part1 [15]);
tran (cceip0_out_ia_wdata[47], \cceip0_out_ia_wdata.f.tdata_lo [15]);
tran (cceip0_out_ia_wdata[46], \cceip0_out_ia_wdata.r.part1 [14]);
tran (cceip0_out_ia_wdata[46], \cceip0_out_ia_wdata.f.tdata_lo [14]);
tran (cceip0_out_ia_wdata[45], \cceip0_out_ia_wdata.r.part1 [13]);
tran (cceip0_out_ia_wdata[45], \cceip0_out_ia_wdata.f.tdata_lo [13]);
tran (cceip0_out_ia_wdata[44], \cceip0_out_ia_wdata.r.part1 [12]);
tran (cceip0_out_ia_wdata[44], \cceip0_out_ia_wdata.f.tdata_lo [12]);
tran (cceip0_out_ia_wdata[43], \cceip0_out_ia_wdata.r.part1 [11]);
tran (cceip0_out_ia_wdata[43], \cceip0_out_ia_wdata.f.tdata_lo [11]);
tran (cceip0_out_ia_wdata[42], \cceip0_out_ia_wdata.r.part1 [10]);
tran (cceip0_out_ia_wdata[42], \cceip0_out_ia_wdata.f.tdata_lo [10]);
tran (cceip0_out_ia_wdata[41], \cceip0_out_ia_wdata.r.part1 [9]);
tran (cceip0_out_ia_wdata[41], \cceip0_out_ia_wdata.f.tdata_lo [9]);
tran (cceip0_out_ia_wdata[40], \cceip0_out_ia_wdata.r.part1 [8]);
tran (cceip0_out_ia_wdata[40], \cceip0_out_ia_wdata.f.tdata_lo [8]);
tran (cceip0_out_ia_wdata[39], \cceip0_out_ia_wdata.r.part1 [7]);
tran (cceip0_out_ia_wdata[39], \cceip0_out_ia_wdata.f.tdata_lo [7]);
tran (cceip0_out_ia_wdata[38], \cceip0_out_ia_wdata.r.part1 [6]);
tran (cceip0_out_ia_wdata[38], \cceip0_out_ia_wdata.f.tdata_lo [6]);
tran (cceip0_out_ia_wdata[37], \cceip0_out_ia_wdata.r.part1 [5]);
tran (cceip0_out_ia_wdata[37], \cceip0_out_ia_wdata.f.tdata_lo [5]);
tran (cceip0_out_ia_wdata[36], \cceip0_out_ia_wdata.r.part1 [4]);
tran (cceip0_out_ia_wdata[36], \cceip0_out_ia_wdata.f.tdata_lo [4]);
tran (cceip0_out_ia_wdata[35], \cceip0_out_ia_wdata.r.part1 [3]);
tran (cceip0_out_ia_wdata[35], \cceip0_out_ia_wdata.f.tdata_lo [3]);
tran (cceip0_out_ia_wdata[34], \cceip0_out_ia_wdata.r.part1 [2]);
tran (cceip0_out_ia_wdata[34], \cceip0_out_ia_wdata.f.tdata_lo [2]);
tran (cceip0_out_ia_wdata[33], \cceip0_out_ia_wdata.r.part1 [1]);
tran (cceip0_out_ia_wdata[33], \cceip0_out_ia_wdata.f.tdata_lo [1]);
tran (cceip0_out_ia_wdata[32], \cceip0_out_ia_wdata.r.part1 [0]);
tran (cceip0_out_ia_wdata[32], \cceip0_out_ia_wdata.f.tdata_lo [0]);
tran (cceip0_out_ia_wdata[95], \cceip0_out_ia_wdata.r.part2 [31]);
tran (cceip0_out_ia_wdata[95], \cceip0_out_ia_wdata.f.tdata_hi [31]);
tran (cceip0_out_ia_wdata[94], \cceip0_out_ia_wdata.r.part2 [30]);
tran (cceip0_out_ia_wdata[94], \cceip0_out_ia_wdata.f.tdata_hi [30]);
tran (cceip0_out_ia_wdata[93], \cceip0_out_ia_wdata.r.part2 [29]);
tran (cceip0_out_ia_wdata[93], \cceip0_out_ia_wdata.f.tdata_hi [29]);
tran (cceip0_out_ia_wdata[92], \cceip0_out_ia_wdata.r.part2 [28]);
tran (cceip0_out_ia_wdata[92], \cceip0_out_ia_wdata.f.tdata_hi [28]);
tran (cceip0_out_ia_wdata[91], \cceip0_out_ia_wdata.r.part2 [27]);
tran (cceip0_out_ia_wdata[91], \cceip0_out_ia_wdata.f.tdata_hi [27]);
tran (cceip0_out_ia_wdata[90], \cceip0_out_ia_wdata.r.part2 [26]);
tran (cceip0_out_ia_wdata[90], \cceip0_out_ia_wdata.f.tdata_hi [26]);
tran (cceip0_out_ia_wdata[89], \cceip0_out_ia_wdata.r.part2 [25]);
tran (cceip0_out_ia_wdata[89], \cceip0_out_ia_wdata.f.tdata_hi [25]);
tran (cceip0_out_ia_wdata[88], \cceip0_out_ia_wdata.r.part2 [24]);
tran (cceip0_out_ia_wdata[88], \cceip0_out_ia_wdata.f.tdata_hi [24]);
tran (cceip0_out_ia_wdata[87], \cceip0_out_ia_wdata.r.part2 [23]);
tran (cceip0_out_ia_wdata[87], \cceip0_out_ia_wdata.f.tdata_hi [23]);
tran (cceip0_out_ia_wdata[86], \cceip0_out_ia_wdata.r.part2 [22]);
tran (cceip0_out_ia_wdata[86], \cceip0_out_ia_wdata.f.tdata_hi [22]);
tran (cceip0_out_ia_wdata[85], \cceip0_out_ia_wdata.r.part2 [21]);
tran (cceip0_out_ia_wdata[85], \cceip0_out_ia_wdata.f.tdata_hi [21]);
tran (cceip0_out_ia_wdata[84], \cceip0_out_ia_wdata.r.part2 [20]);
tran (cceip0_out_ia_wdata[84], \cceip0_out_ia_wdata.f.tdata_hi [20]);
tran (cceip0_out_ia_wdata[83], \cceip0_out_ia_wdata.r.part2 [19]);
tran (cceip0_out_ia_wdata[83], \cceip0_out_ia_wdata.f.tdata_hi [19]);
tran (cceip0_out_ia_wdata[82], \cceip0_out_ia_wdata.r.part2 [18]);
tran (cceip0_out_ia_wdata[82], \cceip0_out_ia_wdata.f.tdata_hi [18]);
tran (cceip0_out_ia_wdata[81], \cceip0_out_ia_wdata.r.part2 [17]);
tran (cceip0_out_ia_wdata[81], \cceip0_out_ia_wdata.f.tdata_hi [17]);
tran (cceip0_out_ia_wdata[80], \cceip0_out_ia_wdata.r.part2 [16]);
tran (cceip0_out_ia_wdata[80], \cceip0_out_ia_wdata.f.tdata_hi [16]);
tran (cceip0_out_ia_wdata[79], \cceip0_out_ia_wdata.r.part2 [15]);
tran (cceip0_out_ia_wdata[79], \cceip0_out_ia_wdata.f.tdata_hi [15]);
tran (cceip0_out_ia_wdata[78], \cceip0_out_ia_wdata.r.part2 [14]);
tran (cceip0_out_ia_wdata[78], \cceip0_out_ia_wdata.f.tdata_hi [14]);
tran (cceip0_out_ia_wdata[77], \cceip0_out_ia_wdata.r.part2 [13]);
tran (cceip0_out_ia_wdata[77], \cceip0_out_ia_wdata.f.tdata_hi [13]);
tran (cceip0_out_ia_wdata[76], \cceip0_out_ia_wdata.r.part2 [12]);
tran (cceip0_out_ia_wdata[76], \cceip0_out_ia_wdata.f.tdata_hi [12]);
tran (cceip0_out_ia_wdata[75], \cceip0_out_ia_wdata.r.part2 [11]);
tran (cceip0_out_ia_wdata[75], \cceip0_out_ia_wdata.f.tdata_hi [11]);
tran (cceip0_out_ia_wdata[74], \cceip0_out_ia_wdata.r.part2 [10]);
tran (cceip0_out_ia_wdata[74], \cceip0_out_ia_wdata.f.tdata_hi [10]);
tran (cceip0_out_ia_wdata[73], \cceip0_out_ia_wdata.r.part2 [9]);
tran (cceip0_out_ia_wdata[73], \cceip0_out_ia_wdata.f.tdata_hi [9]);
tran (cceip0_out_ia_wdata[72], \cceip0_out_ia_wdata.r.part2 [8]);
tran (cceip0_out_ia_wdata[72], \cceip0_out_ia_wdata.f.tdata_hi [8]);
tran (cceip0_out_ia_wdata[71], \cceip0_out_ia_wdata.r.part2 [7]);
tran (cceip0_out_ia_wdata[71], \cceip0_out_ia_wdata.f.tdata_hi [7]);
tran (cceip0_out_ia_wdata[70], \cceip0_out_ia_wdata.r.part2 [6]);
tran (cceip0_out_ia_wdata[70], \cceip0_out_ia_wdata.f.tdata_hi [6]);
tran (cceip0_out_ia_wdata[69], \cceip0_out_ia_wdata.r.part2 [5]);
tran (cceip0_out_ia_wdata[69], \cceip0_out_ia_wdata.f.tdata_hi [5]);
tran (cceip0_out_ia_wdata[68], \cceip0_out_ia_wdata.r.part2 [4]);
tran (cceip0_out_ia_wdata[68], \cceip0_out_ia_wdata.f.tdata_hi [4]);
tran (cceip0_out_ia_wdata[67], \cceip0_out_ia_wdata.r.part2 [3]);
tran (cceip0_out_ia_wdata[67], \cceip0_out_ia_wdata.f.tdata_hi [3]);
tran (cceip0_out_ia_wdata[66], \cceip0_out_ia_wdata.r.part2 [2]);
tran (cceip0_out_ia_wdata[66], \cceip0_out_ia_wdata.f.tdata_hi [2]);
tran (cceip0_out_ia_wdata[65], \cceip0_out_ia_wdata.r.part2 [1]);
tran (cceip0_out_ia_wdata[65], \cceip0_out_ia_wdata.f.tdata_hi [1]);
tran (cceip0_out_ia_wdata[64], \cceip0_out_ia_wdata.r.part2 [0]);
tran (cceip0_out_ia_wdata[64], \cceip0_out_ia_wdata.f.tdata_hi [0]);
tran (cceip0_out_ia_config[12], \cceip0_out_ia_config.r.part0 [12]);
tran (cceip0_out_ia_config[12], \cceip0_out_ia_config.f.op [3]);
tran (cceip0_out_ia_config[11], \cceip0_out_ia_config.r.part0 [11]);
tran (cceip0_out_ia_config[11], \cceip0_out_ia_config.f.op [2]);
tran (cceip0_out_ia_config[10], \cceip0_out_ia_config.r.part0 [10]);
tran (cceip0_out_ia_config[10], \cceip0_out_ia_config.f.op [1]);
tran (cceip0_out_ia_config[9], \cceip0_out_ia_config.r.part0 [9]);
tran (cceip0_out_ia_config[9], \cceip0_out_ia_config.f.op [0]);
tran (cceip0_out_ia_config[8], \cceip0_out_ia_config.r.part0 [8]);
tran (cceip0_out_ia_config[8], \cceip0_out_ia_config.f.addr [8]);
tran (cceip0_out_ia_config[7], \cceip0_out_ia_config.r.part0 [7]);
tran (cceip0_out_ia_config[7], \cceip0_out_ia_config.f.addr [7]);
tran (cceip0_out_ia_config[6], \cceip0_out_ia_config.r.part0 [6]);
tran (cceip0_out_ia_config[6], \cceip0_out_ia_config.f.addr [6]);
tran (cceip0_out_ia_config[5], \cceip0_out_ia_config.r.part0 [5]);
tran (cceip0_out_ia_config[5], \cceip0_out_ia_config.f.addr [5]);
tran (cceip0_out_ia_config[4], \cceip0_out_ia_config.r.part0 [4]);
tran (cceip0_out_ia_config[4], \cceip0_out_ia_config.f.addr [4]);
tran (cceip0_out_ia_config[3], \cceip0_out_ia_config.r.part0 [3]);
tran (cceip0_out_ia_config[3], \cceip0_out_ia_config.f.addr [3]);
tran (cceip0_out_ia_config[2], \cceip0_out_ia_config.r.part0 [2]);
tran (cceip0_out_ia_config[2], \cceip0_out_ia_config.f.addr [2]);
tran (cceip0_out_ia_config[1], \cceip0_out_ia_config.r.part0 [1]);
tran (cceip0_out_ia_config[1], \cceip0_out_ia_config.f.addr [1]);
tran (cceip0_out_ia_config[0], \cceip0_out_ia_config.r.part0 [0]);
tran (cceip0_out_ia_config[0], \cceip0_out_ia_config.f.addr [0]);
tran (cceip0_out_im_config[11], \cceip0_out_im_config.r.part0 [11]);
tran (cceip0_out_im_config[11], \cceip0_out_im_config.f.mode [1]);
tran (cceip0_out_im_config[10], \cceip0_out_im_config.r.part0 [10]);
tran (cceip0_out_im_config[10], \cceip0_out_im_config.f.mode [0]);
tran (cceip0_out_im_config[9], \cceip0_out_im_config.r.part0 [9]);
tran (cceip0_out_im_config[9], \cceip0_out_im_config.f.wr_credit_config [9]);
tran (cceip0_out_im_config[8], \cceip0_out_im_config.r.part0 [8]);
tran (cceip0_out_im_config[8], \cceip0_out_im_config.f.wr_credit_config [8]);
tran (cceip0_out_im_config[7], \cceip0_out_im_config.r.part0 [7]);
tran (cceip0_out_im_config[7], \cceip0_out_im_config.f.wr_credit_config [7]);
tran (cceip0_out_im_config[6], \cceip0_out_im_config.r.part0 [6]);
tran (cceip0_out_im_config[6], \cceip0_out_im_config.f.wr_credit_config [6]);
tran (cceip0_out_im_config[5], \cceip0_out_im_config.r.part0 [5]);
tran (cceip0_out_im_config[5], \cceip0_out_im_config.f.wr_credit_config [5]);
tran (cceip0_out_im_config[4], \cceip0_out_im_config.r.part0 [4]);
tran (cceip0_out_im_config[4], \cceip0_out_im_config.f.wr_credit_config [4]);
tran (cceip0_out_im_config[3], \cceip0_out_im_config.r.part0 [3]);
tran (cceip0_out_im_config[3], \cceip0_out_im_config.f.wr_credit_config [3]);
tran (cceip0_out_im_config[2], \cceip0_out_im_config.r.part0 [2]);
tran (cceip0_out_im_config[2], \cceip0_out_im_config.f.wr_credit_config [2]);
tran (cceip0_out_im_config[1], \cceip0_out_im_config.r.part0 [1]);
tran (cceip0_out_im_config[1], \cceip0_out_im_config.f.wr_credit_config [1]);
tran (cceip0_out_im_config[0], \cceip0_out_im_config.r.part0 [0]);
tran (cceip0_out_im_config[0], \cceip0_out_im_config.f.wr_credit_config [0]);
tran (cceip1_out_ia_wdata[31], \cceip1_out_ia_wdata.r.part0 [31]);
tran (cceip1_out_ia_wdata[31], \cceip1_out_ia_wdata.f.eob );
tran (cceip1_out_ia_wdata[30], \cceip1_out_ia_wdata.r.part0 [30]);
tran (cceip1_out_ia_wdata[30], \cceip1_out_ia_wdata.f.bytes_vld [7]);
tran (cceip1_out_ia_wdata[29], \cceip1_out_ia_wdata.r.part0 [29]);
tran (cceip1_out_ia_wdata[29], \cceip1_out_ia_wdata.f.bytes_vld [6]);
tran (cceip1_out_ia_wdata[28], \cceip1_out_ia_wdata.r.part0 [28]);
tran (cceip1_out_ia_wdata[28], \cceip1_out_ia_wdata.f.bytes_vld [5]);
tran (cceip1_out_ia_wdata[27], \cceip1_out_ia_wdata.r.part0 [27]);
tran (cceip1_out_ia_wdata[27], \cceip1_out_ia_wdata.f.bytes_vld [4]);
tran (cceip1_out_ia_wdata[26], \cceip1_out_ia_wdata.r.part0 [26]);
tran (cceip1_out_ia_wdata[26], \cceip1_out_ia_wdata.f.bytes_vld [3]);
tran (cceip1_out_ia_wdata[25], \cceip1_out_ia_wdata.r.part0 [25]);
tran (cceip1_out_ia_wdata[25], \cceip1_out_ia_wdata.f.bytes_vld [2]);
tran (cceip1_out_ia_wdata[24], \cceip1_out_ia_wdata.r.part0 [24]);
tran (cceip1_out_ia_wdata[24], \cceip1_out_ia_wdata.f.bytes_vld [1]);
tran (cceip1_out_ia_wdata[23], \cceip1_out_ia_wdata.r.part0 [23]);
tran (cceip1_out_ia_wdata[23], \cceip1_out_ia_wdata.f.bytes_vld [0]);
tran (cceip1_out_ia_wdata[22], \cceip1_out_ia_wdata.r.part0 [22]);
tran (cceip1_out_ia_wdata[22], \cceip1_out_ia_wdata.f.unused1 [7]);
tran (cceip1_out_ia_wdata[21], \cceip1_out_ia_wdata.r.part0 [21]);
tran (cceip1_out_ia_wdata[21], \cceip1_out_ia_wdata.f.unused1 [6]);
tran (cceip1_out_ia_wdata[20], \cceip1_out_ia_wdata.r.part0 [20]);
tran (cceip1_out_ia_wdata[20], \cceip1_out_ia_wdata.f.unused1 [5]);
tran (cceip1_out_ia_wdata[19], \cceip1_out_ia_wdata.r.part0 [19]);
tran (cceip1_out_ia_wdata[19], \cceip1_out_ia_wdata.f.unused1 [4]);
tran (cceip1_out_ia_wdata[18], \cceip1_out_ia_wdata.r.part0 [18]);
tran (cceip1_out_ia_wdata[18], \cceip1_out_ia_wdata.f.unused1 [3]);
tran (cceip1_out_ia_wdata[17], \cceip1_out_ia_wdata.r.part0 [17]);
tran (cceip1_out_ia_wdata[17], \cceip1_out_ia_wdata.f.unused1 [2]);
tran (cceip1_out_ia_wdata[16], \cceip1_out_ia_wdata.r.part0 [16]);
tran (cceip1_out_ia_wdata[16], \cceip1_out_ia_wdata.f.unused1 [1]);
tran (cceip1_out_ia_wdata[15], \cceip1_out_ia_wdata.r.part0 [15]);
tran (cceip1_out_ia_wdata[15], \cceip1_out_ia_wdata.f.unused1 [0]);
tran (cceip1_out_ia_wdata[14], \cceip1_out_ia_wdata.r.part0 [14]);
tran (cceip1_out_ia_wdata[14], \cceip1_out_ia_wdata.f.tid );
tran (cceip1_out_ia_wdata[13], \cceip1_out_ia_wdata.r.part0 [13]);
tran (cceip1_out_ia_wdata[13], \cceip1_out_ia_wdata.f.tuser [7]);
tran (cceip1_out_ia_wdata[12], \cceip1_out_ia_wdata.r.part0 [12]);
tran (cceip1_out_ia_wdata[12], \cceip1_out_ia_wdata.f.tuser [6]);
tran (cceip1_out_ia_wdata[11], \cceip1_out_ia_wdata.r.part0 [11]);
tran (cceip1_out_ia_wdata[11], \cceip1_out_ia_wdata.f.tuser [5]);
tran (cceip1_out_ia_wdata[10], \cceip1_out_ia_wdata.r.part0 [10]);
tran (cceip1_out_ia_wdata[10], \cceip1_out_ia_wdata.f.tuser [4]);
tran (cceip1_out_ia_wdata[9], \cceip1_out_ia_wdata.r.part0 [9]);
tran (cceip1_out_ia_wdata[9], \cceip1_out_ia_wdata.f.tuser [3]);
tran (cceip1_out_ia_wdata[8], \cceip1_out_ia_wdata.r.part0 [8]);
tran (cceip1_out_ia_wdata[8], \cceip1_out_ia_wdata.f.tuser [2]);
tran (cceip1_out_ia_wdata[7], \cceip1_out_ia_wdata.r.part0 [7]);
tran (cceip1_out_ia_wdata[7], \cceip1_out_ia_wdata.f.tuser [1]);
tran (cceip1_out_ia_wdata[6], \cceip1_out_ia_wdata.r.part0 [6]);
tran (cceip1_out_ia_wdata[6], \cceip1_out_ia_wdata.f.tuser [0]);
tran (cceip1_out_ia_wdata[5], \cceip1_out_ia_wdata.r.part0 [5]);
tran (cceip1_out_ia_wdata[5], \cceip1_out_ia_wdata.f.unused0 [5]);
tran (cceip1_out_ia_wdata[4], \cceip1_out_ia_wdata.r.part0 [4]);
tran (cceip1_out_ia_wdata[4], \cceip1_out_ia_wdata.f.unused0 [4]);
tran (cceip1_out_ia_wdata[3], \cceip1_out_ia_wdata.r.part0 [3]);
tran (cceip1_out_ia_wdata[3], \cceip1_out_ia_wdata.f.unused0 [3]);
tran (cceip1_out_ia_wdata[2], \cceip1_out_ia_wdata.r.part0 [2]);
tran (cceip1_out_ia_wdata[2], \cceip1_out_ia_wdata.f.unused0 [2]);
tran (cceip1_out_ia_wdata[1], \cceip1_out_ia_wdata.r.part0 [1]);
tran (cceip1_out_ia_wdata[1], \cceip1_out_ia_wdata.f.unused0 [1]);
tran (cceip1_out_ia_wdata[0], \cceip1_out_ia_wdata.r.part0 [0]);
tran (cceip1_out_ia_wdata[0], \cceip1_out_ia_wdata.f.unused0 [0]);
tran (cceip1_out_ia_wdata[63], \cceip1_out_ia_wdata.r.part1 [31]);
tran (cceip1_out_ia_wdata[63], \cceip1_out_ia_wdata.f.tdata_lo [31]);
tran (cceip1_out_ia_wdata[62], \cceip1_out_ia_wdata.r.part1 [30]);
tran (cceip1_out_ia_wdata[62], \cceip1_out_ia_wdata.f.tdata_lo [30]);
tran (cceip1_out_ia_wdata[61], \cceip1_out_ia_wdata.r.part1 [29]);
tran (cceip1_out_ia_wdata[61], \cceip1_out_ia_wdata.f.tdata_lo [29]);
tran (cceip1_out_ia_wdata[60], \cceip1_out_ia_wdata.r.part1 [28]);
tran (cceip1_out_ia_wdata[60], \cceip1_out_ia_wdata.f.tdata_lo [28]);
tran (cceip1_out_ia_wdata[59], \cceip1_out_ia_wdata.r.part1 [27]);
tran (cceip1_out_ia_wdata[59], \cceip1_out_ia_wdata.f.tdata_lo [27]);
tran (cceip1_out_ia_wdata[58], \cceip1_out_ia_wdata.r.part1 [26]);
tran (cceip1_out_ia_wdata[58], \cceip1_out_ia_wdata.f.tdata_lo [26]);
tran (cceip1_out_ia_wdata[57], \cceip1_out_ia_wdata.r.part1 [25]);
tran (cceip1_out_ia_wdata[57], \cceip1_out_ia_wdata.f.tdata_lo [25]);
tran (cceip1_out_ia_wdata[56], \cceip1_out_ia_wdata.r.part1 [24]);
tran (cceip1_out_ia_wdata[56], \cceip1_out_ia_wdata.f.tdata_lo [24]);
tran (cceip1_out_ia_wdata[55], \cceip1_out_ia_wdata.r.part1 [23]);
tran (cceip1_out_ia_wdata[55], \cceip1_out_ia_wdata.f.tdata_lo [23]);
tran (cceip1_out_ia_wdata[54], \cceip1_out_ia_wdata.r.part1 [22]);
tran (cceip1_out_ia_wdata[54], \cceip1_out_ia_wdata.f.tdata_lo [22]);
tran (cceip1_out_ia_wdata[53], \cceip1_out_ia_wdata.r.part1 [21]);
tran (cceip1_out_ia_wdata[53], \cceip1_out_ia_wdata.f.tdata_lo [21]);
tran (cceip1_out_ia_wdata[52], \cceip1_out_ia_wdata.r.part1 [20]);
tran (cceip1_out_ia_wdata[52], \cceip1_out_ia_wdata.f.tdata_lo [20]);
tran (cceip1_out_ia_wdata[51], \cceip1_out_ia_wdata.r.part1 [19]);
tran (cceip1_out_ia_wdata[51], \cceip1_out_ia_wdata.f.tdata_lo [19]);
tran (cceip1_out_ia_wdata[50], \cceip1_out_ia_wdata.r.part1 [18]);
tran (cceip1_out_ia_wdata[50], \cceip1_out_ia_wdata.f.tdata_lo [18]);
tran (cceip1_out_ia_wdata[49], \cceip1_out_ia_wdata.r.part1 [17]);
tran (cceip1_out_ia_wdata[49], \cceip1_out_ia_wdata.f.tdata_lo [17]);
tran (cceip1_out_ia_wdata[48], \cceip1_out_ia_wdata.r.part1 [16]);
tran (cceip1_out_ia_wdata[48], \cceip1_out_ia_wdata.f.tdata_lo [16]);
tran (cceip1_out_ia_wdata[47], \cceip1_out_ia_wdata.r.part1 [15]);
tran (cceip1_out_ia_wdata[47], \cceip1_out_ia_wdata.f.tdata_lo [15]);
tran (cceip1_out_ia_wdata[46], \cceip1_out_ia_wdata.r.part1 [14]);
tran (cceip1_out_ia_wdata[46], \cceip1_out_ia_wdata.f.tdata_lo [14]);
tran (cceip1_out_ia_wdata[45], \cceip1_out_ia_wdata.r.part1 [13]);
tran (cceip1_out_ia_wdata[45], \cceip1_out_ia_wdata.f.tdata_lo [13]);
tran (cceip1_out_ia_wdata[44], \cceip1_out_ia_wdata.r.part1 [12]);
tran (cceip1_out_ia_wdata[44], \cceip1_out_ia_wdata.f.tdata_lo [12]);
tran (cceip1_out_ia_wdata[43], \cceip1_out_ia_wdata.r.part1 [11]);
tran (cceip1_out_ia_wdata[43], \cceip1_out_ia_wdata.f.tdata_lo [11]);
tran (cceip1_out_ia_wdata[42], \cceip1_out_ia_wdata.r.part1 [10]);
tran (cceip1_out_ia_wdata[42], \cceip1_out_ia_wdata.f.tdata_lo [10]);
tran (cceip1_out_ia_wdata[41], \cceip1_out_ia_wdata.r.part1 [9]);
tran (cceip1_out_ia_wdata[41], \cceip1_out_ia_wdata.f.tdata_lo [9]);
tran (cceip1_out_ia_wdata[40], \cceip1_out_ia_wdata.r.part1 [8]);
tran (cceip1_out_ia_wdata[40], \cceip1_out_ia_wdata.f.tdata_lo [8]);
tran (cceip1_out_ia_wdata[39], \cceip1_out_ia_wdata.r.part1 [7]);
tran (cceip1_out_ia_wdata[39], \cceip1_out_ia_wdata.f.tdata_lo [7]);
tran (cceip1_out_ia_wdata[38], \cceip1_out_ia_wdata.r.part1 [6]);
tran (cceip1_out_ia_wdata[38], \cceip1_out_ia_wdata.f.tdata_lo [6]);
tran (cceip1_out_ia_wdata[37], \cceip1_out_ia_wdata.r.part1 [5]);
tran (cceip1_out_ia_wdata[37], \cceip1_out_ia_wdata.f.tdata_lo [5]);
tran (cceip1_out_ia_wdata[36], \cceip1_out_ia_wdata.r.part1 [4]);
tran (cceip1_out_ia_wdata[36], \cceip1_out_ia_wdata.f.tdata_lo [4]);
tran (cceip1_out_ia_wdata[35], \cceip1_out_ia_wdata.r.part1 [3]);
tran (cceip1_out_ia_wdata[35], \cceip1_out_ia_wdata.f.tdata_lo [3]);
tran (cceip1_out_ia_wdata[34], \cceip1_out_ia_wdata.r.part1 [2]);
tran (cceip1_out_ia_wdata[34], \cceip1_out_ia_wdata.f.tdata_lo [2]);
tran (cceip1_out_ia_wdata[33], \cceip1_out_ia_wdata.r.part1 [1]);
tran (cceip1_out_ia_wdata[33], \cceip1_out_ia_wdata.f.tdata_lo [1]);
tran (cceip1_out_ia_wdata[32], \cceip1_out_ia_wdata.r.part1 [0]);
tran (cceip1_out_ia_wdata[32], \cceip1_out_ia_wdata.f.tdata_lo [0]);
tran (cceip1_out_ia_wdata[95], \cceip1_out_ia_wdata.r.part2 [31]);
tran (cceip1_out_ia_wdata[95], \cceip1_out_ia_wdata.f.tdata_hi [31]);
tran (cceip1_out_ia_wdata[94], \cceip1_out_ia_wdata.r.part2 [30]);
tran (cceip1_out_ia_wdata[94], \cceip1_out_ia_wdata.f.tdata_hi [30]);
tran (cceip1_out_ia_wdata[93], \cceip1_out_ia_wdata.r.part2 [29]);
tran (cceip1_out_ia_wdata[93], \cceip1_out_ia_wdata.f.tdata_hi [29]);
tran (cceip1_out_ia_wdata[92], \cceip1_out_ia_wdata.r.part2 [28]);
tran (cceip1_out_ia_wdata[92], \cceip1_out_ia_wdata.f.tdata_hi [28]);
tran (cceip1_out_ia_wdata[91], \cceip1_out_ia_wdata.r.part2 [27]);
tran (cceip1_out_ia_wdata[91], \cceip1_out_ia_wdata.f.tdata_hi [27]);
tran (cceip1_out_ia_wdata[90], \cceip1_out_ia_wdata.r.part2 [26]);
tran (cceip1_out_ia_wdata[90], \cceip1_out_ia_wdata.f.tdata_hi [26]);
tran (cceip1_out_ia_wdata[89], \cceip1_out_ia_wdata.r.part2 [25]);
tran (cceip1_out_ia_wdata[89], \cceip1_out_ia_wdata.f.tdata_hi [25]);
tran (cceip1_out_ia_wdata[88], \cceip1_out_ia_wdata.r.part2 [24]);
tran (cceip1_out_ia_wdata[88], \cceip1_out_ia_wdata.f.tdata_hi [24]);
tran (cceip1_out_ia_wdata[87], \cceip1_out_ia_wdata.r.part2 [23]);
tran (cceip1_out_ia_wdata[87], \cceip1_out_ia_wdata.f.tdata_hi [23]);
tran (cceip1_out_ia_wdata[86], \cceip1_out_ia_wdata.r.part2 [22]);
tran (cceip1_out_ia_wdata[86], \cceip1_out_ia_wdata.f.tdata_hi [22]);
tran (cceip1_out_ia_wdata[85], \cceip1_out_ia_wdata.r.part2 [21]);
tran (cceip1_out_ia_wdata[85], \cceip1_out_ia_wdata.f.tdata_hi [21]);
tran (cceip1_out_ia_wdata[84], \cceip1_out_ia_wdata.r.part2 [20]);
tran (cceip1_out_ia_wdata[84], \cceip1_out_ia_wdata.f.tdata_hi [20]);
tran (cceip1_out_ia_wdata[83], \cceip1_out_ia_wdata.r.part2 [19]);
tran (cceip1_out_ia_wdata[83], \cceip1_out_ia_wdata.f.tdata_hi [19]);
tran (cceip1_out_ia_wdata[82], \cceip1_out_ia_wdata.r.part2 [18]);
tran (cceip1_out_ia_wdata[82], \cceip1_out_ia_wdata.f.tdata_hi [18]);
tran (cceip1_out_ia_wdata[81], \cceip1_out_ia_wdata.r.part2 [17]);
tran (cceip1_out_ia_wdata[81], \cceip1_out_ia_wdata.f.tdata_hi [17]);
tran (cceip1_out_ia_wdata[80], \cceip1_out_ia_wdata.r.part2 [16]);
tran (cceip1_out_ia_wdata[80], \cceip1_out_ia_wdata.f.tdata_hi [16]);
tran (cceip1_out_ia_wdata[79], \cceip1_out_ia_wdata.r.part2 [15]);
tran (cceip1_out_ia_wdata[79], \cceip1_out_ia_wdata.f.tdata_hi [15]);
tran (cceip1_out_ia_wdata[78], \cceip1_out_ia_wdata.r.part2 [14]);
tran (cceip1_out_ia_wdata[78], \cceip1_out_ia_wdata.f.tdata_hi [14]);
tran (cceip1_out_ia_wdata[77], \cceip1_out_ia_wdata.r.part2 [13]);
tran (cceip1_out_ia_wdata[77], \cceip1_out_ia_wdata.f.tdata_hi [13]);
tran (cceip1_out_ia_wdata[76], \cceip1_out_ia_wdata.r.part2 [12]);
tran (cceip1_out_ia_wdata[76], \cceip1_out_ia_wdata.f.tdata_hi [12]);
tran (cceip1_out_ia_wdata[75], \cceip1_out_ia_wdata.r.part2 [11]);
tran (cceip1_out_ia_wdata[75], \cceip1_out_ia_wdata.f.tdata_hi [11]);
tran (cceip1_out_ia_wdata[74], \cceip1_out_ia_wdata.r.part2 [10]);
tran (cceip1_out_ia_wdata[74], \cceip1_out_ia_wdata.f.tdata_hi [10]);
tran (cceip1_out_ia_wdata[73], \cceip1_out_ia_wdata.r.part2 [9]);
tran (cceip1_out_ia_wdata[73], \cceip1_out_ia_wdata.f.tdata_hi [9]);
tran (cceip1_out_ia_wdata[72], \cceip1_out_ia_wdata.r.part2 [8]);
tran (cceip1_out_ia_wdata[72], \cceip1_out_ia_wdata.f.tdata_hi [8]);
tran (cceip1_out_ia_wdata[71], \cceip1_out_ia_wdata.r.part2 [7]);
tran (cceip1_out_ia_wdata[71], \cceip1_out_ia_wdata.f.tdata_hi [7]);
tran (cceip1_out_ia_wdata[70], \cceip1_out_ia_wdata.r.part2 [6]);
tran (cceip1_out_ia_wdata[70], \cceip1_out_ia_wdata.f.tdata_hi [6]);
tran (cceip1_out_ia_wdata[69], \cceip1_out_ia_wdata.r.part2 [5]);
tran (cceip1_out_ia_wdata[69], \cceip1_out_ia_wdata.f.tdata_hi [5]);
tran (cceip1_out_ia_wdata[68], \cceip1_out_ia_wdata.r.part2 [4]);
tran (cceip1_out_ia_wdata[68], \cceip1_out_ia_wdata.f.tdata_hi [4]);
tran (cceip1_out_ia_wdata[67], \cceip1_out_ia_wdata.r.part2 [3]);
tran (cceip1_out_ia_wdata[67], \cceip1_out_ia_wdata.f.tdata_hi [3]);
tran (cceip1_out_ia_wdata[66], \cceip1_out_ia_wdata.r.part2 [2]);
tran (cceip1_out_ia_wdata[66], \cceip1_out_ia_wdata.f.tdata_hi [2]);
tran (cceip1_out_ia_wdata[65], \cceip1_out_ia_wdata.r.part2 [1]);
tran (cceip1_out_ia_wdata[65], \cceip1_out_ia_wdata.f.tdata_hi [1]);
tran (cceip1_out_ia_wdata[64], \cceip1_out_ia_wdata.r.part2 [0]);
tran (cceip1_out_ia_wdata[64], \cceip1_out_ia_wdata.f.tdata_hi [0]);
tran (cceip1_out_ia_config[12], \cceip1_out_ia_config.r.part0 [12]);
tran (cceip1_out_ia_config[12], \cceip1_out_ia_config.f.op [3]);
tran (cceip1_out_ia_config[11], \cceip1_out_ia_config.r.part0 [11]);
tran (cceip1_out_ia_config[11], \cceip1_out_ia_config.f.op [2]);
tran (cceip1_out_ia_config[10], \cceip1_out_ia_config.r.part0 [10]);
tran (cceip1_out_ia_config[10], \cceip1_out_ia_config.f.op [1]);
tran (cceip1_out_ia_config[9], \cceip1_out_ia_config.r.part0 [9]);
tran (cceip1_out_ia_config[9], \cceip1_out_ia_config.f.op [0]);
tran (cceip1_out_ia_config[8], \cceip1_out_ia_config.r.part0 [8]);
tran (cceip1_out_ia_config[8], \cceip1_out_ia_config.f.addr [8]);
tran (cceip1_out_ia_config[7], \cceip1_out_ia_config.r.part0 [7]);
tran (cceip1_out_ia_config[7], \cceip1_out_ia_config.f.addr [7]);
tran (cceip1_out_ia_config[6], \cceip1_out_ia_config.r.part0 [6]);
tran (cceip1_out_ia_config[6], \cceip1_out_ia_config.f.addr [6]);
tran (cceip1_out_ia_config[5], \cceip1_out_ia_config.r.part0 [5]);
tran (cceip1_out_ia_config[5], \cceip1_out_ia_config.f.addr [5]);
tran (cceip1_out_ia_config[4], \cceip1_out_ia_config.r.part0 [4]);
tran (cceip1_out_ia_config[4], \cceip1_out_ia_config.f.addr [4]);
tran (cceip1_out_ia_config[3], \cceip1_out_ia_config.r.part0 [3]);
tran (cceip1_out_ia_config[3], \cceip1_out_ia_config.f.addr [3]);
tran (cceip1_out_ia_config[2], \cceip1_out_ia_config.r.part0 [2]);
tran (cceip1_out_ia_config[2], \cceip1_out_ia_config.f.addr [2]);
tran (cceip1_out_ia_config[1], \cceip1_out_ia_config.r.part0 [1]);
tran (cceip1_out_ia_config[1], \cceip1_out_ia_config.f.addr [1]);
tran (cceip1_out_ia_config[0], \cceip1_out_ia_config.r.part0 [0]);
tran (cceip1_out_ia_config[0], \cceip1_out_ia_config.f.addr [0]);
tran (cceip1_out_im_config[11], \cceip1_out_im_config.r.part0 [11]);
tran (cceip1_out_im_config[11], \cceip1_out_im_config.f.mode [1]);
tran (cceip1_out_im_config[10], \cceip1_out_im_config.r.part0 [10]);
tran (cceip1_out_im_config[10], \cceip1_out_im_config.f.mode [0]);
tran (cceip1_out_im_config[9], \cceip1_out_im_config.r.part0 [9]);
tran (cceip1_out_im_config[9], \cceip1_out_im_config.f.wr_credit_config [9]);
tran (cceip1_out_im_config[8], \cceip1_out_im_config.r.part0 [8]);
tran (cceip1_out_im_config[8], \cceip1_out_im_config.f.wr_credit_config [8]);
tran (cceip1_out_im_config[7], \cceip1_out_im_config.r.part0 [7]);
tran (cceip1_out_im_config[7], \cceip1_out_im_config.f.wr_credit_config [7]);
tran (cceip1_out_im_config[6], \cceip1_out_im_config.r.part0 [6]);
tran (cceip1_out_im_config[6], \cceip1_out_im_config.f.wr_credit_config [6]);
tran (cceip1_out_im_config[5], \cceip1_out_im_config.r.part0 [5]);
tran (cceip1_out_im_config[5], \cceip1_out_im_config.f.wr_credit_config [5]);
tran (cceip1_out_im_config[4], \cceip1_out_im_config.r.part0 [4]);
tran (cceip1_out_im_config[4], \cceip1_out_im_config.f.wr_credit_config [4]);
tran (cceip1_out_im_config[3], \cceip1_out_im_config.r.part0 [3]);
tran (cceip1_out_im_config[3], \cceip1_out_im_config.f.wr_credit_config [3]);
tran (cceip1_out_im_config[2], \cceip1_out_im_config.r.part0 [2]);
tran (cceip1_out_im_config[2], \cceip1_out_im_config.f.wr_credit_config [2]);
tran (cceip1_out_im_config[1], \cceip1_out_im_config.r.part0 [1]);
tran (cceip1_out_im_config[1], \cceip1_out_im_config.f.wr_credit_config [1]);
tran (cceip1_out_im_config[0], \cceip1_out_im_config.r.part0 [0]);
tran (cceip1_out_im_config[0], \cceip1_out_im_config.f.wr_credit_config [0]);
tran (cceip2_out_ia_wdata[31], \cceip2_out_ia_wdata.r.part0 [31]);
tran (cceip2_out_ia_wdata[31], \cceip2_out_ia_wdata.f.eob );
tran (cceip2_out_ia_wdata[30], \cceip2_out_ia_wdata.r.part0 [30]);
tran (cceip2_out_ia_wdata[30], \cceip2_out_ia_wdata.f.bytes_vld [7]);
tran (cceip2_out_ia_wdata[29], \cceip2_out_ia_wdata.r.part0 [29]);
tran (cceip2_out_ia_wdata[29], \cceip2_out_ia_wdata.f.bytes_vld [6]);
tran (cceip2_out_ia_wdata[28], \cceip2_out_ia_wdata.r.part0 [28]);
tran (cceip2_out_ia_wdata[28], \cceip2_out_ia_wdata.f.bytes_vld [5]);
tran (cceip2_out_ia_wdata[27], \cceip2_out_ia_wdata.r.part0 [27]);
tran (cceip2_out_ia_wdata[27], \cceip2_out_ia_wdata.f.bytes_vld [4]);
tran (cceip2_out_ia_wdata[26], \cceip2_out_ia_wdata.r.part0 [26]);
tran (cceip2_out_ia_wdata[26], \cceip2_out_ia_wdata.f.bytes_vld [3]);
tran (cceip2_out_ia_wdata[25], \cceip2_out_ia_wdata.r.part0 [25]);
tran (cceip2_out_ia_wdata[25], \cceip2_out_ia_wdata.f.bytes_vld [2]);
tran (cceip2_out_ia_wdata[24], \cceip2_out_ia_wdata.r.part0 [24]);
tran (cceip2_out_ia_wdata[24], \cceip2_out_ia_wdata.f.bytes_vld [1]);
tran (cceip2_out_ia_wdata[23], \cceip2_out_ia_wdata.r.part0 [23]);
tran (cceip2_out_ia_wdata[23], \cceip2_out_ia_wdata.f.bytes_vld [0]);
tran (cceip2_out_ia_wdata[22], \cceip2_out_ia_wdata.r.part0 [22]);
tran (cceip2_out_ia_wdata[22], \cceip2_out_ia_wdata.f.unused1 [7]);
tran (cceip2_out_ia_wdata[21], \cceip2_out_ia_wdata.r.part0 [21]);
tran (cceip2_out_ia_wdata[21], \cceip2_out_ia_wdata.f.unused1 [6]);
tran (cceip2_out_ia_wdata[20], \cceip2_out_ia_wdata.r.part0 [20]);
tran (cceip2_out_ia_wdata[20], \cceip2_out_ia_wdata.f.unused1 [5]);
tran (cceip2_out_ia_wdata[19], \cceip2_out_ia_wdata.r.part0 [19]);
tran (cceip2_out_ia_wdata[19], \cceip2_out_ia_wdata.f.unused1 [4]);
tran (cceip2_out_ia_wdata[18], \cceip2_out_ia_wdata.r.part0 [18]);
tran (cceip2_out_ia_wdata[18], \cceip2_out_ia_wdata.f.unused1 [3]);
tran (cceip2_out_ia_wdata[17], \cceip2_out_ia_wdata.r.part0 [17]);
tran (cceip2_out_ia_wdata[17], \cceip2_out_ia_wdata.f.unused1 [2]);
tran (cceip2_out_ia_wdata[16], \cceip2_out_ia_wdata.r.part0 [16]);
tran (cceip2_out_ia_wdata[16], \cceip2_out_ia_wdata.f.unused1 [1]);
tran (cceip2_out_ia_wdata[15], \cceip2_out_ia_wdata.r.part0 [15]);
tran (cceip2_out_ia_wdata[15], \cceip2_out_ia_wdata.f.unused1 [0]);
tran (cceip2_out_ia_wdata[14], \cceip2_out_ia_wdata.r.part0 [14]);
tran (cceip2_out_ia_wdata[14], \cceip2_out_ia_wdata.f.tid );
tran (cceip2_out_ia_wdata[13], \cceip2_out_ia_wdata.r.part0 [13]);
tran (cceip2_out_ia_wdata[13], \cceip2_out_ia_wdata.f.tuser [7]);
tran (cceip2_out_ia_wdata[12], \cceip2_out_ia_wdata.r.part0 [12]);
tran (cceip2_out_ia_wdata[12], \cceip2_out_ia_wdata.f.tuser [6]);
tran (cceip2_out_ia_wdata[11], \cceip2_out_ia_wdata.r.part0 [11]);
tran (cceip2_out_ia_wdata[11], \cceip2_out_ia_wdata.f.tuser [5]);
tran (cceip2_out_ia_wdata[10], \cceip2_out_ia_wdata.r.part0 [10]);
tran (cceip2_out_ia_wdata[10], \cceip2_out_ia_wdata.f.tuser [4]);
tran (cceip2_out_ia_wdata[9], \cceip2_out_ia_wdata.r.part0 [9]);
tran (cceip2_out_ia_wdata[9], \cceip2_out_ia_wdata.f.tuser [3]);
tran (cceip2_out_ia_wdata[8], \cceip2_out_ia_wdata.r.part0 [8]);
tran (cceip2_out_ia_wdata[8], \cceip2_out_ia_wdata.f.tuser [2]);
tran (cceip2_out_ia_wdata[7], \cceip2_out_ia_wdata.r.part0 [7]);
tran (cceip2_out_ia_wdata[7], \cceip2_out_ia_wdata.f.tuser [1]);
tran (cceip2_out_ia_wdata[6], \cceip2_out_ia_wdata.r.part0 [6]);
tran (cceip2_out_ia_wdata[6], \cceip2_out_ia_wdata.f.tuser [0]);
tran (cceip2_out_ia_wdata[5], \cceip2_out_ia_wdata.r.part0 [5]);
tran (cceip2_out_ia_wdata[5], \cceip2_out_ia_wdata.f.unused0 [5]);
tran (cceip2_out_ia_wdata[4], \cceip2_out_ia_wdata.r.part0 [4]);
tran (cceip2_out_ia_wdata[4], \cceip2_out_ia_wdata.f.unused0 [4]);
tran (cceip2_out_ia_wdata[3], \cceip2_out_ia_wdata.r.part0 [3]);
tran (cceip2_out_ia_wdata[3], \cceip2_out_ia_wdata.f.unused0 [3]);
tran (cceip2_out_ia_wdata[2], \cceip2_out_ia_wdata.r.part0 [2]);
tran (cceip2_out_ia_wdata[2], \cceip2_out_ia_wdata.f.unused0 [2]);
tran (cceip2_out_ia_wdata[1], \cceip2_out_ia_wdata.r.part0 [1]);
tran (cceip2_out_ia_wdata[1], \cceip2_out_ia_wdata.f.unused0 [1]);
tran (cceip2_out_ia_wdata[0], \cceip2_out_ia_wdata.r.part0 [0]);
tran (cceip2_out_ia_wdata[0], \cceip2_out_ia_wdata.f.unused0 [0]);
tran (cceip2_out_ia_wdata[63], \cceip2_out_ia_wdata.r.part1 [31]);
tran (cceip2_out_ia_wdata[63], \cceip2_out_ia_wdata.f.tdata_lo [31]);
tran (cceip2_out_ia_wdata[62], \cceip2_out_ia_wdata.r.part1 [30]);
tran (cceip2_out_ia_wdata[62], \cceip2_out_ia_wdata.f.tdata_lo [30]);
tran (cceip2_out_ia_wdata[61], \cceip2_out_ia_wdata.r.part1 [29]);
tran (cceip2_out_ia_wdata[61], \cceip2_out_ia_wdata.f.tdata_lo [29]);
tran (cceip2_out_ia_wdata[60], \cceip2_out_ia_wdata.r.part1 [28]);
tran (cceip2_out_ia_wdata[60], \cceip2_out_ia_wdata.f.tdata_lo [28]);
tran (cceip2_out_ia_wdata[59], \cceip2_out_ia_wdata.r.part1 [27]);
tran (cceip2_out_ia_wdata[59], \cceip2_out_ia_wdata.f.tdata_lo [27]);
tran (cceip2_out_ia_wdata[58], \cceip2_out_ia_wdata.r.part1 [26]);
tran (cceip2_out_ia_wdata[58], \cceip2_out_ia_wdata.f.tdata_lo [26]);
tran (cceip2_out_ia_wdata[57], \cceip2_out_ia_wdata.r.part1 [25]);
tran (cceip2_out_ia_wdata[57], \cceip2_out_ia_wdata.f.tdata_lo [25]);
tran (cceip2_out_ia_wdata[56], \cceip2_out_ia_wdata.r.part1 [24]);
tran (cceip2_out_ia_wdata[56], \cceip2_out_ia_wdata.f.tdata_lo [24]);
tran (cceip2_out_ia_wdata[55], \cceip2_out_ia_wdata.r.part1 [23]);
tran (cceip2_out_ia_wdata[55], \cceip2_out_ia_wdata.f.tdata_lo [23]);
tran (cceip2_out_ia_wdata[54], \cceip2_out_ia_wdata.r.part1 [22]);
tran (cceip2_out_ia_wdata[54], \cceip2_out_ia_wdata.f.tdata_lo [22]);
tran (cceip2_out_ia_wdata[53], \cceip2_out_ia_wdata.r.part1 [21]);
tran (cceip2_out_ia_wdata[53], \cceip2_out_ia_wdata.f.tdata_lo [21]);
tran (cceip2_out_ia_wdata[52], \cceip2_out_ia_wdata.r.part1 [20]);
tran (cceip2_out_ia_wdata[52], \cceip2_out_ia_wdata.f.tdata_lo [20]);
tran (cceip2_out_ia_wdata[51], \cceip2_out_ia_wdata.r.part1 [19]);
tran (cceip2_out_ia_wdata[51], \cceip2_out_ia_wdata.f.tdata_lo [19]);
tran (cceip2_out_ia_wdata[50], \cceip2_out_ia_wdata.r.part1 [18]);
tran (cceip2_out_ia_wdata[50], \cceip2_out_ia_wdata.f.tdata_lo [18]);
tran (cceip2_out_ia_wdata[49], \cceip2_out_ia_wdata.r.part1 [17]);
tran (cceip2_out_ia_wdata[49], \cceip2_out_ia_wdata.f.tdata_lo [17]);
tran (cceip2_out_ia_wdata[48], \cceip2_out_ia_wdata.r.part1 [16]);
tran (cceip2_out_ia_wdata[48], \cceip2_out_ia_wdata.f.tdata_lo [16]);
tran (cceip2_out_ia_wdata[47], \cceip2_out_ia_wdata.r.part1 [15]);
tran (cceip2_out_ia_wdata[47], \cceip2_out_ia_wdata.f.tdata_lo [15]);
tran (cceip2_out_ia_wdata[46], \cceip2_out_ia_wdata.r.part1 [14]);
tran (cceip2_out_ia_wdata[46], \cceip2_out_ia_wdata.f.tdata_lo [14]);
tran (cceip2_out_ia_wdata[45], \cceip2_out_ia_wdata.r.part1 [13]);
tran (cceip2_out_ia_wdata[45], \cceip2_out_ia_wdata.f.tdata_lo [13]);
tran (cceip2_out_ia_wdata[44], \cceip2_out_ia_wdata.r.part1 [12]);
tran (cceip2_out_ia_wdata[44], \cceip2_out_ia_wdata.f.tdata_lo [12]);
tran (cceip2_out_ia_wdata[43], \cceip2_out_ia_wdata.r.part1 [11]);
tran (cceip2_out_ia_wdata[43], \cceip2_out_ia_wdata.f.tdata_lo [11]);
tran (cceip2_out_ia_wdata[42], \cceip2_out_ia_wdata.r.part1 [10]);
tran (cceip2_out_ia_wdata[42], \cceip2_out_ia_wdata.f.tdata_lo [10]);
tran (cceip2_out_ia_wdata[41], \cceip2_out_ia_wdata.r.part1 [9]);
tran (cceip2_out_ia_wdata[41], \cceip2_out_ia_wdata.f.tdata_lo [9]);
tran (cceip2_out_ia_wdata[40], \cceip2_out_ia_wdata.r.part1 [8]);
tran (cceip2_out_ia_wdata[40], \cceip2_out_ia_wdata.f.tdata_lo [8]);
tran (cceip2_out_ia_wdata[39], \cceip2_out_ia_wdata.r.part1 [7]);
tran (cceip2_out_ia_wdata[39], \cceip2_out_ia_wdata.f.tdata_lo [7]);
tran (cceip2_out_ia_wdata[38], \cceip2_out_ia_wdata.r.part1 [6]);
tran (cceip2_out_ia_wdata[38], \cceip2_out_ia_wdata.f.tdata_lo [6]);
tran (cceip2_out_ia_wdata[37], \cceip2_out_ia_wdata.r.part1 [5]);
tran (cceip2_out_ia_wdata[37], \cceip2_out_ia_wdata.f.tdata_lo [5]);
tran (cceip2_out_ia_wdata[36], \cceip2_out_ia_wdata.r.part1 [4]);
tran (cceip2_out_ia_wdata[36], \cceip2_out_ia_wdata.f.tdata_lo [4]);
tran (cceip2_out_ia_wdata[35], \cceip2_out_ia_wdata.r.part1 [3]);
tran (cceip2_out_ia_wdata[35], \cceip2_out_ia_wdata.f.tdata_lo [3]);
tran (cceip2_out_ia_wdata[34], \cceip2_out_ia_wdata.r.part1 [2]);
tran (cceip2_out_ia_wdata[34], \cceip2_out_ia_wdata.f.tdata_lo [2]);
tran (cceip2_out_ia_wdata[33], \cceip2_out_ia_wdata.r.part1 [1]);
tran (cceip2_out_ia_wdata[33], \cceip2_out_ia_wdata.f.tdata_lo [1]);
tran (cceip2_out_ia_wdata[32], \cceip2_out_ia_wdata.r.part1 [0]);
tran (cceip2_out_ia_wdata[32], \cceip2_out_ia_wdata.f.tdata_lo [0]);
tran (cceip2_out_ia_wdata[95], \cceip2_out_ia_wdata.r.part2 [31]);
tran (cceip2_out_ia_wdata[95], \cceip2_out_ia_wdata.f.tdata_hi [31]);
tran (cceip2_out_ia_wdata[94], \cceip2_out_ia_wdata.r.part2 [30]);
tran (cceip2_out_ia_wdata[94], \cceip2_out_ia_wdata.f.tdata_hi [30]);
tran (cceip2_out_ia_wdata[93], \cceip2_out_ia_wdata.r.part2 [29]);
tran (cceip2_out_ia_wdata[93], \cceip2_out_ia_wdata.f.tdata_hi [29]);
tran (cceip2_out_ia_wdata[92], \cceip2_out_ia_wdata.r.part2 [28]);
tran (cceip2_out_ia_wdata[92], \cceip2_out_ia_wdata.f.tdata_hi [28]);
tran (cceip2_out_ia_wdata[91], \cceip2_out_ia_wdata.r.part2 [27]);
tran (cceip2_out_ia_wdata[91], \cceip2_out_ia_wdata.f.tdata_hi [27]);
tran (cceip2_out_ia_wdata[90], \cceip2_out_ia_wdata.r.part2 [26]);
tran (cceip2_out_ia_wdata[90], \cceip2_out_ia_wdata.f.tdata_hi [26]);
tran (cceip2_out_ia_wdata[89], \cceip2_out_ia_wdata.r.part2 [25]);
tran (cceip2_out_ia_wdata[89], \cceip2_out_ia_wdata.f.tdata_hi [25]);
tran (cceip2_out_ia_wdata[88], \cceip2_out_ia_wdata.r.part2 [24]);
tran (cceip2_out_ia_wdata[88], \cceip2_out_ia_wdata.f.tdata_hi [24]);
tran (cceip2_out_ia_wdata[87], \cceip2_out_ia_wdata.r.part2 [23]);
tran (cceip2_out_ia_wdata[87], \cceip2_out_ia_wdata.f.tdata_hi [23]);
tran (cceip2_out_ia_wdata[86], \cceip2_out_ia_wdata.r.part2 [22]);
tran (cceip2_out_ia_wdata[86], \cceip2_out_ia_wdata.f.tdata_hi [22]);
tran (cceip2_out_ia_wdata[85], \cceip2_out_ia_wdata.r.part2 [21]);
tran (cceip2_out_ia_wdata[85], \cceip2_out_ia_wdata.f.tdata_hi [21]);
tran (cceip2_out_ia_wdata[84], \cceip2_out_ia_wdata.r.part2 [20]);
tran (cceip2_out_ia_wdata[84], \cceip2_out_ia_wdata.f.tdata_hi [20]);
tran (cceip2_out_ia_wdata[83], \cceip2_out_ia_wdata.r.part2 [19]);
tran (cceip2_out_ia_wdata[83], \cceip2_out_ia_wdata.f.tdata_hi [19]);
tran (cceip2_out_ia_wdata[82], \cceip2_out_ia_wdata.r.part2 [18]);
tran (cceip2_out_ia_wdata[82], \cceip2_out_ia_wdata.f.tdata_hi [18]);
tran (cceip2_out_ia_wdata[81], \cceip2_out_ia_wdata.r.part2 [17]);
tran (cceip2_out_ia_wdata[81], \cceip2_out_ia_wdata.f.tdata_hi [17]);
tran (cceip2_out_ia_wdata[80], \cceip2_out_ia_wdata.r.part2 [16]);
tran (cceip2_out_ia_wdata[80], \cceip2_out_ia_wdata.f.tdata_hi [16]);
tran (cceip2_out_ia_wdata[79], \cceip2_out_ia_wdata.r.part2 [15]);
tran (cceip2_out_ia_wdata[79], \cceip2_out_ia_wdata.f.tdata_hi [15]);
tran (cceip2_out_ia_wdata[78], \cceip2_out_ia_wdata.r.part2 [14]);
tran (cceip2_out_ia_wdata[78], \cceip2_out_ia_wdata.f.tdata_hi [14]);
tran (cceip2_out_ia_wdata[77], \cceip2_out_ia_wdata.r.part2 [13]);
tran (cceip2_out_ia_wdata[77], \cceip2_out_ia_wdata.f.tdata_hi [13]);
tran (cceip2_out_ia_wdata[76], \cceip2_out_ia_wdata.r.part2 [12]);
tran (cceip2_out_ia_wdata[76], \cceip2_out_ia_wdata.f.tdata_hi [12]);
tran (cceip2_out_ia_wdata[75], \cceip2_out_ia_wdata.r.part2 [11]);
tran (cceip2_out_ia_wdata[75], \cceip2_out_ia_wdata.f.tdata_hi [11]);
tran (cceip2_out_ia_wdata[74], \cceip2_out_ia_wdata.r.part2 [10]);
tran (cceip2_out_ia_wdata[74], \cceip2_out_ia_wdata.f.tdata_hi [10]);
tran (cceip2_out_ia_wdata[73], \cceip2_out_ia_wdata.r.part2 [9]);
tran (cceip2_out_ia_wdata[73], \cceip2_out_ia_wdata.f.tdata_hi [9]);
tran (cceip2_out_ia_wdata[72], \cceip2_out_ia_wdata.r.part2 [8]);
tran (cceip2_out_ia_wdata[72], \cceip2_out_ia_wdata.f.tdata_hi [8]);
tran (cceip2_out_ia_wdata[71], \cceip2_out_ia_wdata.r.part2 [7]);
tran (cceip2_out_ia_wdata[71], \cceip2_out_ia_wdata.f.tdata_hi [7]);
tran (cceip2_out_ia_wdata[70], \cceip2_out_ia_wdata.r.part2 [6]);
tran (cceip2_out_ia_wdata[70], \cceip2_out_ia_wdata.f.tdata_hi [6]);
tran (cceip2_out_ia_wdata[69], \cceip2_out_ia_wdata.r.part2 [5]);
tran (cceip2_out_ia_wdata[69], \cceip2_out_ia_wdata.f.tdata_hi [5]);
tran (cceip2_out_ia_wdata[68], \cceip2_out_ia_wdata.r.part2 [4]);
tran (cceip2_out_ia_wdata[68], \cceip2_out_ia_wdata.f.tdata_hi [4]);
tran (cceip2_out_ia_wdata[67], \cceip2_out_ia_wdata.r.part2 [3]);
tran (cceip2_out_ia_wdata[67], \cceip2_out_ia_wdata.f.tdata_hi [3]);
tran (cceip2_out_ia_wdata[66], \cceip2_out_ia_wdata.r.part2 [2]);
tran (cceip2_out_ia_wdata[66], \cceip2_out_ia_wdata.f.tdata_hi [2]);
tran (cceip2_out_ia_wdata[65], \cceip2_out_ia_wdata.r.part2 [1]);
tran (cceip2_out_ia_wdata[65], \cceip2_out_ia_wdata.f.tdata_hi [1]);
tran (cceip2_out_ia_wdata[64], \cceip2_out_ia_wdata.r.part2 [0]);
tran (cceip2_out_ia_wdata[64], \cceip2_out_ia_wdata.f.tdata_hi [0]);
tran (cceip2_out_ia_config[12], \cceip2_out_ia_config.r.part0 [12]);
tran (cceip2_out_ia_config[12], \cceip2_out_ia_config.f.op [3]);
tran (cceip2_out_ia_config[11], \cceip2_out_ia_config.r.part0 [11]);
tran (cceip2_out_ia_config[11], \cceip2_out_ia_config.f.op [2]);
tran (cceip2_out_ia_config[10], \cceip2_out_ia_config.r.part0 [10]);
tran (cceip2_out_ia_config[10], \cceip2_out_ia_config.f.op [1]);
tran (cceip2_out_ia_config[9], \cceip2_out_ia_config.r.part0 [9]);
tran (cceip2_out_ia_config[9], \cceip2_out_ia_config.f.op [0]);
tran (cceip2_out_ia_config[8], \cceip2_out_ia_config.r.part0 [8]);
tran (cceip2_out_ia_config[8], \cceip2_out_ia_config.f.addr [8]);
tran (cceip2_out_ia_config[7], \cceip2_out_ia_config.r.part0 [7]);
tran (cceip2_out_ia_config[7], \cceip2_out_ia_config.f.addr [7]);
tran (cceip2_out_ia_config[6], \cceip2_out_ia_config.r.part0 [6]);
tran (cceip2_out_ia_config[6], \cceip2_out_ia_config.f.addr [6]);
tran (cceip2_out_ia_config[5], \cceip2_out_ia_config.r.part0 [5]);
tran (cceip2_out_ia_config[5], \cceip2_out_ia_config.f.addr [5]);
tran (cceip2_out_ia_config[4], \cceip2_out_ia_config.r.part0 [4]);
tran (cceip2_out_ia_config[4], \cceip2_out_ia_config.f.addr [4]);
tran (cceip2_out_ia_config[3], \cceip2_out_ia_config.r.part0 [3]);
tran (cceip2_out_ia_config[3], \cceip2_out_ia_config.f.addr [3]);
tran (cceip2_out_ia_config[2], \cceip2_out_ia_config.r.part0 [2]);
tran (cceip2_out_ia_config[2], \cceip2_out_ia_config.f.addr [2]);
tran (cceip2_out_ia_config[1], \cceip2_out_ia_config.r.part0 [1]);
tran (cceip2_out_ia_config[1], \cceip2_out_ia_config.f.addr [1]);
tran (cceip2_out_ia_config[0], \cceip2_out_ia_config.r.part0 [0]);
tran (cceip2_out_ia_config[0], \cceip2_out_ia_config.f.addr [0]);
tran (cceip2_out_im_config[11], \cceip2_out_im_config.r.part0 [11]);
tran (cceip2_out_im_config[11], \cceip2_out_im_config.f.mode [1]);
tran (cceip2_out_im_config[10], \cceip2_out_im_config.r.part0 [10]);
tran (cceip2_out_im_config[10], \cceip2_out_im_config.f.mode [0]);
tran (cceip2_out_im_config[9], \cceip2_out_im_config.r.part0 [9]);
tran (cceip2_out_im_config[9], \cceip2_out_im_config.f.wr_credit_config [9]);
tran (cceip2_out_im_config[8], \cceip2_out_im_config.r.part0 [8]);
tran (cceip2_out_im_config[8], \cceip2_out_im_config.f.wr_credit_config [8]);
tran (cceip2_out_im_config[7], \cceip2_out_im_config.r.part0 [7]);
tran (cceip2_out_im_config[7], \cceip2_out_im_config.f.wr_credit_config [7]);
tran (cceip2_out_im_config[6], \cceip2_out_im_config.r.part0 [6]);
tran (cceip2_out_im_config[6], \cceip2_out_im_config.f.wr_credit_config [6]);
tran (cceip2_out_im_config[5], \cceip2_out_im_config.r.part0 [5]);
tran (cceip2_out_im_config[5], \cceip2_out_im_config.f.wr_credit_config [5]);
tran (cceip2_out_im_config[4], \cceip2_out_im_config.r.part0 [4]);
tran (cceip2_out_im_config[4], \cceip2_out_im_config.f.wr_credit_config [4]);
tran (cceip2_out_im_config[3], \cceip2_out_im_config.r.part0 [3]);
tran (cceip2_out_im_config[3], \cceip2_out_im_config.f.wr_credit_config [3]);
tran (cceip2_out_im_config[2], \cceip2_out_im_config.r.part0 [2]);
tran (cceip2_out_im_config[2], \cceip2_out_im_config.f.wr_credit_config [2]);
tran (cceip2_out_im_config[1], \cceip2_out_im_config.r.part0 [1]);
tran (cceip2_out_im_config[1], \cceip2_out_im_config.f.wr_credit_config [1]);
tran (cceip2_out_im_config[0], \cceip2_out_im_config.r.part0 [0]);
tran (cceip2_out_im_config[0], \cceip2_out_im_config.f.wr_credit_config [0]);
tran (cceip3_out_ia_wdata[31], \cceip3_out_ia_wdata.r.part0 [31]);
tran (cceip3_out_ia_wdata[31], \cceip3_out_ia_wdata.f.eob );
tran (cceip3_out_ia_wdata[30], \cceip3_out_ia_wdata.r.part0 [30]);
tran (cceip3_out_ia_wdata[30], \cceip3_out_ia_wdata.f.bytes_vld [7]);
tran (cceip3_out_ia_wdata[29], \cceip3_out_ia_wdata.r.part0 [29]);
tran (cceip3_out_ia_wdata[29], \cceip3_out_ia_wdata.f.bytes_vld [6]);
tran (cceip3_out_ia_wdata[28], \cceip3_out_ia_wdata.r.part0 [28]);
tran (cceip3_out_ia_wdata[28], \cceip3_out_ia_wdata.f.bytes_vld [5]);
tran (cceip3_out_ia_wdata[27], \cceip3_out_ia_wdata.r.part0 [27]);
tran (cceip3_out_ia_wdata[27], \cceip3_out_ia_wdata.f.bytes_vld [4]);
tran (cceip3_out_ia_wdata[26], \cceip3_out_ia_wdata.r.part0 [26]);
tran (cceip3_out_ia_wdata[26], \cceip3_out_ia_wdata.f.bytes_vld [3]);
tran (cceip3_out_ia_wdata[25], \cceip3_out_ia_wdata.r.part0 [25]);
tran (cceip3_out_ia_wdata[25], \cceip3_out_ia_wdata.f.bytes_vld [2]);
tran (cceip3_out_ia_wdata[24], \cceip3_out_ia_wdata.r.part0 [24]);
tran (cceip3_out_ia_wdata[24], \cceip3_out_ia_wdata.f.bytes_vld [1]);
tran (cceip3_out_ia_wdata[23], \cceip3_out_ia_wdata.r.part0 [23]);
tran (cceip3_out_ia_wdata[23], \cceip3_out_ia_wdata.f.bytes_vld [0]);
tran (cceip3_out_ia_wdata[22], \cceip3_out_ia_wdata.r.part0 [22]);
tran (cceip3_out_ia_wdata[22], \cceip3_out_ia_wdata.f.unused1 [7]);
tran (cceip3_out_ia_wdata[21], \cceip3_out_ia_wdata.r.part0 [21]);
tran (cceip3_out_ia_wdata[21], \cceip3_out_ia_wdata.f.unused1 [6]);
tran (cceip3_out_ia_wdata[20], \cceip3_out_ia_wdata.r.part0 [20]);
tran (cceip3_out_ia_wdata[20], \cceip3_out_ia_wdata.f.unused1 [5]);
tran (cceip3_out_ia_wdata[19], \cceip3_out_ia_wdata.r.part0 [19]);
tran (cceip3_out_ia_wdata[19], \cceip3_out_ia_wdata.f.unused1 [4]);
tran (cceip3_out_ia_wdata[18], \cceip3_out_ia_wdata.r.part0 [18]);
tran (cceip3_out_ia_wdata[18], \cceip3_out_ia_wdata.f.unused1 [3]);
tran (cceip3_out_ia_wdata[17], \cceip3_out_ia_wdata.r.part0 [17]);
tran (cceip3_out_ia_wdata[17], \cceip3_out_ia_wdata.f.unused1 [2]);
tran (cceip3_out_ia_wdata[16], \cceip3_out_ia_wdata.r.part0 [16]);
tran (cceip3_out_ia_wdata[16], \cceip3_out_ia_wdata.f.unused1 [1]);
tran (cceip3_out_ia_wdata[15], \cceip3_out_ia_wdata.r.part0 [15]);
tran (cceip3_out_ia_wdata[15], \cceip3_out_ia_wdata.f.unused1 [0]);
tran (cceip3_out_ia_wdata[14], \cceip3_out_ia_wdata.r.part0 [14]);
tran (cceip3_out_ia_wdata[14], \cceip3_out_ia_wdata.f.tid );
tran (cceip3_out_ia_wdata[13], \cceip3_out_ia_wdata.r.part0 [13]);
tran (cceip3_out_ia_wdata[13], \cceip3_out_ia_wdata.f.tuser [7]);
tran (cceip3_out_ia_wdata[12], \cceip3_out_ia_wdata.r.part0 [12]);
tran (cceip3_out_ia_wdata[12], \cceip3_out_ia_wdata.f.tuser [6]);
tran (cceip3_out_ia_wdata[11], \cceip3_out_ia_wdata.r.part0 [11]);
tran (cceip3_out_ia_wdata[11], \cceip3_out_ia_wdata.f.tuser [5]);
tran (cceip3_out_ia_wdata[10], \cceip3_out_ia_wdata.r.part0 [10]);
tran (cceip3_out_ia_wdata[10], \cceip3_out_ia_wdata.f.tuser [4]);
tran (cceip3_out_ia_wdata[9], \cceip3_out_ia_wdata.r.part0 [9]);
tran (cceip3_out_ia_wdata[9], \cceip3_out_ia_wdata.f.tuser [3]);
tran (cceip3_out_ia_wdata[8], \cceip3_out_ia_wdata.r.part0 [8]);
tran (cceip3_out_ia_wdata[8], \cceip3_out_ia_wdata.f.tuser [2]);
tran (cceip3_out_ia_wdata[7], \cceip3_out_ia_wdata.r.part0 [7]);
tran (cceip3_out_ia_wdata[7], \cceip3_out_ia_wdata.f.tuser [1]);
tran (cceip3_out_ia_wdata[6], \cceip3_out_ia_wdata.r.part0 [6]);
tran (cceip3_out_ia_wdata[6], \cceip3_out_ia_wdata.f.tuser [0]);
tran (cceip3_out_ia_wdata[5], \cceip3_out_ia_wdata.r.part0 [5]);
tran (cceip3_out_ia_wdata[5], \cceip3_out_ia_wdata.f.unused0 [5]);
tran (cceip3_out_ia_wdata[4], \cceip3_out_ia_wdata.r.part0 [4]);
tran (cceip3_out_ia_wdata[4], \cceip3_out_ia_wdata.f.unused0 [4]);
tran (cceip3_out_ia_wdata[3], \cceip3_out_ia_wdata.r.part0 [3]);
tran (cceip3_out_ia_wdata[3], \cceip3_out_ia_wdata.f.unused0 [3]);
tran (cceip3_out_ia_wdata[2], \cceip3_out_ia_wdata.r.part0 [2]);
tran (cceip3_out_ia_wdata[2], \cceip3_out_ia_wdata.f.unused0 [2]);
tran (cceip3_out_ia_wdata[1], \cceip3_out_ia_wdata.r.part0 [1]);
tran (cceip3_out_ia_wdata[1], \cceip3_out_ia_wdata.f.unused0 [1]);
tran (cceip3_out_ia_wdata[0], \cceip3_out_ia_wdata.r.part0 [0]);
tran (cceip3_out_ia_wdata[0], \cceip3_out_ia_wdata.f.unused0 [0]);
tran (cceip3_out_ia_wdata[63], \cceip3_out_ia_wdata.r.part1 [31]);
tran (cceip3_out_ia_wdata[63], \cceip3_out_ia_wdata.f.tdata_lo [31]);
tran (cceip3_out_ia_wdata[62], \cceip3_out_ia_wdata.r.part1 [30]);
tran (cceip3_out_ia_wdata[62], \cceip3_out_ia_wdata.f.tdata_lo [30]);
tran (cceip3_out_ia_wdata[61], \cceip3_out_ia_wdata.r.part1 [29]);
tran (cceip3_out_ia_wdata[61], \cceip3_out_ia_wdata.f.tdata_lo [29]);
tran (cceip3_out_ia_wdata[60], \cceip3_out_ia_wdata.r.part1 [28]);
tran (cceip3_out_ia_wdata[60], \cceip3_out_ia_wdata.f.tdata_lo [28]);
tran (cceip3_out_ia_wdata[59], \cceip3_out_ia_wdata.r.part1 [27]);
tran (cceip3_out_ia_wdata[59], \cceip3_out_ia_wdata.f.tdata_lo [27]);
tran (cceip3_out_ia_wdata[58], \cceip3_out_ia_wdata.r.part1 [26]);
tran (cceip3_out_ia_wdata[58], \cceip3_out_ia_wdata.f.tdata_lo [26]);
tran (cceip3_out_ia_wdata[57], \cceip3_out_ia_wdata.r.part1 [25]);
tran (cceip3_out_ia_wdata[57], \cceip3_out_ia_wdata.f.tdata_lo [25]);
tran (cceip3_out_ia_wdata[56], \cceip3_out_ia_wdata.r.part1 [24]);
tran (cceip3_out_ia_wdata[56], \cceip3_out_ia_wdata.f.tdata_lo [24]);
tran (cceip3_out_ia_wdata[55], \cceip3_out_ia_wdata.r.part1 [23]);
tran (cceip3_out_ia_wdata[55], \cceip3_out_ia_wdata.f.tdata_lo [23]);
tran (cceip3_out_ia_wdata[54], \cceip3_out_ia_wdata.r.part1 [22]);
tran (cceip3_out_ia_wdata[54], \cceip3_out_ia_wdata.f.tdata_lo [22]);
tran (cceip3_out_ia_wdata[53], \cceip3_out_ia_wdata.r.part1 [21]);
tran (cceip3_out_ia_wdata[53], \cceip3_out_ia_wdata.f.tdata_lo [21]);
tran (cceip3_out_ia_wdata[52], \cceip3_out_ia_wdata.r.part1 [20]);
tran (cceip3_out_ia_wdata[52], \cceip3_out_ia_wdata.f.tdata_lo [20]);
tran (cceip3_out_ia_wdata[51], \cceip3_out_ia_wdata.r.part1 [19]);
tran (cceip3_out_ia_wdata[51], \cceip3_out_ia_wdata.f.tdata_lo [19]);
tran (cceip3_out_ia_wdata[50], \cceip3_out_ia_wdata.r.part1 [18]);
tran (cceip3_out_ia_wdata[50], \cceip3_out_ia_wdata.f.tdata_lo [18]);
tran (cceip3_out_ia_wdata[49], \cceip3_out_ia_wdata.r.part1 [17]);
tran (cceip3_out_ia_wdata[49], \cceip3_out_ia_wdata.f.tdata_lo [17]);
tran (cceip3_out_ia_wdata[48], \cceip3_out_ia_wdata.r.part1 [16]);
tran (cceip3_out_ia_wdata[48], \cceip3_out_ia_wdata.f.tdata_lo [16]);
tran (cceip3_out_ia_wdata[47], \cceip3_out_ia_wdata.r.part1 [15]);
tran (cceip3_out_ia_wdata[47], \cceip3_out_ia_wdata.f.tdata_lo [15]);
tran (cceip3_out_ia_wdata[46], \cceip3_out_ia_wdata.r.part1 [14]);
tran (cceip3_out_ia_wdata[46], \cceip3_out_ia_wdata.f.tdata_lo [14]);
tran (cceip3_out_ia_wdata[45], \cceip3_out_ia_wdata.r.part1 [13]);
tran (cceip3_out_ia_wdata[45], \cceip3_out_ia_wdata.f.tdata_lo [13]);
tran (cceip3_out_ia_wdata[44], \cceip3_out_ia_wdata.r.part1 [12]);
tran (cceip3_out_ia_wdata[44], \cceip3_out_ia_wdata.f.tdata_lo [12]);
tran (cceip3_out_ia_wdata[43], \cceip3_out_ia_wdata.r.part1 [11]);
tran (cceip3_out_ia_wdata[43], \cceip3_out_ia_wdata.f.tdata_lo [11]);
tran (cceip3_out_ia_wdata[42], \cceip3_out_ia_wdata.r.part1 [10]);
tran (cceip3_out_ia_wdata[42], \cceip3_out_ia_wdata.f.tdata_lo [10]);
tran (cceip3_out_ia_wdata[41], \cceip3_out_ia_wdata.r.part1 [9]);
tran (cceip3_out_ia_wdata[41], \cceip3_out_ia_wdata.f.tdata_lo [9]);
tran (cceip3_out_ia_wdata[40], \cceip3_out_ia_wdata.r.part1 [8]);
tran (cceip3_out_ia_wdata[40], \cceip3_out_ia_wdata.f.tdata_lo [8]);
tran (cceip3_out_ia_wdata[39], \cceip3_out_ia_wdata.r.part1 [7]);
tran (cceip3_out_ia_wdata[39], \cceip3_out_ia_wdata.f.tdata_lo [7]);
tran (cceip3_out_ia_wdata[38], \cceip3_out_ia_wdata.r.part1 [6]);
tran (cceip3_out_ia_wdata[38], \cceip3_out_ia_wdata.f.tdata_lo [6]);
tran (cceip3_out_ia_wdata[37], \cceip3_out_ia_wdata.r.part1 [5]);
tran (cceip3_out_ia_wdata[37], \cceip3_out_ia_wdata.f.tdata_lo [5]);
tran (cceip3_out_ia_wdata[36], \cceip3_out_ia_wdata.r.part1 [4]);
tran (cceip3_out_ia_wdata[36], \cceip3_out_ia_wdata.f.tdata_lo [4]);
tran (cceip3_out_ia_wdata[35], \cceip3_out_ia_wdata.r.part1 [3]);
tran (cceip3_out_ia_wdata[35], \cceip3_out_ia_wdata.f.tdata_lo [3]);
tran (cceip3_out_ia_wdata[34], \cceip3_out_ia_wdata.r.part1 [2]);
tran (cceip3_out_ia_wdata[34], \cceip3_out_ia_wdata.f.tdata_lo [2]);
tran (cceip3_out_ia_wdata[33], \cceip3_out_ia_wdata.r.part1 [1]);
tran (cceip3_out_ia_wdata[33], \cceip3_out_ia_wdata.f.tdata_lo [1]);
tran (cceip3_out_ia_wdata[32], \cceip3_out_ia_wdata.r.part1 [0]);
tran (cceip3_out_ia_wdata[32], \cceip3_out_ia_wdata.f.tdata_lo [0]);
tran (cceip3_out_ia_wdata[95], \cceip3_out_ia_wdata.r.part2 [31]);
tran (cceip3_out_ia_wdata[95], \cceip3_out_ia_wdata.f.tdata_hi [31]);
tran (cceip3_out_ia_wdata[94], \cceip3_out_ia_wdata.r.part2 [30]);
tran (cceip3_out_ia_wdata[94], \cceip3_out_ia_wdata.f.tdata_hi [30]);
tran (cceip3_out_ia_wdata[93], \cceip3_out_ia_wdata.r.part2 [29]);
tran (cceip3_out_ia_wdata[93], \cceip3_out_ia_wdata.f.tdata_hi [29]);
tran (cceip3_out_ia_wdata[92], \cceip3_out_ia_wdata.r.part2 [28]);
tran (cceip3_out_ia_wdata[92], \cceip3_out_ia_wdata.f.tdata_hi [28]);
tran (cceip3_out_ia_wdata[91], \cceip3_out_ia_wdata.r.part2 [27]);
tran (cceip3_out_ia_wdata[91], \cceip3_out_ia_wdata.f.tdata_hi [27]);
tran (cceip3_out_ia_wdata[90], \cceip3_out_ia_wdata.r.part2 [26]);
tran (cceip3_out_ia_wdata[90], \cceip3_out_ia_wdata.f.tdata_hi [26]);
tran (cceip3_out_ia_wdata[89], \cceip3_out_ia_wdata.r.part2 [25]);
tran (cceip3_out_ia_wdata[89], \cceip3_out_ia_wdata.f.tdata_hi [25]);
tran (cceip3_out_ia_wdata[88], \cceip3_out_ia_wdata.r.part2 [24]);
tran (cceip3_out_ia_wdata[88], \cceip3_out_ia_wdata.f.tdata_hi [24]);
tran (cceip3_out_ia_wdata[87], \cceip3_out_ia_wdata.r.part2 [23]);
tran (cceip3_out_ia_wdata[87], \cceip3_out_ia_wdata.f.tdata_hi [23]);
tran (cceip3_out_ia_wdata[86], \cceip3_out_ia_wdata.r.part2 [22]);
tran (cceip3_out_ia_wdata[86], \cceip3_out_ia_wdata.f.tdata_hi [22]);
tran (cceip3_out_ia_wdata[85], \cceip3_out_ia_wdata.r.part2 [21]);
tran (cceip3_out_ia_wdata[85], \cceip3_out_ia_wdata.f.tdata_hi [21]);
tran (cceip3_out_ia_wdata[84], \cceip3_out_ia_wdata.r.part2 [20]);
tran (cceip3_out_ia_wdata[84], \cceip3_out_ia_wdata.f.tdata_hi [20]);
tran (cceip3_out_ia_wdata[83], \cceip3_out_ia_wdata.r.part2 [19]);
tran (cceip3_out_ia_wdata[83], \cceip3_out_ia_wdata.f.tdata_hi [19]);
tran (cceip3_out_ia_wdata[82], \cceip3_out_ia_wdata.r.part2 [18]);
tran (cceip3_out_ia_wdata[82], \cceip3_out_ia_wdata.f.tdata_hi [18]);
tran (cceip3_out_ia_wdata[81], \cceip3_out_ia_wdata.r.part2 [17]);
tran (cceip3_out_ia_wdata[81], \cceip3_out_ia_wdata.f.tdata_hi [17]);
tran (cceip3_out_ia_wdata[80], \cceip3_out_ia_wdata.r.part2 [16]);
tran (cceip3_out_ia_wdata[80], \cceip3_out_ia_wdata.f.tdata_hi [16]);
tran (cceip3_out_ia_wdata[79], \cceip3_out_ia_wdata.r.part2 [15]);
tran (cceip3_out_ia_wdata[79], \cceip3_out_ia_wdata.f.tdata_hi [15]);
tran (cceip3_out_ia_wdata[78], \cceip3_out_ia_wdata.r.part2 [14]);
tran (cceip3_out_ia_wdata[78], \cceip3_out_ia_wdata.f.tdata_hi [14]);
tran (cceip3_out_ia_wdata[77], \cceip3_out_ia_wdata.r.part2 [13]);
tran (cceip3_out_ia_wdata[77], \cceip3_out_ia_wdata.f.tdata_hi [13]);
tran (cceip3_out_ia_wdata[76], \cceip3_out_ia_wdata.r.part2 [12]);
tran (cceip3_out_ia_wdata[76], \cceip3_out_ia_wdata.f.tdata_hi [12]);
tran (cceip3_out_ia_wdata[75], \cceip3_out_ia_wdata.r.part2 [11]);
tran (cceip3_out_ia_wdata[75], \cceip3_out_ia_wdata.f.tdata_hi [11]);
tran (cceip3_out_ia_wdata[74], \cceip3_out_ia_wdata.r.part2 [10]);
tran (cceip3_out_ia_wdata[74], \cceip3_out_ia_wdata.f.tdata_hi [10]);
tran (cceip3_out_ia_wdata[73], \cceip3_out_ia_wdata.r.part2 [9]);
tran (cceip3_out_ia_wdata[73], \cceip3_out_ia_wdata.f.tdata_hi [9]);
tran (cceip3_out_ia_wdata[72], \cceip3_out_ia_wdata.r.part2 [8]);
tran (cceip3_out_ia_wdata[72], \cceip3_out_ia_wdata.f.tdata_hi [8]);
tran (cceip3_out_ia_wdata[71], \cceip3_out_ia_wdata.r.part2 [7]);
tran (cceip3_out_ia_wdata[71], \cceip3_out_ia_wdata.f.tdata_hi [7]);
tran (cceip3_out_ia_wdata[70], \cceip3_out_ia_wdata.r.part2 [6]);
tran (cceip3_out_ia_wdata[70], \cceip3_out_ia_wdata.f.tdata_hi [6]);
tran (cceip3_out_ia_wdata[69], \cceip3_out_ia_wdata.r.part2 [5]);
tran (cceip3_out_ia_wdata[69], \cceip3_out_ia_wdata.f.tdata_hi [5]);
tran (cceip3_out_ia_wdata[68], \cceip3_out_ia_wdata.r.part2 [4]);
tran (cceip3_out_ia_wdata[68], \cceip3_out_ia_wdata.f.tdata_hi [4]);
tran (cceip3_out_ia_wdata[67], \cceip3_out_ia_wdata.r.part2 [3]);
tran (cceip3_out_ia_wdata[67], \cceip3_out_ia_wdata.f.tdata_hi [3]);
tran (cceip3_out_ia_wdata[66], \cceip3_out_ia_wdata.r.part2 [2]);
tran (cceip3_out_ia_wdata[66], \cceip3_out_ia_wdata.f.tdata_hi [2]);
tran (cceip3_out_ia_wdata[65], \cceip3_out_ia_wdata.r.part2 [1]);
tran (cceip3_out_ia_wdata[65], \cceip3_out_ia_wdata.f.tdata_hi [1]);
tran (cceip3_out_ia_wdata[64], \cceip3_out_ia_wdata.r.part2 [0]);
tran (cceip3_out_ia_wdata[64], \cceip3_out_ia_wdata.f.tdata_hi [0]);
tran (cceip3_out_ia_config[12], \cceip3_out_ia_config.r.part0 [12]);
tran (cceip3_out_ia_config[12], \cceip3_out_ia_config.f.op [3]);
tran (cceip3_out_ia_config[11], \cceip3_out_ia_config.r.part0 [11]);
tran (cceip3_out_ia_config[11], \cceip3_out_ia_config.f.op [2]);
tran (cceip3_out_ia_config[10], \cceip3_out_ia_config.r.part0 [10]);
tran (cceip3_out_ia_config[10], \cceip3_out_ia_config.f.op [1]);
tran (cceip3_out_ia_config[9], \cceip3_out_ia_config.r.part0 [9]);
tran (cceip3_out_ia_config[9], \cceip3_out_ia_config.f.op [0]);
tran (cceip3_out_ia_config[8], \cceip3_out_ia_config.r.part0 [8]);
tran (cceip3_out_ia_config[8], \cceip3_out_ia_config.f.addr [8]);
tran (cceip3_out_ia_config[7], \cceip3_out_ia_config.r.part0 [7]);
tran (cceip3_out_ia_config[7], \cceip3_out_ia_config.f.addr [7]);
tran (cceip3_out_ia_config[6], \cceip3_out_ia_config.r.part0 [6]);
tran (cceip3_out_ia_config[6], \cceip3_out_ia_config.f.addr [6]);
tran (cceip3_out_ia_config[5], \cceip3_out_ia_config.r.part0 [5]);
tran (cceip3_out_ia_config[5], \cceip3_out_ia_config.f.addr [5]);
tran (cceip3_out_ia_config[4], \cceip3_out_ia_config.r.part0 [4]);
tran (cceip3_out_ia_config[4], \cceip3_out_ia_config.f.addr [4]);
tran (cceip3_out_ia_config[3], \cceip3_out_ia_config.r.part0 [3]);
tran (cceip3_out_ia_config[3], \cceip3_out_ia_config.f.addr [3]);
tran (cceip3_out_ia_config[2], \cceip3_out_ia_config.r.part0 [2]);
tran (cceip3_out_ia_config[2], \cceip3_out_ia_config.f.addr [2]);
tran (cceip3_out_ia_config[1], \cceip3_out_ia_config.r.part0 [1]);
tran (cceip3_out_ia_config[1], \cceip3_out_ia_config.f.addr [1]);
tran (cceip3_out_ia_config[0], \cceip3_out_ia_config.r.part0 [0]);
tran (cceip3_out_ia_config[0], \cceip3_out_ia_config.f.addr [0]);
tran (cceip3_out_im_config[11], \cceip3_out_im_config.r.part0 [11]);
tran (cceip3_out_im_config[11], \cceip3_out_im_config.f.mode [1]);
tran (cceip3_out_im_config[10], \cceip3_out_im_config.r.part0 [10]);
tran (cceip3_out_im_config[10], \cceip3_out_im_config.f.mode [0]);
tran (cceip3_out_im_config[9], \cceip3_out_im_config.r.part0 [9]);
tran (cceip3_out_im_config[9], \cceip3_out_im_config.f.wr_credit_config [9]);
tran (cceip3_out_im_config[8], \cceip3_out_im_config.r.part0 [8]);
tran (cceip3_out_im_config[8], \cceip3_out_im_config.f.wr_credit_config [8]);
tran (cceip3_out_im_config[7], \cceip3_out_im_config.r.part0 [7]);
tran (cceip3_out_im_config[7], \cceip3_out_im_config.f.wr_credit_config [7]);
tran (cceip3_out_im_config[6], \cceip3_out_im_config.r.part0 [6]);
tran (cceip3_out_im_config[6], \cceip3_out_im_config.f.wr_credit_config [6]);
tran (cceip3_out_im_config[5], \cceip3_out_im_config.r.part0 [5]);
tran (cceip3_out_im_config[5], \cceip3_out_im_config.f.wr_credit_config [5]);
tran (cceip3_out_im_config[4], \cceip3_out_im_config.r.part0 [4]);
tran (cceip3_out_im_config[4], \cceip3_out_im_config.f.wr_credit_config [4]);
tran (cceip3_out_im_config[3], \cceip3_out_im_config.r.part0 [3]);
tran (cceip3_out_im_config[3], \cceip3_out_im_config.f.wr_credit_config [3]);
tran (cceip3_out_im_config[2], \cceip3_out_im_config.r.part0 [2]);
tran (cceip3_out_im_config[2], \cceip3_out_im_config.f.wr_credit_config [2]);
tran (cceip3_out_im_config[1], \cceip3_out_im_config.r.part0 [1]);
tran (cceip3_out_im_config[1], \cceip3_out_im_config.f.wr_credit_config [1]);
tran (cceip3_out_im_config[0], \cceip3_out_im_config.r.part0 [0]);
tran (cceip3_out_im_config[0], \cceip3_out_im_config.f.wr_credit_config [0]);
tran (cddip0_out_ia_wdata[31], \cddip0_out_ia_wdata.r.part0 [31]);
tran (cddip0_out_ia_wdata[31], \cddip0_out_ia_wdata.f.eob );
tran (cddip0_out_ia_wdata[30], \cddip0_out_ia_wdata.r.part0 [30]);
tran (cddip0_out_ia_wdata[30], \cddip0_out_ia_wdata.f.bytes_vld [7]);
tran (cddip0_out_ia_wdata[29], \cddip0_out_ia_wdata.r.part0 [29]);
tran (cddip0_out_ia_wdata[29], \cddip0_out_ia_wdata.f.bytes_vld [6]);
tran (cddip0_out_ia_wdata[28], \cddip0_out_ia_wdata.r.part0 [28]);
tran (cddip0_out_ia_wdata[28], \cddip0_out_ia_wdata.f.bytes_vld [5]);
tran (cddip0_out_ia_wdata[27], \cddip0_out_ia_wdata.r.part0 [27]);
tran (cddip0_out_ia_wdata[27], \cddip0_out_ia_wdata.f.bytes_vld [4]);
tran (cddip0_out_ia_wdata[26], \cddip0_out_ia_wdata.r.part0 [26]);
tran (cddip0_out_ia_wdata[26], \cddip0_out_ia_wdata.f.bytes_vld [3]);
tran (cddip0_out_ia_wdata[25], \cddip0_out_ia_wdata.r.part0 [25]);
tran (cddip0_out_ia_wdata[25], \cddip0_out_ia_wdata.f.bytes_vld [2]);
tran (cddip0_out_ia_wdata[24], \cddip0_out_ia_wdata.r.part0 [24]);
tran (cddip0_out_ia_wdata[24], \cddip0_out_ia_wdata.f.bytes_vld [1]);
tran (cddip0_out_ia_wdata[23], \cddip0_out_ia_wdata.r.part0 [23]);
tran (cddip0_out_ia_wdata[23], \cddip0_out_ia_wdata.f.bytes_vld [0]);
tran (cddip0_out_ia_wdata[22], \cddip0_out_ia_wdata.r.part0 [22]);
tran (cddip0_out_ia_wdata[22], \cddip0_out_ia_wdata.f.unused1 [7]);
tran (cddip0_out_ia_wdata[21], \cddip0_out_ia_wdata.r.part0 [21]);
tran (cddip0_out_ia_wdata[21], \cddip0_out_ia_wdata.f.unused1 [6]);
tran (cddip0_out_ia_wdata[20], \cddip0_out_ia_wdata.r.part0 [20]);
tran (cddip0_out_ia_wdata[20], \cddip0_out_ia_wdata.f.unused1 [5]);
tran (cddip0_out_ia_wdata[19], \cddip0_out_ia_wdata.r.part0 [19]);
tran (cddip0_out_ia_wdata[19], \cddip0_out_ia_wdata.f.unused1 [4]);
tran (cddip0_out_ia_wdata[18], \cddip0_out_ia_wdata.r.part0 [18]);
tran (cddip0_out_ia_wdata[18], \cddip0_out_ia_wdata.f.unused1 [3]);
tran (cddip0_out_ia_wdata[17], \cddip0_out_ia_wdata.r.part0 [17]);
tran (cddip0_out_ia_wdata[17], \cddip0_out_ia_wdata.f.unused1 [2]);
tran (cddip0_out_ia_wdata[16], \cddip0_out_ia_wdata.r.part0 [16]);
tran (cddip0_out_ia_wdata[16], \cddip0_out_ia_wdata.f.unused1 [1]);
tran (cddip0_out_ia_wdata[15], \cddip0_out_ia_wdata.r.part0 [15]);
tran (cddip0_out_ia_wdata[15], \cddip0_out_ia_wdata.f.unused1 [0]);
tran (cddip0_out_ia_wdata[14], \cddip0_out_ia_wdata.r.part0 [14]);
tran (cddip0_out_ia_wdata[14], \cddip0_out_ia_wdata.f.tid );
tran (cddip0_out_ia_wdata[13], \cddip0_out_ia_wdata.r.part0 [13]);
tran (cddip0_out_ia_wdata[13], \cddip0_out_ia_wdata.f.tuser [7]);
tran (cddip0_out_ia_wdata[12], \cddip0_out_ia_wdata.r.part0 [12]);
tran (cddip0_out_ia_wdata[12], \cddip0_out_ia_wdata.f.tuser [6]);
tran (cddip0_out_ia_wdata[11], \cddip0_out_ia_wdata.r.part0 [11]);
tran (cddip0_out_ia_wdata[11], \cddip0_out_ia_wdata.f.tuser [5]);
tran (cddip0_out_ia_wdata[10], \cddip0_out_ia_wdata.r.part0 [10]);
tran (cddip0_out_ia_wdata[10], \cddip0_out_ia_wdata.f.tuser [4]);
tran (cddip0_out_ia_wdata[9], \cddip0_out_ia_wdata.r.part0 [9]);
tran (cddip0_out_ia_wdata[9], \cddip0_out_ia_wdata.f.tuser [3]);
tran (cddip0_out_ia_wdata[8], \cddip0_out_ia_wdata.r.part0 [8]);
tran (cddip0_out_ia_wdata[8], \cddip0_out_ia_wdata.f.tuser [2]);
tran (cddip0_out_ia_wdata[7], \cddip0_out_ia_wdata.r.part0 [7]);
tran (cddip0_out_ia_wdata[7], \cddip0_out_ia_wdata.f.tuser [1]);
tran (cddip0_out_ia_wdata[6], \cddip0_out_ia_wdata.r.part0 [6]);
tran (cddip0_out_ia_wdata[6], \cddip0_out_ia_wdata.f.tuser [0]);
tran (cddip0_out_ia_wdata[5], \cddip0_out_ia_wdata.r.part0 [5]);
tran (cddip0_out_ia_wdata[5], \cddip0_out_ia_wdata.f.unused0 [5]);
tran (cddip0_out_ia_wdata[4], \cddip0_out_ia_wdata.r.part0 [4]);
tran (cddip0_out_ia_wdata[4], \cddip0_out_ia_wdata.f.unused0 [4]);
tran (cddip0_out_ia_wdata[3], \cddip0_out_ia_wdata.r.part0 [3]);
tran (cddip0_out_ia_wdata[3], \cddip0_out_ia_wdata.f.unused0 [3]);
tran (cddip0_out_ia_wdata[2], \cddip0_out_ia_wdata.r.part0 [2]);
tran (cddip0_out_ia_wdata[2], \cddip0_out_ia_wdata.f.unused0 [2]);
tran (cddip0_out_ia_wdata[1], \cddip0_out_ia_wdata.r.part0 [1]);
tran (cddip0_out_ia_wdata[1], \cddip0_out_ia_wdata.f.unused0 [1]);
tran (cddip0_out_ia_wdata[0], \cddip0_out_ia_wdata.r.part0 [0]);
tran (cddip0_out_ia_wdata[0], \cddip0_out_ia_wdata.f.unused0 [0]);
tran (cddip0_out_ia_wdata[63], \cddip0_out_ia_wdata.r.part1 [31]);
tran (cddip0_out_ia_wdata[63], \cddip0_out_ia_wdata.f.tdata_lo [31]);
tran (cddip0_out_ia_wdata[62], \cddip0_out_ia_wdata.r.part1 [30]);
tran (cddip0_out_ia_wdata[62], \cddip0_out_ia_wdata.f.tdata_lo [30]);
tran (cddip0_out_ia_wdata[61], \cddip0_out_ia_wdata.r.part1 [29]);
tran (cddip0_out_ia_wdata[61], \cddip0_out_ia_wdata.f.tdata_lo [29]);
tran (cddip0_out_ia_wdata[60], \cddip0_out_ia_wdata.r.part1 [28]);
tran (cddip0_out_ia_wdata[60], \cddip0_out_ia_wdata.f.tdata_lo [28]);
tran (cddip0_out_ia_wdata[59], \cddip0_out_ia_wdata.r.part1 [27]);
tran (cddip0_out_ia_wdata[59], \cddip0_out_ia_wdata.f.tdata_lo [27]);
tran (cddip0_out_ia_wdata[58], \cddip0_out_ia_wdata.r.part1 [26]);
tran (cddip0_out_ia_wdata[58], \cddip0_out_ia_wdata.f.tdata_lo [26]);
tran (cddip0_out_ia_wdata[57], \cddip0_out_ia_wdata.r.part1 [25]);
tran (cddip0_out_ia_wdata[57], \cddip0_out_ia_wdata.f.tdata_lo [25]);
tran (cddip0_out_ia_wdata[56], \cddip0_out_ia_wdata.r.part1 [24]);
tran (cddip0_out_ia_wdata[56], \cddip0_out_ia_wdata.f.tdata_lo [24]);
tran (cddip0_out_ia_wdata[55], \cddip0_out_ia_wdata.r.part1 [23]);
tran (cddip0_out_ia_wdata[55], \cddip0_out_ia_wdata.f.tdata_lo [23]);
tran (cddip0_out_ia_wdata[54], \cddip0_out_ia_wdata.r.part1 [22]);
tran (cddip0_out_ia_wdata[54], \cddip0_out_ia_wdata.f.tdata_lo [22]);
tran (cddip0_out_ia_wdata[53], \cddip0_out_ia_wdata.r.part1 [21]);
tran (cddip0_out_ia_wdata[53], \cddip0_out_ia_wdata.f.tdata_lo [21]);
tran (cddip0_out_ia_wdata[52], \cddip0_out_ia_wdata.r.part1 [20]);
tran (cddip0_out_ia_wdata[52], \cddip0_out_ia_wdata.f.tdata_lo [20]);
tran (cddip0_out_ia_wdata[51], \cddip0_out_ia_wdata.r.part1 [19]);
tran (cddip0_out_ia_wdata[51], \cddip0_out_ia_wdata.f.tdata_lo [19]);
tran (cddip0_out_ia_wdata[50], \cddip0_out_ia_wdata.r.part1 [18]);
tran (cddip0_out_ia_wdata[50], \cddip0_out_ia_wdata.f.tdata_lo [18]);
tran (cddip0_out_ia_wdata[49], \cddip0_out_ia_wdata.r.part1 [17]);
tran (cddip0_out_ia_wdata[49], \cddip0_out_ia_wdata.f.tdata_lo [17]);
tran (cddip0_out_ia_wdata[48], \cddip0_out_ia_wdata.r.part1 [16]);
tran (cddip0_out_ia_wdata[48], \cddip0_out_ia_wdata.f.tdata_lo [16]);
tran (cddip0_out_ia_wdata[47], \cddip0_out_ia_wdata.r.part1 [15]);
tran (cddip0_out_ia_wdata[47], \cddip0_out_ia_wdata.f.tdata_lo [15]);
tran (cddip0_out_ia_wdata[46], \cddip0_out_ia_wdata.r.part1 [14]);
tran (cddip0_out_ia_wdata[46], \cddip0_out_ia_wdata.f.tdata_lo [14]);
tran (cddip0_out_ia_wdata[45], \cddip0_out_ia_wdata.r.part1 [13]);
tran (cddip0_out_ia_wdata[45], \cddip0_out_ia_wdata.f.tdata_lo [13]);
tran (cddip0_out_ia_wdata[44], \cddip0_out_ia_wdata.r.part1 [12]);
tran (cddip0_out_ia_wdata[44], \cddip0_out_ia_wdata.f.tdata_lo [12]);
tran (cddip0_out_ia_wdata[43], \cddip0_out_ia_wdata.r.part1 [11]);
tran (cddip0_out_ia_wdata[43], \cddip0_out_ia_wdata.f.tdata_lo [11]);
tran (cddip0_out_ia_wdata[42], \cddip0_out_ia_wdata.r.part1 [10]);
tran (cddip0_out_ia_wdata[42], \cddip0_out_ia_wdata.f.tdata_lo [10]);
tran (cddip0_out_ia_wdata[41], \cddip0_out_ia_wdata.r.part1 [9]);
tran (cddip0_out_ia_wdata[41], \cddip0_out_ia_wdata.f.tdata_lo [9]);
tran (cddip0_out_ia_wdata[40], \cddip0_out_ia_wdata.r.part1 [8]);
tran (cddip0_out_ia_wdata[40], \cddip0_out_ia_wdata.f.tdata_lo [8]);
tran (cddip0_out_ia_wdata[39], \cddip0_out_ia_wdata.r.part1 [7]);
tran (cddip0_out_ia_wdata[39], \cddip0_out_ia_wdata.f.tdata_lo [7]);
tran (cddip0_out_ia_wdata[38], \cddip0_out_ia_wdata.r.part1 [6]);
tran (cddip0_out_ia_wdata[38], \cddip0_out_ia_wdata.f.tdata_lo [6]);
tran (cddip0_out_ia_wdata[37], \cddip0_out_ia_wdata.r.part1 [5]);
tran (cddip0_out_ia_wdata[37], \cddip0_out_ia_wdata.f.tdata_lo [5]);
tran (cddip0_out_ia_wdata[36], \cddip0_out_ia_wdata.r.part1 [4]);
tran (cddip0_out_ia_wdata[36], \cddip0_out_ia_wdata.f.tdata_lo [4]);
tran (cddip0_out_ia_wdata[35], \cddip0_out_ia_wdata.r.part1 [3]);
tran (cddip0_out_ia_wdata[35], \cddip0_out_ia_wdata.f.tdata_lo [3]);
tran (cddip0_out_ia_wdata[34], \cddip0_out_ia_wdata.r.part1 [2]);
tran (cddip0_out_ia_wdata[34], \cddip0_out_ia_wdata.f.tdata_lo [2]);
tran (cddip0_out_ia_wdata[33], \cddip0_out_ia_wdata.r.part1 [1]);
tran (cddip0_out_ia_wdata[33], \cddip0_out_ia_wdata.f.tdata_lo [1]);
tran (cddip0_out_ia_wdata[32], \cddip0_out_ia_wdata.r.part1 [0]);
tran (cddip0_out_ia_wdata[32], \cddip0_out_ia_wdata.f.tdata_lo [0]);
tran (cddip0_out_ia_wdata[95], \cddip0_out_ia_wdata.r.part2 [31]);
tran (cddip0_out_ia_wdata[95], \cddip0_out_ia_wdata.f.tdata_hi [31]);
tran (cddip0_out_ia_wdata[94], \cddip0_out_ia_wdata.r.part2 [30]);
tran (cddip0_out_ia_wdata[94], \cddip0_out_ia_wdata.f.tdata_hi [30]);
tran (cddip0_out_ia_wdata[93], \cddip0_out_ia_wdata.r.part2 [29]);
tran (cddip0_out_ia_wdata[93], \cddip0_out_ia_wdata.f.tdata_hi [29]);
tran (cddip0_out_ia_wdata[92], \cddip0_out_ia_wdata.r.part2 [28]);
tran (cddip0_out_ia_wdata[92], \cddip0_out_ia_wdata.f.tdata_hi [28]);
tran (cddip0_out_ia_wdata[91], \cddip0_out_ia_wdata.r.part2 [27]);
tran (cddip0_out_ia_wdata[91], \cddip0_out_ia_wdata.f.tdata_hi [27]);
tran (cddip0_out_ia_wdata[90], \cddip0_out_ia_wdata.r.part2 [26]);
tran (cddip0_out_ia_wdata[90], \cddip0_out_ia_wdata.f.tdata_hi [26]);
tran (cddip0_out_ia_wdata[89], \cddip0_out_ia_wdata.r.part2 [25]);
tran (cddip0_out_ia_wdata[89], \cddip0_out_ia_wdata.f.tdata_hi [25]);
tran (cddip0_out_ia_wdata[88], \cddip0_out_ia_wdata.r.part2 [24]);
tran (cddip0_out_ia_wdata[88], \cddip0_out_ia_wdata.f.tdata_hi [24]);
tran (cddip0_out_ia_wdata[87], \cddip0_out_ia_wdata.r.part2 [23]);
tran (cddip0_out_ia_wdata[87], \cddip0_out_ia_wdata.f.tdata_hi [23]);
tran (cddip0_out_ia_wdata[86], \cddip0_out_ia_wdata.r.part2 [22]);
tran (cddip0_out_ia_wdata[86], \cddip0_out_ia_wdata.f.tdata_hi [22]);
tran (cddip0_out_ia_wdata[85], \cddip0_out_ia_wdata.r.part2 [21]);
tran (cddip0_out_ia_wdata[85], \cddip0_out_ia_wdata.f.tdata_hi [21]);
tran (cddip0_out_ia_wdata[84], \cddip0_out_ia_wdata.r.part2 [20]);
tran (cddip0_out_ia_wdata[84], \cddip0_out_ia_wdata.f.tdata_hi [20]);
tran (cddip0_out_ia_wdata[83], \cddip0_out_ia_wdata.r.part2 [19]);
tran (cddip0_out_ia_wdata[83], \cddip0_out_ia_wdata.f.tdata_hi [19]);
tran (cddip0_out_ia_wdata[82], \cddip0_out_ia_wdata.r.part2 [18]);
tran (cddip0_out_ia_wdata[82], \cddip0_out_ia_wdata.f.tdata_hi [18]);
tran (cddip0_out_ia_wdata[81], \cddip0_out_ia_wdata.r.part2 [17]);
tran (cddip0_out_ia_wdata[81], \cddip0_out_ia_wdata.f.tdata_hi [17]);
tran (cddip0_out_ia_wdata[80], \cddip0_out_ia_wdata.r.part2 [16]);
tran (cddip0_out_ia_wdata[80], \cddip0_out_ia_wdata.f.tdata_hi [16]);
tran (cddip0_out_ia_wdata[79], \cddip0_out_ia_wdata.r.part2 [15]);
tran (cddip0_out_ia_wdata[79], \cddip0_out_ia_wdata.f.tdata_hi [15]);
tran (cddip0_out_ia_wdata[78], \cddip0_out_ia_wdata.r.part2 [14]);
tran (cddip0_out_ia_wdata[78], \cddip0_out_ia_wdata.f.tdata_hi [14]);
tran (cddip0_out_ia_wdata[77], \cddip0_out_ia_wdata.r.part2 [13]);
tran (cddip0_out_ia_wdata[77], \cddip0_out_ia_wdata.f.tdata_hi [13]);
tran (cddip0_out_ia_wdata[76], \cddip0_out_ia_wdata.r.part2 [12]);
tran (cddip0_out_ia_wdata[76], \cddip0_out_ia_wdata.f.tdata_hi [12]);
tran (cddip0_out_ia_wdata[75], \cddip0_out_ia_wdata.r.part2 [11]);
tran (cddip0_out_ia_wdata[75], \cddip0_out_ia_wdata.f.tdata_hi [11]);
tran (cddip0_out_ia_wdata[74], \cddip0_out_ia_wdata.r.part2 [10]);
tran (cddip0_out_ia_wdata[74], \cddip0_out_ia_wdata.f.tdata_hi [10]);
tran (cddip0_out_ia_wdata[73], \cddip0_out_ia_wdata.r.part2 [9]);
tran (cddip0_out_ia_wdata[73], \cddip0_out_ia_wdata.f.tdata_hi [9]);
tran (cddip0_out_ia_wdata[72], \cddip0_out_ia_wdata.r.part2 [8]);
tran (cddip0_out_ia_wdata[72], \cddip0_out_ia_wdata.f.tdata_hi [8]);
tran (cddip0_out_ia_wdata[71], \cddip0_out_ia_wdata.r.part2 [7]);
tran (cddip0_out_ia_wdata[71], \cddip0_out_ia_wdata.f.tdata_hi [7]);
tran (cddip0_out_ia_wdata[70], \cddip0_out_ia_wdata.r.part2 [6]);
tran (cddip0_out_ia_wdata[70], \cddip0_out_ia_wdata.f.tdata_hi [6]);
tran (cddip0_out_ia_wdata[69], \cddip0_out_ia_wdata.r.part2 [5]);
tran (cddip0_out_ia_wdata[69], \cddip0_out_ia_wdata.f.tdata_hi [5]);
tran (cddip0_out_ia_wdata[68], \cddip0_out_ia_wdata.r.part2 [4]);
tran (cddip0_out_ia_wdata[68], \cddip0_out_ia_wdata.f.tdata_hi [4]);
tran (cddip0_out_ia_wdata[67], \cddip0_out_ia_wdata.r.part2 [3]);
tran (cddip0_out_ia_wdata[67], \cddip0_out_ia_wdata.f.tdata_hi [3]);
tran (cddip0_out_ia_wdata[66], \cddip0_out_ia_wdata.r.part2 [2]);
tran (cddip0_out_ia_wdata[66], \cddip0_out_ia_wdata.f.tdata_hi [2]);
tran (cddip0_out_ia_wdata[65], \cddip0_out_ia_wdata.r.part2 [1]);
tran (cddip0_out_ia_wdata[65], \cddip0_out_ia_wdata.f.tdata_hi [1]);
tran (cddip0_out_ia_wdata[64], \cddip0_out_ia_wdata.r.part2 [0]);
tran (cddip0_out_ia_wdata[64], \cddip0_out_ia_wdata.f.tdata_hi [0]);
tran (cddip0_out_ia_config[12], \cddip0_out_ia_config.r.part0 [12]);
tran (cddip0_out_ia_config[12], \cddip0_out_ia_config.f.op [3]);
tran (cddip0_out_ia_config[11], \cddip0_out_ia_config.r.part0 [11]);
tran (cddip0_out_ia_config[11], \cddip0_out_ia_config.f.op [2]);
tran (cddip0_out_ia_config[10], \cddip0_out_ia_config.r.part0 [10]);
tran (cddip0_out_ia_config[10], \cddip0_out_ia_config.f.op [1]);
tran (cddip0_out_ia_config[9], \cddip0_out_ia_config.r.part0 [9]);
tran (cddip0_out_ia_config[9], \cddip0_out_ia_config.f.op [0]);
tran (cddip0_out_ia_config[8], \cddip0_out_ia_config.r.part0 [8]);
tran (cddip0_out_ia_config[8], \cddip0_out_ia_config.f.addr [8]);
tran (cddip0_out_ia_config[7], \cddip0_out_ia_config.r.part0 [7]);
tran (cddip0_out_ia_config[7], \cddip0_out_ia_config.f.addr [7]);
tran (cddip0_out_ia_config[6], \cddip0_out_ia_config.r.part0 [6]);
tran (cddip0_out_ia_config[6], \cddip0_out_ia_config.f.addr [6]);
tran (cddip0_out_ia_config[5], \cddip0_out_ia_config.r.part0 [5]);
tran (cddip0_out_ia_config[5], \cddip0_out_ia_config.f.addr [5]);
tran (cddip0_out_ia_config[4], \cddip0_out_ia_config.r.part0 [4]);
tran (cddip0_out_ia_config[4], \cddip0_out_ia_config.f.addr [4]);
tran (cddip0_out_ia_config[3], \cddip0_out_ia_config.r.part0 [3]);
tran (cddip0_out_ia_config[3], \cddip0_out_ia_config.f.addr [3]);
tran (cddip0_out_ia_config[2], \cddip0_out_ia_config.r.part0 [2]);
tran (cddip0_out_ia_config[2], \cddip0_out_ia_config.f.addr [2]);
tran (cddip0_out_ia_config[1], \cddip0_out_ia_config.r.part0 [1]);
tran (cddip0_out_ia_config[1], \cddip0_out_ia_config.f.addr [1]);
tran (cddip0_out_ia_config[0], \cddip0_out_ia_config.r.part0 [0]);
tran (cddip0_out_ia_config[0], \cddip0_out_ia_config.f.addr [0]);
tran (cddip0_out_im_config[11], \cddip0_out_im_config.r.part0 [11]);
tran (cddip0_out_im_config[11], \cddip0_out_im_config.f.mode [1]);
tran (cddip0_out_im_config[10], \cddip0_out_im_config.r.part0 [10]);
tran (cddip0_out_im_config[10], \cddip0_out_im_config.f.mode [0]);
tran (cddip0_out_im_config[9], \cddip0_out_im_config.r.part0 [9]);
tran (cddip0_out_im_config[9], \cddip0_out_im_config.f.wr_credit_config [9]);
tran (cddip0_out_im_config[8], \cddip0_out_im_config.r.part0 [8]);
tran (cddip0_out_im_config[8], \cddip0_out_im_config.f.wr_credit_config [8]);
tran (cddip0_out_im_config[7], \cddip0_out_im_config.r.part0 [7]);
tran (cddip0_out_im_config[7], \cddip0_out_im_config.f.wr_credit_config [7]);
tran (cddip0_out_im_config[6], \cddip0_out_im_config.r.part0 [6]);
tran (cddip0_out_im_config[6], \cddip0_out_im_config.f.wr_credit_config [6]);
tran (cddip0_out_im_config[5], \cddip0_out_im_config.r.part0 [5]);
tran (cddip0_out_im_config[5], \cddip0_out_im_config.f.wr_credit_config [5]);
tran (cddip0_out_im_config[4], \cddip0_out_im_config.r.part0 [4]);
tran (cddip0_out_im_config[4], \cddip0_out_im_config.f.wr_credit_config [4]);
tran (cddip0_out_im_config[3], \cddip0_out_im_config.r.part0 [3]);
tran (cddip0_out_im_config[3], \cddip0_out_im_config.f.wr_credit_config [3]);
tran (cddip0_out_im_config[2], \cddip0_out_im_config.r.part0 [2]);
tran (cddip0_out_im_config[2], \cddip0_out_im_config.f.wr_credit_config [2]);
tran (cddip0_out_im_config[1], \cddip0_out_im_config.r.part0 [1]);
tran (cddip0_out_im_config[1], \cddip0_out_im_config.f.wr_credit_config [1]);
tran (cddip0_out_im_config[0], \cddip0_out_im_config.r.part0 [0]);
tran (cddip0_out_im_config[0], \cddip0_out_im_config.f.wr_credit_config [0]);
tran (cddip1_out_ia_wdata[31], \cddip1_out_ia_wdata.r.part0 [31]);
tran (cddip1_out_ia_wdata[31], \cddip1_out_ia_wdata.f.eob );
tran (cddip1_out_ia_wdata[30], \cddip1_out_ia_wdata.r.part0 [30]);
tran (cddip1_out_ia_wdata[30], \cddip1_out_ia_wdata.f.bytes_vld [7]);
tran (cddip1_out_ia_wdata[29], \cddip1_out_ia_wdata.r.part0 [29]);
tran (cddip1_out_ia_wdata[29], \cddip1_out_ia_wdata.f.bytes_vld [6]);
tran (cddip1_out_ia_wdata[28], \cddip1_out_ia_wdata.r.part0 [28]);
tran (cddip1_out_ia_wdata[28], \cddip1_out_ia_wdata.f.bytes_vld [5]);
tran (cddip1_out_ia_wdata[27], \cddip1_out_ia_wdata.r.part0 [27]);
tran (cddip1_out_ia_wdata[27], \cddip1_out_ia_wdata.f.bytes_vld [4]);
tran (cddip1_out_ia_wdata[26], \cddip1_out_ia_wdata.r.part0 [26]);
tran (cddip1_out_ia_wdata[26], \cddip1_out_ia_wdata.f.bytes_vld [3]);
tran (cddip1_out_ia_wdata[25], \cddip1_out_ia_wdata.r.part0 [25]);
tran (cddip1_out_ia_wdata[25], \cddip1_out_ia_wdata.f.bytes_vld [2]);
tran (cddip1_out_ia_wdata[24], \cddip1_out_ia_wdata.r.part0 [24]);
tran (cddip1_out_ia_wdata[24], \cddip1_out_ia_wdata.f.bytes_vld [1]);
tran (cddip1_out_ia_wdata[23], \cddip1_out_ia_wdata.r.part0 [23]);
tran (cddip1_out_ia_wdata[23], \cddip1_out_ia_wdata.f.bytes_vld [0]);
tran (cddip1_out_ia_wdata[22], \cddip1_out_ia_wdata.r.part0 [22]);
tran (cddip1_out_ia_wdata[22], \cddip1_out_ia_wdata.f.unused1 [7]);
tran (cddip1_out_ia_wdata[21], \cddip1_out_ia_wdata.r.part0 [21]);
tran (cddip1_out_ia_wdata[21], \cddip1_out_ia_wdata.f.unused1 [6]);
tran (cddip1_out_ia_wdata[20], \cddip1_out_ia_wdata.r.part0 [20]);
tran (cddip1_out_ia_wdata[20], \cddip1_out_ia_wdata.f.unused1 [5]);
tran (cddip1_out_ia_wdata[19], \cddip1_out_ia_wdata.r.part0 [19]);
tran (cddip1_out_ia_wdata[19], \cddip1_out_ia_wdata.f.unused1 [4]);
tran (cddip1_out_ia_wdata[18], \cddip1_out_ia_wdata.r.part0 [18]);
tran (cddip1_out_ia_wdata[18], \cddip1_out_ia_wdata.f.unused1 [3]);
tran (cddip1_out_ia_wdata[17], \cddip1_out_ia_wdata.r.part0 [17]);
tran (cddip1_out_ia_wdata[17], \cddip1_out_ia_wdata.f.unused1 [2]);
tran (cddip1_out_ia_wdata[16], \cddip1_out_ia_wdata.r.part0 [16]);
tran (cddip1_out_ia_wdata[16], \cddip1_out_ia_wdata.f.unused1 [1]);
tran (cddip1_out_ia_wdata[15], \cddip1_out_ia_wdata.r.part0 [15]);
tran (cddip1_out_ia_wdata[15], \cddip1_out_ia_wdata.f.unused1 [0]);
tran (cddip1_out_ia_wdata[14], \cddip1_out_ia_wdata.r.part0 [14]);
tran (cddip1_out_ia_wdata[14], \cddip1_out_ia_wdata.f.tid );
tran (cddip1_out_ia_wdata[13], \cddip1_out_ia_wdata.r.part0 [13]);
tran (cddip1_out_ia_wdata[13], \cddip1_out_ia_wdata.f.tuser [7]);
tran (cddip1_out_ia_wdata[12], \cddip1_out_ia_wdata.r.part0 [12]);
tran (cddip1_out_ia_wdata[12], \cddip1_out_ia_wdata.f.tuser [6]);
tran (cddip1_out_ia_wdata[11], \cddip1_out_ia_wdata.r.part0 [11]);
tran (cddip1_out_ia_wdata[11], \cddip1_out_ia_wdata.f.tuser [5]);
tran (cddip1_out_ia_wdata[10], \cddip1_out_ia_wdata.r.part0 [10]);
tran (cddip1_out_ia_wdata[10], \cddip1_out_ia_wdata.f.tuser [4]);
tran (cddip1_out_ia_wdata[9], \cddip1_out_ia_wdata.r.part0 [9]);
tran (cddip1_out_ia_wdata[9], \cddip1_out_ia_wdata.f.tuser [3]);
tran (cddip1_out_ia_wdata[8], \cddip1_out_ia_wdata.r.part0 [8]);
tran (cddip1_out_ia_wdata[8], \cddip1_out_ia_wdata.f.tuser [2]);
tran (cddip1_out_ia_wdata[7], \cddip1_out_ia_wdata.r.part0 [7]);
tran (cddip1_out_ia_wdata[7], \cddip1_out_ia_wdata.f.tuser [1]);
tran (cddip1_out_ia_wdata[6], \cddip1_out_ia_wdata.r.part0 [6]);
tran (cddip1_out_ia_wdata[6], \cddip1_out_ia_wdata.f.tuser [0]);
tran (cddip1_out_ia_wdata[5], \cddip1_out_ia_wdata.r.part0 [5]);
tran (cddip1_out_ia_wdata[5], \cddip1_out_ia_wdata.f.unused0 [5]);
tran (cddip1_out_ia_wdata[4], \cddip1_out_ia_wdata.r.part0 [4]);
tran (cddip1_out_ia_wdata[4], \cddip1_out_ia_wdata.f.unused0 [4]);
tran (cddip1_out_ia_wdata[3], \cddip1_out_ia_wdata.r.part0 [3]);
tran (cddip1_out_ia_wdata[3], \cddip1_out_ia_wdata.f.unused0 [3]);
tran (cddip1_out_ia_wdata[2], \cddip1_out_ia_wdata.r.part0 [2]);
tran (cddip1_out_ia_wdata[2], \cddip1_out_ia_wdata.f.unused0 [2]);
tran (cddip1_out_ia_wdata[1], \cddip1_out_ia_wdata.r.part0 [1]);
tran (cddip1_out_ia_wdata[1], \cddip1_out_ia_wdata.f.unused0 [1]);
tran (cddip1_out_ia_wdata[0], \cddip1_out_ia_wdata.r.part0 [0]);
tran (cddip1_out_ia_wdata[0], \cddip1_out_ia_wdata.f.unused0 [0]);
tran (cddip1_out_ia_wdata[63], \cddip1_out_ia_wdata.r.part1 [31]);
tran (cddip1_out_ia_wdata[63], \cddip1_out_ia_wdata.f.tdata_lo [31]);
tran (cddip1_out_ia_wdata[62], \cddip1_out_ia_wdata.r.part1 [30]);
tran (cddip1_out_ia_wdata[62], \cddip1_out_ia_wdata.f.tdata_lo [30]);
tran (cddip1_out_ia_wdata[61], \cddip1_out_ia_wdata.r.part1 [29]);
tran (cddip1_out_ia_wdata[61], \cddip1_out_ia_wdata.f.tdata_lo [29]);
tran (cddip1_out_ia_wdata[60], \cddip1_out_ia_wdata.r.part1 [28]);
tran (cddip1_out_ia_wdata[60], \cddip1_out_ia_wdata.f.tdata_lo [28]);
tran (cddip1_out_ia_wdata[59], \cddip1_out_ia_wdata.r.part1 [27]);
tran (cddip1_out_ia_wdata[59], \cddip1_out_ia_wdata.f.tdata_lo [27]);
tran (cddip1_out_ia_wdata[58], \cddip1_out_ia_wdata.r.part1 [26]);
tran (cddip1_out_ia_wdata[58], \cddip1_out_ia_wdata.f.tdata_lo [26]);
tran (cddip1_out_ia_wdata[57], \cddip1_out_ia_wdata.r.part1 [25]);
tran (cddip1_out_ia_wdata[57], \cddip1_out_ia_wdata.f.tdata_lo [25]);
tran (cddip1_out_ia_wdata[56], \cddip1_out_ia_wdata.r.part1 [24]);
tran (cddip1_out_ia_wdata[56], \cddip1_out_ia_wdata.f.tdata_lo [24]);
tran (cddip1_out_ia_wdata[55], \cddip1_out_ia_wdata.r.part1 [23]);
tran (cddip1_out_ia_wdata[55], \cddip1_out_ia_wdata.f.tdata_lo [23]);
tran (cddip1_out_ia_wdata[54], \cddip1_out_ia_wdata.r.part1 [22]);
tran (cddip1_out_ia_wdata[54], \cddip1_out_ia_wdata.f.tdata_lo [22]);
tran (cddip1_out_ia_wdata[53], \cddip1_out_ia_wdata.r.part1 [21]);
tran (cddip1_out_ia_wdata[53], \cddip1_out_ia_wdata.f.tdata_lo [21]);
tran (cddip1_out_ia_wdata[52], \cddip1_out_ia_wdata.r.part1 [20]);
tran (cddip1_out_ia_wdata[52], \cddip1_out_ia_wdata.f.tdata_lo [20]);
tran (cddip1_out_ia_wdata[51], \cddip1_out_ia_wdata.r.part1 [19]);
tran (cddip1_out_ia_wdata[51], \cddip1_out_ia_wdata.f.tdata_lo [19]);
tran (cddip1_out_ia_wdata[50], \cddip1_out_ia_wdata.r.part1 [18]);
tran (cddip1_out_ia_wdata[50], \cddip1_out_ia_wdata.f.tdata_lo [18]);
tran (cddip1_out_ia_wdata[49], \cddip1_out_ia_wdata.r.part1 [17]);
tran (cddip1_out_ia_wdata[49], \cddip1_out_ia_wdata.f.tdata_lo [17]);
tran (cddip1_out_ia_wdata[48], \cddip1_out_ia_wdata.r.part1 [16]);
tran (cddip1_out_ia_wdata[48], \cddip1_out_ia_wdata.f.tdata_lo [16]);
tran (cddip1_out_ia_wdata[47], \cddip1_out_ia_wdata.r.part1 [15]);
tran (cddip1_out_ia_wdata[47], \cddip1_out_ia_wdata.f.tdata_lo [15]);
tran (cddip1_out_ia_wdata[46], \cddip1_out_ia_wdata.r.part1 [14]);
tran (cddip1_out_ia_wdata[46], \cddip1_out_ia_wdata.f.tdata_lo [14]);
tran (cddip1_out_ia_wdata[45], \cddip1_out_ia_wdata.r.part1 [13]);
tran (cddip1_out_ia_wdata[45], \cddip1_out_ia_wdata.f.tdata_lo [13]);
tran (cddip1_out_ia_wdata[44], \cddip1_out_ia_wdata.r.part1 [12]);
tran (cddip1_out_ia_wdata[44], \cddip1_out_ia_wdata.f.tdata_lo [12]);
tran (cddip1_out_ia_wdata[43], \cddip1_out_ia_wdata.r.part1 [11]);
tran (cddip1_out_ia_wdata[43], \cddip1_out_ia_wdata.f.tdata_lo [11]);
tran (cddip1_out_ia_wdata[42], \cddip1_out_ia_wdata.r.part1 [10]);
tran (cddip1_out_ia_wdata[42], \cddip1_out_ia_wdata.f.tdata_lo [10]);
tran (cddip1_out_ia_wdata[41], \cddip1_out_ia_wdata.r.part1 [9]);
tran (cddip1_out_ia_wdata[41], \cddip1_out_ia_wdata.f.tdata_lo [9]);
tran (cddip1_out_ia_wdata[40], \cddip1_out_ia_wdata.r.part1 [8]);
tran (cddip1_out_ia_wdata[40], \cddip1_out_ia_wdata.f.tdata_lo [8]);
tran (cddip1_out_ia_wdata[39], \cddip1_out_ia_wdata.r.part1 [7]);
tran (cddip1_out_ia_wdata[39], \cddip1_out_ia_wdata.f.tdata_lo [7]);
tran (cddip1_out_ia_wdata[38], \cddip1_out_ia_wdata.r.part1 [6]);
tran (cddip1_out_ia_wdata[38], \cddip1_out_ia_wdata.f.tdata_lo [6]);
tran (cddip1_out_ia_wdata[37], \cddip1_out_ia_wdata.r.part1 [5]);
tran (cddip1_out_ia_wdata[37], \cddip1_out_ia_wdata.f.tdata_lo [5]);
tran (cddip1_out_ia_wdata[36], \cddip1_out_ia_wdata.r.part1 [4]);
tran (cddip1_out_ia_wdata[36], \cddip1_out_ia_wdata.f.tdata_lo [4]);
tran (cddip1_out_ia_wdata[35], \cddip1_out_ia_wdata.r.part1 [3]);
tran (cddip1_out_ia_wdata[35], \cddip1_out_ia_wdata.f.tdata_lo [3]);
tran (cddip1_out_ia_wdata[34], \cddip1_out_ia_wdata.r.part1 [2]);
tran (cddip1_out_ia_wdata[34], \cddip1_out_ia_wdata.f.tdata_lo [2]);
tran (cddip1_out_ia_wdata[33], \cddip1_out_ia_wdata.r.part1 [1]);
tran (cddip1_out_ia_wdata[33], \cddip1_out_ia_wdata.f.tdata_lo [1]);
tran (cddip1_out_ia_wdata[32], \cddip1_out_ia_wdata.r.part1 [0]);
tran (cddip1_out_ia_wdata[32], \cddip1_out_ia_wdata.f.tdata_lo [0]);
tran (cddip1_out_ia_wdata[95], \cddip1_out_ia_wdata.r.part2 [31]);
tran (cddip1_out_ia_wdata[95], \cddip1_out_ia_wdata.f.tdata_hi [31]);
tran (cddip1_out_ia_wdata[94], \cddip1_out_ia_wdata.r.part2 [30]);
tran (cddip1_out_ia_wdata[94], \cddip1_out_ia_wdata.f.tdata_hi [30]);
tran (cddip1_out_ia_wdata[93], \cddip1_out_ia_wdata.r.part2 [29]);
tran (cddip1_out_ia_wdata[93], \cddip1_out_ia_wdata.f.tdata_hi [29]);
tran (cddip1_out_ia_wdata[92], \cddip1_out_ia_wdata.r.part2 [28]);
tran (cddip1_out_ia_wdata[92], \cddip1_out_ia_wdata.f.tdata_hi [28]);
tran (cddip1_out_ia_wdata[91], \cddip1_out_ia_wdata.r.part2 [27]);
tran (cddip1_out_ia_wdata[91], \cddip1_out_ia_wdata.f.tdata_hi [27]);
tran (cddip1_out_ia_wdata[90], \cddip1_out_ia_wdata.r.part2 [26]);
tran (cddip1_out_ia_wdata[90], \cddip1_out_ia_wdata.f.tdata_hi [26]);
tran (cddip1_out_ia_wdata[89], \cddip1_out_ia_wdata.r.part2 [25]);
tran (cddip1_out_ia_wdata[89], \cddip1_out_ia_wdata.f.tdata_hi [25]);
tran (cddip1_out_ia_wdata[88], \cddip1_out_ia_wdata.r.part2 [24]);
tran (cddip1_out_ia_wdata[88], \cddip1_out_ia_wdata.f.tdata_hi [24]);
tran (cddip1_out_ia_wdata[87], \cddip1_out_ia_wdata.r.part2 [23]);
tran (cddip1_out_ia_wdata[87], \cddip1_out_ia_wdata.f.tdata_hi [23]);
tran (cddip1_out_ia_wdata[86], \cddip1_out_ia_wdata.r.part2 [22]);
tran (cddip1_out_ia_wdata[86], \cddip1_out_ia_wdata.f.tdata_hi [22]);
tran (cddip1_out_ia_wdata[85], \cddip1_out_ia_wdata.r.part2 [21]);
tran (cddip1_out_ia_wdata[85], \cddip1_out_ia_wdata.f.tdata_hi [21]);
tran (cddip1_out_ia_wdata[84], \cddip1_out_ia_wdata.r.part2 [20]);
tran (cddip1_out_ia_wdata[84], \cddip1_out_ia_wdata.f.tdata_hi [20]);
tran (cddip1_out_ia_wdata[83], \cddip1_out_ia_wdata.r.part2 [19]);
tran (cddip1_out_ia_wdata[83], \cddip1_out_ia_wdata.f.tdata_hi [19]);
tran (cddip1_out_ia_wdata[82], \cddip1_out_ia_wdata.r.part2 [18]);
tran (cddip1_out_ia_wdata[82], \cddip1_out_ia_wdata.f.tdata_hi [18]);
tran (cddip1_out_ia_wdata[81], \cddip1_out_ia_wdata.r.part2 [17]);
tran (cddip1_out_ia_wdata[81], \cddip1_out_ia_wdata.f.tdata_hi [17]);
tran (cddip1_out_ia_wdata[80], \cddip1_out_ia_wdata.r.part2 [16]);
tran (cddip1_out_ia_wdata[80], \cddip1_out_ia_wdata.f.tdata_hi [16]);
tran (cddip1_out_ia_wdata[79], \cddip1_out_ia_wdata.r.part2 [15]);
tran (cddip1_out_ia_wdata[79], \cddip1_out_ia_wdata.f.tdata_hi [15]);
tran (cddip1_out_ia_wdata[78], \cddip1_out_ia_wdata.r.part2 [14]);
tran (cddip1_out_ia_wdata[78], \cddip1_out_ia_wdata.f.tdata_hi [14]);
tran (cddip1_out_ia_wdata[77], \cddip1_out_ia_wdata.r.part2 [13]);
tran (cddip1_out_ia_wdata[77], \cddip1_out_ia_wdata.f.tdata_hi [13]);
tran (cddip1_out_ia_wdata[76], \cddip1_out_ia_wdata.r.part2 [12]);
tran (cddip1_out_ia_wdata[76], \cddip1_out_ia_wdata.f.tdata_hi [12]);
tran (cddip1_out_ia_wdata[75], \cddip1_out_ia_wdata.r.part2 [11]);
tran (cddip1_out_ia_wdata[75], \cddip1_out_ia_wdata.f.tdata_hi [11]);
tran (cddip1_out_ia_wdata[74], \cddip1_out_ia_wdata.r.part2 [10]);
tran (cddip1_out_ia_wdata[74], \cddip1_out_ia_wdata.f.tdata_hi [10]);
tran (cddip1_out_ia_wdata[73], \cddip1_out_ia_wdata.r.part2 [9]);
tran (cddip1_out_ia_wdata[73], \cddip1_out_ia_wdata.f.tdata_hi [9]);
tran (cddip1_out_ia_wdata[72], \cddip1_out_ia_wdata.r.part2 [8]);
tran (cddip1_out_ia_wdata[72], \cddip1_out_ia_wdata.f.tdata_hi [8]);
tran (cddip1_out_ia_wdata[71], \cddip1_out_ia_wdata.r.part2 [7]);
tran (cddip1_out_ia_wdata[71], \cddip1_out_ia_wdata.f.tdata_hi [7]);
tran (cddip1_out_ia_wdata[70], \cddip1_out_ia_wdata.r.part2 [6]);
tran (cddip1_out_ia_wdata[70], \cddip1_out_ia_wdata.f.tdata_hi [6]);
tran (cddip1_out_ia_wdata[69], \cddip1_out_ia_wdata.r.part2 [5]);
tran (cddip1_out_ia_wdata[69], \cddip1_out_ia_wdata.f.tdata_hi [5]);
tran (cddip1_out_ia_wdata[68], \cddip1_out_ia_wdata.r.part2 [4]);
tran (cddip1_out_ia_wdata[68], \cddip1_out_ia_wdata.f.tdata_hi [4]);
tran (cddip1_out_ia_wdata[67], \cddip1_out_ia_wdata.r.part2 [3]);
tran (cddip1_out_ia_wdata[67], \cddip1_out_ia_wdata.f.tdata_hi [3]);
tran (cddip1_out_ia_wdata[66], \cddip1_out_ia_wdata.r.part2 [2]);
tran (cddip1_out_ia_wdata[66], \cddip1_out_ia_wdata.f.tdata_hi [2]);
tran (cddip1_out_ia_wdata[65], \cddip1_out_ia_wdata.r.part2 [1]);
tran (cddip1_out_ia_wdata[65], \cddip1_out_ia_wdata.f.tdata_hi [1]);
tran (cddip1_out_ia_wdata[64], \cddip1_out_ia_wdata.r.part2 [0]);
tran (cddip1_out_ia_wdata[64], \cddip1_out_ia_wdata.f.tdata_hi [0]);
tran (cddip1_out_ia_config[12], \cddip1_out_ia_config.r.part0 [12]);
tran (cddip1_out_ia_config[12], \cddip1_out_ia_config.f.op [3]);
tran (cddip1_out_ia_config[11], \cddip1_out_ia_config.r.part0 [11]);
tran (cddip1_out_ia_config[11], \cddip1_out_ia_config.f.op [2]);
tran (cddip1_out_ia_config[10], \cddip1_out_ia_config.r.part0 [10]);
tran (cddip1_out_ia_config[10], \cddip1_out_ia_config.f.op [1]);
tran (cddip1_out_ia_config[9], \cddip1_out_ia_config.r.part0 [9]);
tran (cddip1_out_ia_config[9], \cddip1_out_ia_config.f.op [0]);
tran (cddip1_out_ia_config[8], \cddip1_out_ia_config.r.part0 [8]);
tran (cddip1_out_ia_config[8], \cddip1_out_ia_config.f.addr [8]);
tran (cddip1_out_ia_config[7], \cddip1_out_ia_config.r.part0 [7]);
tran (cddip1_out_ia_config[7], \cddip1_out_ia_config.f.addr [7]);
tran (cddip1_out_ia_config[6], \cddip1_out_ia_config.r.part0 [6]);
tran (cddip1_out_ia_config[6], \cddip1_out_ia_config.f.addr [6]);
tran (cddip1_out_ia_config[5], \cddip1_out_ia_config.r.part0 [5]);
tran (cddip1_out_ia_config[5], \cddip1_out_ia_config.f.addr [5]);
tran (cddip1_out_ia_config[4], \cddip1_out_ia_config.r.part0 [4]);
tran (cddip1_out_ia_config[4], \cddip1_out_ia_config.f.addr [4]);
tran (cddip1_out_ia_config[3], \cddip1_out_ia_config.r.part0 [3]);
tran (cddip1_out_ia_config[3], \cddip1_out_ia_config.f.addr [3]);
tran (cddip1_out_ia_config[2], \cddip1_out_ia_config.r.part0 [2]);
tran (cddip1_out_ia_config[2], \cddip1_out_ia_config.f.addr [2]);
tran (cddip1_out_ia_config[1], \cddip1_out_ia_config.r.part0 [1]);
tran (cddip1_out_ia_config[1], \cddip1_out_ia_config.f.addr [1]);
tran (cddip1_out_ia_config[0], \cddip1_out_ia_config.r.part0 [0]);
tran (cddip1_out_ia_config[0], \cddip1_out_ia_config.f.addr [0]);
tran (cddip1_out_im_config[11], \cddip1_out_im_config.r.part0 [11]);
tran (cddip1_out_im_config[11], \cddip1_out_im_config.f.mode [1]);
tran (cddip1_out_im_config[10], \cddip1_out_im_config.r.part0 [10]);
tran (cddip1_out_im_config[10], \cddip1_out_im_config.f.mode [0]);
tran (cddip1_out_im_config[9], \cddip1_out_im_config.r.part0 [9]);
tran (cddip1_out_im_config[9], \cddip1_out_im_config.f.wr_credit_config [9]);
tran (cddip1_out_im_config[8], \cddip1_out_im_config.r.part0 [8]);
tran (cddip1_out_im_config[8], \cddip1_out_im_config.f.wr_credit_config [8]);
tran (cddip1_out_im_config[7], \cddip1_out_im_config.r.part0 [7]);
tran (cddip1_out_im_config[7], \cddip1_out_im_config.f.wr_credit_config [7]);
tran (cddip1_out_im_config[6], \cddip1_out_im_config.r.part0 [6]);
tran (cddip1_out_im_config[6], \cddip1_out_im_config.f.wr_credit_config [6]);
tran (cddip1_out_im_config[5], \cddip1_out_im_config.r.part0 [5]);
tran (cddip1_out_im_config[5], \cddip1_out_im_config.f.wr_credit_config [5]);
tran (cddip1_out_im_config[4], \cddip1_out_im_config.r.part0 [4]);
tran (cddip1_out_im_config[4], \cddip1_out_im_config.f.wr_credit_config [4]);
tran (cddip1_out_im_config[3], \cddip1_out_im_config.r.part0 [3]);
tran (cddip1_out_im_config[3], \cddip1_out_im_config.f.wr_credit_config [3]);
tran (cddip1_out_im_config[2], \cddip1_out_im_config.r.part0 [2]);
tran (cddip1_out_im_config[2], \cddip1_out_im_config.f.wr_credit_config [2]);
tran (cddip1_out_im_config[1], \cddip1_out_im_config.r.part0 [1]);
tran (cddip1_out_im_config[1], \cddip1_out_im_config.f.wr_credit_config [1]);
tran (cddip1_out_im_config[0], \cddip1_out_im_config.r.part0 [0]);
tran (cddip1_out_im_config[0], \cddip1_out_im_config.f.wr_credit_config [0]);
tran (cddip2_out_ia_wdata[31], \cddip2_out_ia_wdata.r.part0 [31]);
tran (cddip2_out_ia_wdata[31], \cddip2_out_ia_wdata.f.eob );
tran (cddip2_out_ia_wdata[30], \cddip2_out_ia_wdata.r.part0 [30]);
tran (cddip2_out_ia_wdata[30], \cddip2_out_ia_wdata.f.bytes_vld [7]);
tran (cddip2_out_ia_wdata[29], \cddip2_out_ia_wdata.r.part0 [29]);
tran (cddip2_out_ia_wdata[29], \cddip2_out_ia_wdata.f.bytes_vld [6]);
tran (cddip2_out_ia_wdata[28], \cddip2_out_ia_wdata.r.part0 [28]);
tran (cddip2_out_ia_wdata[28], \cddip2_out_ia_wdata.f.bytes_vld [5]);
tran (cddip2_out_ia_wdata[27], \cddip2_out_ia_wdata.r.part0 [27]);
tran (cddip2_out_ia_wdata[27], \cddip2_out_ia_wdata.f.bytes_vld [4]);
tran (cddip2_out_ia_wdata[26], \cddip2_out_ia_wdata.r.part0 [26]);
tran (cddip2_out_ia_wdata[26], \cddip2_out_ia_wdata.f.bytes_vld [3]);
tran (cddip2_out_ia_wdata[25], \cddip2_out_ia_wdata.r.part0 [25]);
tran (cddip2_out_ia_wdata[25], \cddip2_out_ia_wdata.f.bytes_vld [2]);
tran (cddip2_out_ia_wdata[24], \cddip2_out_ia_wdata.r.part0 [24]);
tran (cddip2_out_ia_wdata[24], \cddip2_out_ia_wdata.f.bytes_vld [1]);
tran (cddip2_out_ia_wdata[23], \cddip2_out_ia_wdata.r.part0 [23]);
tran (cddip2_out_ia_wdata[23], \cddip2_out_ia_wdata.f.bytes_vld [0]);
tran (cddip2_out_ia_wdata[22], \cddip2_out_ia_wdata.r.part0 [22]);
tran (cddip2_out_ia_wdata[22], \cddip2_out_ia_wdata.f.unused1 [7]);
tran (cddip2_out_ia_wdata[21], \cddip2_out_ia_wdata.r.part0 [21]);
tran (cddip2_out_ia_wdata[21], \cddip2_out_ia_wdata.f.unused1 [6]);
tran (cddip2_out_ia_wdata[20], \cddip2_out_ia_wdata.r.part0 [20]);
tran (cddip2_out_ia_wdata[20], \cddip2_out_ia_wdata.f.unused1 [5]);
tran (cddip2_out_ia_wdata[19], \cddip2_out_ia_wdata.r.part0 [19]);
tran (cddip2_out_ia_wdata[19], \cddip2_out_ia_wdata.f.unused1 [4]);
tran (cddip2_out_ia_wdata[18], \cddip2_out_ia_wdata.r.part0 [18]);
tran (cddip2_out_ia_wdata[18], \cddip2_out_ia_wdata.f.unused1 [3]);
tran (cddip2_out_ia_wdata[17], \cddip2_out_ia_wdata.r.part0 [17]);
tran (cddip2_out_ia_wdata[17], \cddip2_out_ia_wdata.f.unused1 [2]);
tran (cddip2_out_ia_wdata[16], \cddip2_out_ia_wdata.r.part0 [16]);
tran (cddip2_out_ia_wdata[16], \cddip2_out_ia_wdata.f.unused1 [1]);
tran (cddip2_out_ia_wdata[15], \cddip2_out_ia_wdata.r.part0 [15]);
tran (cddip2_out_ia_wdata[15], \cddip2_out_ia_wdata.f.unused1 [0]);
tran (cddip2_out_ia_wdata[14], \cddip2_out_ia_wdata.r.part0 [14]);
tran (cddip2_out_ia_wdata[14], \cddip2_out_ia_wdata.f.tid );
tran (cddip2_out_ia_wdata[13], \cddip2_out_ia_wdata.r.part0 [13]);
tran (cddip2_out_ia_wdata[13], \cddip2_out_ia_wdata.f.tuser [7]);
tran (cddip2_out_ia_wdata[12], \cddip2_out_ia_wdata.r.part0 [12]);
tran (cddip2_out_ia_wdata[12], \cddip2_out_ia_wdata.f.tuser [6]);
tran (cddip2_out_ia_wdata[11], \cddip2_out_ia_wdata.r.part0 [11]);
tran (cddip2_out_ia_wdata[11], \cddip2_out_ia_wdata.f.tuser [5]);
tran (cddip2_out_ia_wdata[10], \cddip2_out_ia_wdata.r.part0 [10]);
tran (cddip2_out_ia_wdata[10], \cddip2_out_ia_wdata.f.tuser [4]);
tran (cddip2_out_ia_wdata[9], \cddip2_out_ia_wdata.r.part0 [9]);
tran (cddip2_out_ia_wdata[9], \cddip2_out_ia_wdata.f.tuser [3]);
tran (cddip2_out_ia_wdata[8], \cddip2_out_ia_wdata.r.part0 [8]);
tran (cddip2_out_ia_wdata[8], \cddip2_out_ia_wdata.f.tuser [2]);
tran (cddip2_out_ia_wdata[7], \cddip2_out_ia_wdata.r.part0 [7]);
tran (cddip2_out_ia_wdata[7], \cddip2_out_ia_wdata.f.tuser [1]);
tran (cddip2_out_ia_wdata[6], \cddip2_out_ia_wdata.r.part0 [6]);
tran (cddip2_out_ia_wdata[6], \cddip2_out_ia_wdata.f.tuser [0]);
tran (cddip2_out_ia_wdata[5], \cddip2_out_ia_wdata.r.part0 [5]);
tran (cddip2_out_ia_wdata[5], \cddip2_out_ia_wdata.f.unused0 [5]);
tran (cddip2_out_ia_wdata[4], \cddip2_out_ia_wdata.r.part0 [4]);
tran (cddip2_out_ia_wdata[4], \cddip2_out_ia_wdata.f.unused0 [4]);
tran (cddip2_out_ia_wdata[3], \cddip2_out_ia_wdata.r.part0 [3]);
tran (cddip2_out_ia_wdata[3], \cddip2_out_ia_wdata.f.unused0 [3]);
tran (cddip2_out_ia_wdata[2], \cddip2_out_ia_wdata.r.part0 [2]);
tran (cddip2_out_ia_wdata[2], \cddip2_out_ia_wdata.f.unused0 [2]);
tran (cddip2_out_ia_wdata[1], \cddip2_out_ia_wdata.r.part0 [1]);
tran (cddip2_out_ia_wdata[1], \cddip2_out_ia_wdata.f.unused0 [1]);
tran (cddip2_out_ia_wdata[0], \cddip2_out_ia_wdata.r.part0 [0]);
tran (cddip2_out_ia_wdata[0], \cddip2_out_ia_wdata.f.unused0 [0]);
tran (cddip2_out_ia_wdata[63], \cddip2_out_ia_wdata.r.part1 [31]);
tran (cddip2_out_ia_wdata[63], \cddip2_out_ia_wdata.f.tdata_lo [31]);
tran (cddip2_out_ia_wdata[62], \cddip2_out_ia_wdata.r.part1 [30]);
tran (cddip2_out_ia_wdata[62], \cddip2_out_ia_wdata.f.tdata_lo [30]);
tran (cddip2_out_ia_wdata[61], \cddip2_out_ia_wdata.r.part1 [29]);
tran (cddip2_out_ia_wdata[61], \cddip2_out_ia_wdata.f.tdata_lo [29]);
tran (cddip2_out_ia_wdata[60], \cddip2_out_ia_wdata.r.part1 [28]);
tran (cddip2_out_ia_wdata[60], \cddip2_out_ia_wdata.f.tdata_lo [28]);
tran (cddip2_out_ia_wdata[59], \cddip2_out_ia_wdata.r.part1 [27]);
tran (cddip2_out_ia_wdata[59], \cddip2_out_ia_wdata.f.tdata_lo [27]);
tran (cddip2_out_ia_wdata[58], \cddip2_out_ia_wdata.r.part1 [26]);
tran (cddip2_out_ia_wdata[58], \cddip2_out_ia_wdata.f.tdata_lo [26]);
tran (cddip2_out_ia_wdata[57], \cddip2_out_ia_wdata.r.part1 [25]);
tran (cddip2_out_ia_wdata[57], \cddip2_out_ia_wdata.f.tdata_lo [25]);
tran (cddip2_out_ia_wdata[56], \cddip2_out_ia_wdata.r.part1 [24]);
tran (cddip2_out_ia_wdata[56], \cddip2_out_ia_wdata.f.tdata_lo [24]);
tran (cddip2_out_ia_wdata[55], \cddip2_out_ia_wdata.r.part1 [23]);
tran (cddip2_out_ia_wdata[55], \cddip2_out_ia_wdata.f.tdata_lo [23]);
tran (cddip2_out_ia_wdata[54], \cddip2_out_ia_wdata.r.part1 [22]);
tran (cddip2_out_ia_wdata[54], \cddip2_out_ia_wdata.f.tdata_lo [22]);
tran (cddip2_out_ia_wdata[53], \cddip2_out_ia_wdata.r.part1 [21]);
tran (cddip2_out_ia_wdata[53], \cddip2_out_ia_wdata.f.tdata_lo [21]);
tran (cddip2_out_ia_wdata[52], \cddip2_out_ia_wdata.r.part1 [20]);
tran (cddip2_out_ia_wdata[52], \cddip2_out_ia_wdata.f.tdata_lo [20]);
tran (cddip2_out_ia_wdata[51], \cddip2_out_ia_wdata.r.part1 [19]);
tran (cddip2_out_ia_wdata[51], \cddip2_out_ia_wdata.f.tdata_lo [19]);
tran (cddip2_out_ia_wdata[50], \cddip2_out_ia_wdata.r.part1 [18]);
tran (cddip2_out_ia_wdata[50], \cddip2_out_ia_wdata.f.tdata_lo [18]);
tran (cddip2_out_ia_wdata[49], \cddip2_out_ia_wdata.r.part1 [17]);
tran (cddip2_out_ia_wdata[49], \cddip2_out_ia_wdata.f.tdata_lo [17]);
tran (cddip2_out_ia_wdata[48], \cddip2_out_ia_wdata.r.part1 [16]);
tran (cddip2_out_ia_wdata[48], \cddip2_out_ia_wdata.f.tdata_lo [16]);
tran (cddip2_out_ia_wdata[47], \cddip2_out_ia_wdata.r.part1 [15]);
tran (cddip2_out_ia_wdata[47], \cddip2_out_ia_wdata.f.tdata_lo [15]);
tran (cddip2_out_ia_wdata[46], \cddip2_out_ia_wdata.r.part1 [14]);
tran (cddip2_out_ia_wdata[46], \cddip2_out_ia_wdata.f.tdata_lo [14]);
tran (cddip2_out_ia_wdata[45], \cddip2_out_ia_wdata.r.part1 [13]);
tran (cddip2_out_ia_wdata[45], \cddip2_out_ia_wdata.f.tdata_lo [13]);
tran (cddip2_out_ia_wdata[44], \cddip2_out_ia_wdata.r.part1 [12]);
tran (cddip2_out_ia_wdata[44], \cddip2_out_ia_wdata.f.tdata_lo [12]);
tran (cddip2_out_ia_wdata[43], \cddip2_out_ia_wdata.r.part1 [11]);
tran (cddip2_out_ia_wdata[43], \cddip2_out_ia_wdata.f.tdata_lo [11]);
tran (cddip2_out_ia_wdata[42], \cddip2_out_ia_wdata.r.part1 [10]);
tran (cddip2_out_ia_wdata[42], \cddip2_out_ia_wdata.f.tdata_lo [10]);
tran (cddip2_out_ia_wdata[41], \cddip2_out_ia_wdata.r.part1 [9]);
tran (cddip2_out_ia_wdata[41], \cddip2_out_ia_wdata.f.tdata_lo [9]);
tran (cddip2_out_ia_wdata[40], \cddip2_out_ia_wdata.r.part1 [8]);
tran (cddip2_out_ia_wdata[40], \cddip2_out_ia_wdata.f.tdata_lo [8]);
tran (cddip2_out_ia_wdata[39], \cddip2_out_ia_wdata.r.part1 [7]);
tran (cddip2_out_ia_wdata[39], \cddip2_out_ia_wdata.f.tdata_lo [7]);
tran (cddip2_out_ia_wdata[38], \cddip2_out_ia_wdata.r.part1 [6]);
tran (cddip2_out_ia_wdata[38], \cddip2_out_ia_wdata.f.tdata_lo [6]);
tran (cddip2_out_ia_wdata[37], \cddip2_out_ia_wdata.r.part1 [5]);
tran (cddip2_out_ia_wdata[37], \cddip2_out_ia_wdata.f.tdata_lo [5]);
tran (cddip2_out_ia_wdata[36], \cddip2_out_ia_wdata.r.part1 [4]);
tran (cddip2_out_ia_wdata[36], \cddip2_out_ia_wdata.f.tdata_lo [4]);
tran (cddip2_out_ia_wdata[35], \cddip2_out_ia_wdata.r.part1 [3]);
tran (cddip2_out_ia_wdata[35], \cddip2_out_ia_wdata.f.tdata_lo [3]);
tran (cddip2_out_ia_wdata[34], \cddip2_out_ia_wdata.r.part1 [2]);
tran (cddip2_out_ia_wdata[34], \cddip2_out_ia_wdata.f.tdata_lo [2]);
tran (cddip2_out_ia_wdata[33], \cddip2_out_ia_wdata.r.part1 [1]);
tran (cddip2_out_ia_wdata[33], \cddip2_out_ia_wdata.f.tdata_lo [1]);
tran (cddip2_out_ia_wdata[32], \cddip2_out_ia_wdata.r.part1 [0]);
tran (cddip2_out_ia_wdata[32], \cddip2_out_ia_wdata.f.tdata_lo [0]);
tran (cddip2_out_ia_wdata[95], \cddip2_out_ia_wdata.r.part2 [31]);
tran (cddip2_out_ia_wdata[95], \cddip2_out_ia_wdata.f.tdata_hi [31]);
tran (cddip2_out_ia_wdata[94], \cddip2_out_ia_wdata.r.part2 [30]);
tran (cddip2_out_ia_wdata[94], \cddip2_out_ia_wdata.f.tdata_hi [30]);
tran (cddip2_out_ia_wdata[93], \cddip2_out_ia_wdata.r.part2 [29]);
tran (cddip2_out_ia_wdata[93], \cddip2_out_ia_wdata.f.tdata_hi [29]);
tran (cddip2_out_ia_wdata[92], \cddip2_out_ia_wdata.r.part2 [28]);
tran (cddip2_out_ia_wdata[92], \cddip2_out_ia_wdata.f.tdata_hi [28]);
tran (cddip2_out_ia_wdata[91], \cddip2_out_ia_wdata.r.part2 [27]);
tran (cddip2_out_ia_wdata[91], \cddip2_out_ia_wdata.f.tdata_hi [27]);
tran (cddip2_out_ia_wdata[90], \cddip2_out_ia_wdata.r.part2 [26]);
tran (cddip2_out_ia_wdata[90], \cddip2_out_ia_wdata.f.tdata_hi [26]);
tran (cddip2_out_ia_wdata[89], \cddip2_out_ia_wdata.r.part2 [25]);
tran (cddip2_out_ia_wdata[89], \cddip2_out_ia_wdata.f.tdata_hi [25]);
tran (cddip2_out_ia_wdata[88], \cddip2_out_ia_wdata.r.part2 [24]);
tran (cddip2_out_ia_wdata[88], \cddip2_out_ia_wdata.f.tdata_hi [24]);
tran (cddip2_out_ia_wdata[87], \cddip2_out_ia_wdata.r.part2 [23]);
tran (cddip2_out_ia_wdata[87], \cddip2_out_ia_wdata.f.tdata_hi [23]);
tran (cddip2_out_ia_wdata[86], \cddip2_out_ia_wdata.r.part2 [22]);
tran (cddip2_out_ia_wdata[86], \cddip2_out_ia_wdata.f.tdata_hi [22]);
tran (cddip2_out_ia_wdata[85], \cddip2_out_ia_wdata.r.part2 [21]);
tran (cddip2_out_ia_wdata[85], \cddip2_out_ia_wdata.f.tdata_hi [21]);
tran (cddip2_out_ia_wdata[84], \cddip2_out_ia_wdata.r.part2 [20]);
tran (cddip2_out_ia_wdata[84], \cddip2_out_ia_wdata.f.tdata_hi [20]);
tran (cddip2_out_ia_wdata[83], \cddip2_out_ia_wdata.r.part2 [19]);
tran (cddip2_out_ia_wdata[83], \cddip2_out_ia_wdata.f.tdata_hi [19]);
tran (cddip2_out_ia_wdata[82], \cddip2_out_ia_wdata.r.part2 [18]);
tran (cddip2_out_ia_wdata[82], \cddip2_out_ia_wdata.f.tdata_hi [18]);
tran (cddip2_out_ia_wdata[81], \cddip2_out_ia_wdata.r.part2 [17]);
tran (cddip2_out_ia_wdata[81], \cddip2_out_ia_wdata.f.tdata_hi [17]);
tran (cddip2_out_ia_wdata[80], \cddip2_out_ia_wdata.r.part2 [16]);
tran (cddip2_out_ia_wdata[80], \cddip2_out_ia_wdata.f.tdata_hi [16]);
tran (cddip2_out_ia_wdata[79], \cddip2_out_ia_wdata.r.part2 [15]);
tran (cddip2_out_ia_wdata[79], \cddip2_out_ia_wdata.f.tdata_hi [15]);
tran (cddip2_out_ia_wdata[78], \cddip2_out_ia_wdata.r.part2 [14]);
tran (cddip2_out_ia_wdata[78], \cddip2_out_ia_wdata.f.tdata_hi [14]);
tran (cddip2_out_ia_wdata[77], \cddip2_out_ia_wdata.r.part2 [13]);
tran (cddip2_out_ia_wdata[77], \cddip2_out_ia_wdata.f.tdata_hi [13]);
tran (cddip2_out_ia_wdata[76], \cddip2_out_ia_wdata.r.part2 [12]);
tran (cddip2_out_ia_wdata[76], \cddip2_out_ia_wdata.f.tdata_hi [12]);
tran (cddip2_out_ia_wdata[75], \cddip2_out_ia_wdata.r.part2 [11]);
tran (cddip2_out_ia_wdata[75], \cddip2_out_ia_wdata.f.tdata_hi [11]);
tran (cddip2_out_ia_wdata[74], \cddip2_out_ia_wdata.r.part2 [10]);
tran (cddip2_out_ia_wdata[74], \cddip2_out_ia_wdata.f.tdata_hi [10]);
tran (cddip2_out_ia_wdata[73], \cddip2_out_ia_wdata.r.part2 [9]);
tran (cddip2_out_ia_wdata[73], \cddip2_out_ia_wdata.f.tdata_hi [9]);
tran (cddip2_out_ia_wdata[72], \cddip2_out_ia_wdata.r.part2 [8]);
tran (cddip2_out_ia_wdata[72], \cddip2_out_ia_wdata.f.tdata_hi [8]);
tran (cddip2_out_ia_wdata[71], \cddip2_out_ia_wdata.r.part2 [7]);
tran (cddip2_out_ia_wdata[71], \cddip2_out_ia_wdata.f.tdata_hi [7]);
tran (cddip2_out_ia_wdata[70], \cddip2_out_ia_wdata.r.part2 [6]);
tran (cddip2_out_ia_wdata[70], \cddip2_out_ia_wdata.f.tdata_hi [6]);
tran (cddip2_out_ia_wdata[69], \cddip2_out_ia_wdata.r.part2 [5]);
tran (cddip2_out_ia_wdata[69], \cddip2_out_ia_wdata.f.tdata_hi [5]);
tran (cddip2_out_ia_wdata[68], \cddip2_out_ia_wdata.r.part2 [4]);
tran (cddip2_out_ia_wdata[68], \cddip2_out_ia_wdata.f.tdata_hi [4]);
tran (cddip2_out_ia_wdata[67], \cddip2_out_ia_wdata.r.part2 [3]);
tran (cddip2_out_ia_wdata[67], \cddip2_out_ia_wdata.f.tdata_hi [3]);
tran (cddip2_out_ia_wdata[66], \cddip2_out_ia_wdata.r.part2 [2]);
tran (cddip2_out_ia_wdata[66], \cddip2_out_ia_wdata.f.tdata_hi [2]);
tran (cddip2_out_ia_wdata[65], \cddip2_out_ia_wdata.r.part2 [1]);
tran (cddip2_out_ia_wdata[65], \cddip2_out_ia_wdata.f.tdata_hi [1]);
tran (cddip2_out_ia_wdata[64], \cddip2_out_ia_wdata.r.part2 [0]);
tran (cddip2_out_ia_wdata[64], \cddip2_out_ia_wdata.f.tdata_hi [0]);
tran (cddip2_out_ia_config[12], \cddip2_out_ia_config.r.part0 [12]);
tran (cddip2_out_ia_config[12], \cddip2_out_ia_config.f.op [3]);
tran (cddip2_out_ia_config[11], \cddip2_out_ia_config.r.part0 [11]);
tran (cddip2_out_ia_config[11], \cddip2_out_ia_config.f.op [2]);
tran (cddip2_out_ia_config[10], \cddip2_out_ia_config.r.part0 [10]);
tran (cddip2_out_ia_config[10], \cddip2_out_ia_config.f.op [1]);
tran (cddip2_out_ia_config[9], \cddip2_out_ia_config.r.part0 [9]);
tran (cddip2_out_ia_config[9], \cddip2_out_ia_config.f.op [0]);
tran (cddip2_out_ia_config[8], \cddip2_out_ia_config.r.part0 [8]);
tran (cddip2_out_ia_config[8], \cddip2_out_ia_config.f.addr [8]);
tran (cddip2_out_ia_config[7], \cddip2_out_ia_config.r.part0 [7]);
tran (cddip2_out_ia_config[7], \cddip2_out_ia_config.f.addr [7]);
tran (cddip2_out_ia_config[6], \cddip2_out_ia_config.r.part0 [6]);
tran (cddip2_out_ia_config[6], \cddip2_out_ia_config.f.addr [6]);
tran (cddip2_out_ia_config[5], \cddip2_out_ia_config.r.part0 [5]);
tran (cddip2_out_ia_config[5], \cddip2_out_ia_config.f.addr [5]);
tran (cddip2_out_ia_config[4], \cddip2_out_ia_config.r.part0 [4]);
tran (cddip2_out_ia_config[4], \cddip2_out_ia_config.f.addr [4]);
tran (cddip2_out_ia_config[3], \cddip2_out_ia_config.r.part0 [3]);
tran (cddip2_out_ia_config[3], \cddip2_out_ia_config.f.addr [3]);
tran (cddip2_out_ia_config[2], \cddip2_out_ia_config.r.part0 [2]);
tran (cddip2_out_ia_config[2], \cddip2_out_ia_config.f.addr [2]);
tran (cddip2_out_ia_config[1], \cddip2_out_ia_config.r.part0 [1]);
tran (cddip2_out_ia_config[1], \cddip2_out_ia_config.f.addr [1]);
tran (cddip2_out_ia_config[0], \cddip2_out_ia_config.r.part0 [0]);
tran (cddip2_out_ia_config[0], \cddip2_out_ia_config.f.addr [0]);
tran (cddip2_out_im_config[11], \cddip2_out_im_config.r.part0 [11]);
tran (cddip2_out_im_config[11], \cddip2_out_im_config.f.mode [1]);
tran (cddip2_out_im_config[10], \cddip2_out_im_config.r.part0 [10]);
tran (cddip2_out_im_config[10], \cddip2_out_im_config.f.mode [0]);
tran (cddip2_out_im_config[9], \cddip2_out_im_config.r.part0 [9]);
tran (cddip2_out_im_config[9], \cddip2_out_im_config.f.wr_credit_config [9]);
tran (cddip2_out_im_config[8], \cddip2_out_im_config.r.part0 [8]);
tran (cddip2_out_im_config[8], \cddip2_out_im_config.f.wr_credit_config [8]);
tran (cddip2_out_im_config[7], \cddip2_out_im_config.r.part0 [7]);
tran (cddip2_out_im_config[7], \cddip2_out_im_config.f.wr_credit_config [7]);
tran (cddip2_out_im_config[6], \cddip2_out_im_config.r.part0 [6]);
tran (cddip2_out_im_config[6], \cddip2_out_im_config.f.wr_credit_config [6]);
tran (cddip2_out_im_config[5], \cddip2_out_im_config.r.part0 [5]);
tran (cddip2_out_im_config[5], \cddip2_out_im_config.f.wr_credit_config [5]);
tran (cddip2_out_im_config[4], \cddip2_out_im_config.r.part0 [4]);
tran (cddip2_out_im_config[4], \cddip2_out_im_config.f.wr_credit_config [4]);
tran (cddip2_out_im_config[3], \cddip2_out_im_config.r.part0 [3]);
tran (cddip2_out_im_config[3], \cddip2_out_im_config.f.wr_credit_config [3]);
tran (cddip2_out_im_config[2], \cddip2_out_im_config.r.part0 [2]);
tran (cddip2_out_im_config[2], \cddip2_out_im_config.f.wr_credit_config [2]);
tran (cddip2_out_im_config[1], \cddip2_out_im_config.r.part0 [1]);
tran (cddip2_out_im_config[1], \cddip2_out_im_config.f.wr_credit_config [1]);
tran (cddip2_out_im_config[0], \cddip2_out_im_config.r.part0 [0]);
tran (cddip2_out_im_config[0], \cddip2_out_im_config.f.wr_credit_config [0]);
tran (cddip3_out_ia_wdata[31], \cddip3_out_ia_wdata.r.part0 [31]);
tran (cddip3_out_ia_wdata[31], \cddip3_out_ia_wdata.f.eob );
tran (cddip3_out_ia_wdata[30], \cddip3_out_ia_wdata.r.part0 [30]);
tran (cddip3_out_ia_wdata[30], \cddip3_out_ia_wdata.f.bytes_vld [7]);
tran (cddip3_out_ia_wdata[29], \cddip3_out_ia_wdata.r.part0 [29]);
tran (cddip3_out_ia_wdata[29], \cddip3_out_ia_wdata.f.bytes_vld [6]);
tran (cddip3_out_ia_wdata[28], \cddip3_out_ia_wdata.r.part0 [28]);
tran (cddip3_out_ia_wdata[28], \cddip3_out_ia_wdata.f.bytes_vld [5]);
tran (cddip3_out_ia_wdata[27], \cddip3_out_ia_wdata.r.part0 [27]);
tran (cddip3_out_ia_wdata[27], \cddip3_out_ia_wdata.f.bytes_vld [4]);
tran (cddip3_out_ia_wdata[26], \cddip3_out_ia_wdata.r.part0 [26]);
tran (cddip3_out_ia_wdata[26], \cddip3_out_ia_wdata.f.bytes_vld [3]);
tran (cddip3_out_ia_wdata[25], \cddip3_out_ia_wdata.r.part0 [25]);
tran (cddip3_out_ia_wdata[25], \cddip3_out_ia_wdata.f.bytes_vld [2]);
tran (cddip3_out_ia_wdata[24], \cddip3_out_ia_wdata.r.part0 [24]);
tran (cddip3_out_ia_wdata[24], \cddip3_out_ia_wdata.f.bytes_vld [1]);
tran (cddip3_out_ia_wdata[23], \cddip3_out_ia_wdata.r.part0 [23]);
tran (cddip3_out_ia_wdata[23], \cddip3_out_ia_wdata.f.bytes_vld [0]);
tran (cddip3_out_ia_wdata[22], \cddip3_out_ia_wdata.r.part0 [22]);
tran (cddip3_out_ia_wdata[22], \cddip3_out_ia_wdata.f.unused1 [7]);
tran (cddip3_out_ia_wdata[21], \cddip3_out_ia_wdata.r.part0 [21]);
tran (cddip3_out_ia_wdata[21], \cddip3_out_ia_wdata.f.unused1 [6]);
tran (cddip3_out_ia_wdata[20], \cddip3_out_ia_wdata.r.part0 [20]);
tran (cddip3_out_ia_wdata[20], \cddip3_out_ia_wdata.f.unused1 [5]);
tran (cddip3_out_ia_wdata[19], \cddip3_out_ia_wdata.r.part0 [19]);
tran (cddip3_out_ia_wdata[19], \cddip3_out_ia_wdata.f.unused1 [4]);
tran (cddip3_out_ia_wdata[18], \cddip3_out_ia_wdata.r.part0 [18]);
tran (cddip3_out_ia_wdata[18], \cddip3_out_ia_wdata.f.unused1 [3]);
tran (cddip3_out_ia_wdata[17], \cddip3_out_ia_wdata.r.part0 [17]);
tran (cddip3_out_ia_wdata[17], \cddip3_out_ia_wdata.f.unused1 [2]);
tran (cddip3_out_ia_wdata[16], \cddip3_out_ia_wdata.r.part0 [16]);
tran (cddip3_out_ia_wdata[16], \cddip3_out_ia_wdata.f.unused1 [1]);
tran (cddip3_out_ia_wdata[15], \cddip3_out_ia_wdata.r.part0 [15]);
tran (cddip3_out_ia_wdata[15], \cddip3_out_ia_wdata.f.unused1 [0]);
tran (cddip3_out_ia_wdata[14], \cddip3_out_ia_wdata.r.part0 [14]);
tran (cddip3_out_ia_wdata[14], \cddip3_out_ia_wdata.f.tid );
tran (cddip3_out_ia_wdata[13], \cddip3_out_ia_wdata.r.part0 [13]);
tran (cddip3_out_ia_wdata[13], \cddip3_out_ia_wdata.f.tuser [7]);
tran (cddip3_out_ia_wdata[12], \cddip3_out_ia_wdata.r.part0 [12]);
tran (cddip3_out_ia_wdata[12], \cddip3_out_ia_wdata.f.tuser [6]);
tran (cddip3_out_ia_wdata[11], \cddip3_out_ia_wdata.r.part0 [11]);
tran (cddip3_out_ia_wdata[11], \cddip3_out_ia_wdata.f.tuser [5]);
tran (cddip3_out_ia_wdata[10], \cddip3_out_ia_wdata.r.part0 [10]);
tran (cddip3_out_ia_wdata[10], \cddip3_out_ia_wdata.f.tuser [4]);
tran (cddip3_out_ia_wdata[9], \cddip3_out_ia_wdata.r.part0 [9]);
tran (cddip3_out_ia_wdata[9], \cddip3_out_ia_wdata.f.tuser [3]);
tran (cddip3_out_ia_wdata[8], \cddip3_out_ia_wdata.r.part0 [8]);
tran (cddip3_out_ia_wdata[8], \cddip3_out_ia_wdata.f.tuser [2]);
tran (cddip3_out_ia_wdata[7], \cddip3_out_ia_wdata.r.part0 [7]);
tran (cddip3_out_ia_wdata[7], \cddip3_out_ia_wdata.f.tuser [1]);
tran (cddip3_out_ia_wdata[6], \cddip3_out_ia_wdata.r.part0 [6]);
tran (cddip3_out_ia_wdata[6], \cddip3_out_ia_wdata.f.tuser [0]);
tran (cddip3_out_ia_wdata[5], \cddip3_out_ia_wdata.r.part0 [5]);
tran (cddip3_out_ia_wdata[5], \cddip3_out_ia_wdata.f.unused0 [5]);
tran (cddip3_out_ia_wdata[4], \cddip3_out_ia_wdata.r.part0 [4]);
tran (cddip3_out_ia_wdata[4], \cddip3_out_ia_wdata.f.unused0 [4]);
tran (cddip3_out_ia_wdata[3], \cddip3_out_ia_wdata.r.part0 [3]);
tran (cddip3_out_ia_wdata[3], \cddip3_out_ia_wdata.f.unused0 [3]);
tran (cddip3_out_ia_wdata[2], \cddip3_out_ia_wdata.r.part0 [2]);
tran (cddip3_out_ia_wdata[2], \cddip3_out_ia_wdata.f.unused0 [2]);
tran (cddip3_out_ia_wdata[1], \cddip3_out_ia_wdata.r.part0 [1]);
tran (cddip3_out_ia_wdata[1], \cddip3_out_ia_wdata.f.unused0 [1]);
tran (cddip3_out_ia_wdata[0], \cddip3_out_ia_wdata.r.part0 [0]);
tran (cddip3_out_ia_wdata[0], \cddip3_out_ia_wdata.f.unused0 [0]);
tran (cddip3_out_ia_wdata[63], \cddip3_out_ia_wdata.r.part1 [31]);
tran (cddip3_out_ia_wdata[63], \cddip3_out_ia_wdata.f.tdata_lo [31]);
tran (cddip3_out_ia_wdata[62], \cddip3_out_ia_wdata.r.part1 [30]);
tran (cddip3_out_ia_wdata[62], \cddip3_out_ia_wdata.f.tdata_lo [30]);
tran (cddip3_out_ia_wdata[61], \cddip3_out_ia_wdata.r.part1 [29]);
tran (cddip3_out_ia_wdata[61], \cddip3_out_ia_wdata.f.tdata_lo [29]);
tran (cddip3_out_ia_wdata[60], \cddip3_out_ia_wdata.r.part1 [28]);
tran (cddip3_out_ia_wdata[60], \cddip3_out_ia_wdata.f.tdata_lo [28]);
tran (cddip3_out_ia_wdata[59], \cddip3_out_ia_wdata.r.part1 [27]);
tran (cddip3_out_ia_wdata[59], \cddip3_out_ia_wdata.f.tdata_lo [27]);
tran (cddip3_out_ia_wdata[58], \cddip3_out_ia_wdata.r.part1 [26]);
tran (cddip3_out_ia_wdata[58], \cddip3_out_ia_wdata.f.tdata_lo [26]);
tran (cddip3_out_ia_wdata[57], \cddip3_out_ia_wdata.r.part1 [25]);
tran (cddip3_out_ia_wdata[57], \cddip3_out_ia_wdata.f.tdata_lo [25]);
tran (cddip3_out_ia_wdata[56], \cddip3_out_ia_wdata.r.part1 [24]);
tran (cddip3_out_ia_wdata[56], \cddip3_out_ia_wdata.f.tdata_lo [24]);
tran (cddip3_out_ia_wdata[55], \cddip3_out_ia_wdata.r.part1 [23]);
tran (cddip3_out_ia_wdata[55], \cddip3_out_ia_wdata.f.tdata_lo [23]);
tran (cddip3_out_ia_wdata[54], \cddip3_out_ia_wdata.r.part1 [22]);
tran (cddip3_out_ia_wdata[54], \cddip3_out_ia_wdata.f.tdata_lo [22]);
tran (cddip3_out_ia_wdata[53], \cddip3_out_ia_wdata.r.part1 [21]);
tran (cddip3_out_ia_wdata[53], \cddip3_out_ia_wdata.f.tdata_lo [21]);
tran (cddip3_out_ia_wdata[52], \cddip3_out_ia_wdata.r.part1 [20]);
tran (cddip3_out_ia_wdata[52], \cddip3_out_ia_wdata.f.tdata_lo [20]);
tran (cddip3_out_ia_wdata[51], \cddip3_out_ia_wdata.r.part1 [19]);
tran (cddip3_out_ia_wdata[51], \cddip3_out_ia_wdata.f.tdata_lo [19]);
tran (cddip3_out_ia_wdata[50], \cddip3_out_ia_wdata.r.part1 [18]);
tran (cddip3_out_ia_wdata[50], \cddip3_out_ia_wdata.f.tdata_lo [18]);
tran (cddip3_out_ia_wdata[49], \cddip3_out_ia_wdata.r.part1 [17]);
tran (cddip3_out_ia_wdata[49], \cddip3_out_ia_wdata.f.tdata_lo [17]);
tran (cddip3_out_ia_wdata[48], \cddip3_out_ia_wdata.r.part1 [16]);
tran (cddip3_out_ia_wdata[48], \cddip3_out_ia_wdata.f.tdata_lo [16]);
tran (cddip3_out_ia_wdata[47], \cddip3_out_ia_wdata.r.part1 [15]);
tran (cddip3_out_ia_wdata[47], \cddip3_out_ia_wdata.f.tdata_lo [15]);
tran (cddip3_out_ia_wdata[46], \cddip3_out_ia_wdata.r.part1 [14]);
tran (cddip3_out_ia_wdata[46], \cddip3_out_ia_wdata.f.tdata_lo [14]);
tran (cddip3_out_ia_wdata[45], \cddip3_out_ia_wdata.r.part1 [13]);
tran (cddip3_out_ia_wdata[45], \cddip3_out_ia_wdata.f.tdata_lo [13]);
tran (cddip3_out_ia_wdata[44], \cddip3_out_ia_wdata.r.part1 [12]);
tran (cddip3_out_ia_wdata[44], \cddip3_out_ia_wdata.f.tdata_lo [12]);
tran (cddip3_out_ia_wdata[43], \cddip3_out_ia_wdata.r.part1 [11]);
tran (cddip3_out_ia_wdata[43], \cddip3_out_ia_wdata.f.tdata_lo [11]);
tran (cddip3_out_ia_wdata[42], \cddip3_out_ia_wdata.r.part1 [10]);
tran (cddip3_out_ia_wdata[42], \cddip3_out_ia_wdata.f.tdata_lo [10]);
tran (cddip3_out_ia_wdata[41], \cddip3_out_ia_wdata.r.part1 [9]);
tran (cddip3_out_ia_wdata[41], \cddip3_out_ia_wdata.f.tdata_lo [9]);
tran (cddip3_out_ia_wdata[40], \cddip3_out_ia_wdata.r.part1 [8]);
tran (cddip3_out_ia_wdata[40], \cddip3_out_ia_wdata.f.tdata_lo [8]);
tran (cddip3_out_ia_wdata[39], \cddip3_out_ia_wdata.r.part1 [7]);
tran (cddip3_out_ia_wdata[39], \cddip3_out_ia_wdata.f.tdata_lo [7]);
tran (cddip3_out_ia_wdata[38], \cddip3_out_ia_wdata.r.part1 [6]);
tran (cddip3_out_ia_wdata[38], \cddip3_out_ia_wdata.f.tdata_lo [6]);
tran (cddip3_out_ia_wdata[37], \cddip3_out_ia_wdata.r.part1 [5]);
tran (cddip3_out_ia_wdata[37], \cddip3_out_ia_wdata.f.tdata_lo [5]);
tran (cddip3_out_ia_wdata[36], \cddip3_out_ia_wdata.r.part1 [4]);
tran (cddip3_out_ia_wdata[36], \cddip3_out_ia_wdata.f.tdata_lo [4]);
tran (cddip3_out_ia_wdata[35], \cddip3_out_ia_wdata.r.part1 [3]);
tran (cddip3_out_ia_wdata[35], \cddip3_out_ia_wdata.f.tdata_lo [3]);
tran (cddip3_out_ia_wdata[34], \cddip3_out_ia_wdata.r.part1 [2]);
tran (cddip3_out_ia_wdata[34], \cddip3_out_ia_wdata.f.tdata_lo [2]);
tran (cddip3_out_ia_wdata[33], \cddip3_out_ia_wdata.r.part1 [1]);
tran (cddip3_out_ia_wdata[33], \cddip3_out_ia_wdata.f.tdata_lo [1]);
tran (cddip3_out_ia_wdata[32], \cddip3_out_ia_wdata.r.part1 [0]);
tran (cddip3_out_ia_wdata[32], \cddip3_out_ia_wdata.f.tdata_lo [0]);
tran (cddip3_out_ia_wdata[95], \cddip3_out_ia_wdata.r.part2 [31]);
tran (cddip3_out_ia_wdata[95], \cddip3_out_ia_wdata.f.tdata_hi [31]);
tran (cddip3_out_ia_wdata[94], \cddip3_out_ia_wdata.r.part2 [30]);
tran (cddip3_out_ia_wdata[94], \cddip3_out_ia_wdata.f.tdata_hi [30]);
tran (cddip3_out_ia_wdata[93], \cddip3_out_ia_wdata.r.part2 [29]);
tran (cddip3_out_ia_wdata[93], \cddip3_out_ia_wdata.f.tdata_hi [29]);
tran (cddip3_out_ia_wdata[92], \cddip3_out_ia_wdata.r.part2 [28]);
tran (cddip3_out_ia_wdata[92], \cddip3_out_ia_wdata.f.tdata_hi [28]);
tran (cddip3_out_ia_wdata[91], \cddip3_out_ia_wdata.r.part2 [27]);
tran (cddip3_out_ia_wdata[91], \cddip3_out_ia_wdata.f.tdata_hi [27]);
tran (cddip3_out_ia_wdata[90], \cddip3_out_ia_wdata.r.part2 [26]);
tran (cddip3_out_ia_wdata[90], \cddip3_out_ia_wdata.f.tdata_hi [26]);
tran (cddip3_out_ia_wdata[89], \cddip3_out_ia_wdata.r.part2 [25]);
tran (cddip3_out_ia_wdata[89], \cddip3_out_ia_wdata.f.tdata_hi [25]);
tran (cddip3_out_ia_wdata[88], \cddip3_out_ia_wdata.r.part2 [24]);
tran (cddip3_out_ia_wdata[88], \cddip3_out_ia_wdata.f.tdata_hi [24]);
tran (cddip3_out_ia_wdata[87], \cddip3_out_ia_wdata.r.part2 [23]);
tran (cddip3_out_ia_wdata[87], \cddip3_out_ia_wdata.f.tdata_hi [23]);
tran (cddip3_out_ia_wdata[86], \cddip3_out_ia_wdata.r.part2 [22]);
tran (cddip3_out_ia_wdata[86], \cddip3_out_ia_wdata.f.tdata_hi [22]);
tran (cddip3_out_ia_wdata[85], \cddip3_out_ia_wdata.r.part2 [21]);
tran (cddip3_out_ia_wdata[85], \cddip3_out_ia_wdata.f.tdata_hi [21]);
tran (cddip3_out_ia_wdata[84], \cddip3_out_ia_wdata.r.part2 [20]);
tran (cddip3_out_ia_wdata[84], \cddip3_out_ia_wdata.f.tdata_hi [20]);
tran (cddip3_out_ia_wdata[83], \cddip3_out_ia_wdata.r.part2 [19]);
tran (cddip3_out_ia_wdata[83], \cddip3_out_ia_wdata.f.tdata_hi [19]);
tran (cddip3_out_ia_wdata[82], \cddip3_out_ia_wdata.r.part2 [18]);
tran (cddip3_out_ia_wdata[82], \cddip3_out_ia_wdata.f.tdata_hi [18]);
tran (cddip3_out_ia_wdata[81], \cddip3_out_ia_wdata.r.part2 [17]);
tran (cddip3_out_ia_wdata[81], \cddip3_out_ia_wdata.f.tdata_hi [17]);
tran (cddip3_out_ia_wdata[80], \cddip3_out_ia_wdata.r.part2 [16]);
tran (cddip3_out_ia_wdata[80], \cddip3_out_ia_wdata.f.tdata_hi [16]);
tran (cddip3_out_ia_wdata[79], \cddip3_out_ia_wdata.r.part2 [15]);
tran (cddip3_out_ia_wdata[79], \cddip3_out_ia_wdata.f.tdata_hi [15]);
tran (cddip3_out_ia_wdata[78], \cddip3_out_ia_wdata.r.part2 [14]);
tran (cddip3_out_ia_wdata[78], \cddip3_out_ia_wdata.f.tdata_hi [14]);
tran (cddip3_out_ia_wdata[77], \cddip3_out_ia_wdata.r.part2 [13]);
tran (cddip3_out_ia_wdata[77], \cddip3_out_ia_wdata.f.tdata_hi [13]);
tran (cddip3_out_ia_wdata[76], \cddip3_out_ia_wdata.r.part2 [12]);
tran (cddip3_out_ia_wdata[76], \cddip3_out_ia_wdata.f.tdata_hi [12]);
tran (cddip3_out_ia_wdata[75], \cddip3_out_ia_wdata.r.part2 [11]);
tran (cddip3_out_ia_wdata[75], \cddip3_out_ia_wdata.f.tdata_hi [11]);
tran (cddip3_out_ia_wdata[74], \cddip3_out_ia_wdata.r.part2 [10]);
tran (cddip3_out_ia_wdata[74], \cddip3_out_ia_wdata.f.tdata_hi [10]);
tran (cddip3_out_ia_wdata[73], \cddip3_out_ia_wdata.r.part2 [9]);
tran (cddip3_out_ia_wdata[73], \cddip3_out_ia_wdata.f.tdata_hi [9]);
tran (cddip3_out_ia_wdata[72], \cddip3_out_ia_wdata.r.part2 [8]);
tran (cddip3_out_ia_wdata[72], \cddip3_out_ia_wdata.f.tdata_hi [8]);
tran (cddip3_out_ia_wdata[71], \cddip3_out_ia_wdata.r.part2 [7]);
tran (cddip3_out_ia_wdata[71], \cddip3_out_ia_wdata.f.tdata_hi [7]);
tran (cddip3_out_ia_wdata[70], \cddip3_out_ia_wdata.r.part2 [6]);
tran (cddip3_out_ia_wdata[70], \cddip3_out_ia_wdata.f.tdata_hi [6]);
tran (cddip3_out_ia_wdata[69], \cddip3_out_ia_wdata.r.part2 [5]);
tran (cddip3_out_ia_wdata[69], \cddip3_out_ia_wdata.f.tdata_hi [5]);
tran (cddip3_out_ia_wdata[68], \cddip3_out_ia_wdata.r.part2 [4]);
tran (cddip3_out_ia_wdata[68], \cddip3_out_ia_wdata.f.tdata_hi [4]);
tran (cddip3_out_ia_wdata[67], \cddip3_out_ia_wdata.r.part2 [3]);
tran (cddip3_out_ia_wdata[67], \cddip3_out_ia_wdata.f.tdata_hi [3]);
tran (cddip3_out_ia_wdata[66], \cddip3_out_ia_wdata.r.part2 [2]);
tran (cddip3_out_ia_wdata[66], \cddip3_out_ia_wdata.f.tdata_hi [2]);
tran (cddip3_out_ia_wdata[65], \cddip3_out_ia_wdata.r.part2 [1]);
tran (cddip3_out_ia_wdata[65], \cddip3_out_ia_wdata.f.tdata_hi [1]);
tran (cddip3_out_ia_wdata[64], \cddip3_out_ia_wdata.r.part2 [0]);
tran (cddip3_out_ia_wdata[64], \cddip3_out_ia_wdata.f.tdata_hi [0]);
tran (cddip3_out_ia_config[12], \cddip3_out_ia_config.r.part0 [12]);
tran (cddip3_out_ia_config[12], \cddip3_out_ia_config.f.op [3]);
tran (cddip3_out_ia_config[11], \cddip3_out_ia_config.r.part0 [11]);
tran (cddip3_out_ia_config[11], \cddip3_out_ia_config.f.op [2]);
tran (cddip3_out_ia_config[10], \cddip3_out_ia_config.r.part0 [10]);
tran (cddip3_out_ia_config[10], \cddip3_out_ia_config.f.op [1]);
tran (cddip3_out_ia_config[9], \cddip3_out_ia_config.r.part0 [9]);
tran (cddip3_out_ia_config[9], \cddip3_out_ia_config.f.op [0]);
tran (cddip3_out_ia_config[8], \cddip3_out_ia_config.r.part0 [8]);
tran (cddip3_out_ia_config[8], \cddip3_out_ia_config.f.addr [8]);
tran (cddip3_out_ia_config[7], \cddip3_out_ia_config.r.part0 [7]);
tran (cddip3_out_ia_config[7], \cddip3_out_ia_config.f.addr [7]);
tran (cddip3_out_ia_config[6], \cddip3_out_ia_config.r.part0 [6]);
tran (cddip3_out_ia_config[6], \cddip3_out_ia_config.f.addr [6]);
tran (cddip3_out_ia_config[5], \cddip3_out_ia_config.r.part0 [5]);
tran (cddip3_out_ia_config[5], \cddip3_out_ia_config.f.addr [5]);
tran (cddip3_out_ia_config[4], \cddip3_out_ia_config.r.part0 [4]);
tran (cddip3_out_ia_config[4], \cddip3_out_ia_config.f.addr [4]);
tran (cddip3_out_ia_config[3], \cddip3_out_ia_config.r.part0 [3]);
tran (cddip3_out_ia_config[3], \cddip3_out_ia_config.f.addr [3]);
tran (cddip3_out_ia_config[2], \cddip3_out_ia_config.r.part0 [2]);
tran (cddip3_out_ia_config[2], \cddip3_out_ia_config.f.addr [2]);
tran (cddip3_out_ia_config[1], \cddip3_out_ia_config.r.part0 [1]);
tran (cddip3_out_ia_config[1], \cddip3_out_ia_config.f.addr [1]);
tran (cddip3_out_ia_config[0], \cddip3_out_ia_config.r.part0 [0]);
tran (cddip3_out_ia_config[0], \cddip3_out_ia_config.f.addr [0]);
tran (cddip3_out_im_config[11], \cddip3_out_im_config.r.part0 [11]);
tran (cddip3_out_im_config[11], \cddip3_out_im_config.f.mode [1]);
tran (cddip3_out_im_config[10], \cddip3_out_im_config.r.part0 [10]);
tran (cddip3_out_im_config[10], \cddip3_out_im_config.f.mode [0]);
tran (cddip3_out_im_config[9], \cddip3_out_im_config.r.part0 [9]);
tran (cddip3_out_im_config[9], \cddip3_out_im_config.f.wr_credit_config [9]);
tran (cddip3_out_im_config[8], \cddip3_out_im_config.r.part0 [8]);
tran (cddip3_out_im_config[8], \cddip3_out_im_config.f.wr_credit_config [8]);
tran (cddip3_out_im_config[7], \cddip3_out_im_config.r.part0 [7]);
tran (cddip3_out_im_config[7], \cddip3_out_im_config.f.wr_credit_config [7]);
tran (cddip3_out_im_config[6], \cddip3_out_im_config.r.part0 [6]);
tran (cddip3_out_im_config[6], \cddip3_out_im_config.f.wr_credit_config [6]);
tran (cddip3_out_im_config[5], \cddip3_out_im_config.r.part0 [5]);
tran (cddip3_out_im_config[5], \cddip3_out_im_config.f.wr_credit_config [5]);
tran (cddip3_out_im_config[4], \cddip3_out_im_config.r.part0 [4]);
tran (cddip3_out_im_config[4], \cddip3_out_im_config.f.wr_credit_config [4]);
tran (cddip3_out_im_config[3], \cddip3_out_im_config.r.part0 [3]);
tran (cddip3_out_im_config[3], \cddip3_out_im_config.f.wr_credit_config [3]);
tran (cddip3_out_im_config[2], \cddip3_out_im_config.r.part0 [2]);
tran (cddip3_out_im_config[2], \cddip3_out_im_config.f.wr_credit_config [2]);
tran (cddip3_out_im_config[1], \cddip3_out_im_config.r.part0 [1]);
tran (cddip3_out_im_config[1], \cddip3_out_im_config.f.wr_credit_config [1]);
tran (cddip3_out_im_config[0], \cddip3_out_im_config.r.part0 [0]);
tran (cddip3_out_im_config[0], \cddip3_out_im_config.f.wr_credit_config [0]);
tran (sa_snapshot_ia_wdata[31], \sa_snapshot_ia_wdata.r.part0 [31]);
tran (sa_snapshot_ia_wdata[31], \sa_snapshot_ia_wdata.f.lower [31]);
tran (sa_snapshot_ia_wdata[30], \sa_snapshot_ia_wdata.r.part0 [30]);
tran (sa_snapshot_ia_wdata[30], \sa_snapshot_ia_wdata.f.lower [30]);
tran (sa_snapshot_ia_wdata[29], \sa_snapshot_ia_wdata.r.part0 [29]);
tran (sa_snapshot_ia_wdata[29], \sa_snapshot_ia_wdata.f.lower [29]);
tran (sa_snapshot_ia_wdata[28], \sa_snapshot_ia_wdata.r.part0 [28]);
tran (sa_snapshot_ia_wdata[28], \sa_snapshot_ia_wdata.f.lower [28]);
tran (sa_snapshot_ia_wdata[27], \sa_snapshot_ia_wdata.r.part0 [27]);
tran (sa_snapshot_ia_wdata[27], \sa_snapshot_ia_wdata.f.lower [27]);
tran (sa_snapshot_ia_wdata[26], \sa_snapshot_ia_wdata.r.part0 [26]);
tran (sa_snapshot_ia_wdata[26], \sa_snapshot_ia_wdata.f.lower [26]);
tran (sa_snapshot_ia_wdata[25], \sa_snapshot_ia_wdata.r.part0 [25]);
tran (sa_snapshot_ia_wdata[25], \sa_snapshot_ia_wdata.f.lower [25]);
tran (sa_snapshot_ia_wdata[24], \sa_snapshot_ia_wdata.r.part0 [24]);
tran (sa_snapshot_ia_wdata[24], \sa_snapshot_ia_wdata.f.lower [24]);
tran (sa_snapshot_ia_wdata[23], \sa_snapshot_ia_wdata.r.part0 [23]);
tran (sa_snapshot_ia_wdata[23], \sa_snapshot_ia_wdata.f.lower [23]);
tran (sa_snapshot_ia_wdata[22], \sa_snapshot_ia_wdata.r.part0 [22]);
tran (sa_snapshot_ia_wdata[22], \sa_snapshot_ia_wdata.f.lower [22]);
tran (sa_snapshot_ia_wdata[21], \sa_snapshot_ia_wdata.r.part0 [21]);
tran (sa_snapshot_ia_wdata[21], \sa_snapshot_ia_wdata.f.lower [21]);
tran (sa_snapshot_ia_wdata[20], \sa_snapshot_ia_wdata.r.part0 [20]);
tran (sa_snapshot_ia_wdata[20], \sa_snapshot_ia_wdata.f.lower [20]);
tran (sa_snapshot_ia_wdata[19], \sa_snapshot_ia_wdata.r.part0 [19]);
tran (sa_snapshot_ia_wdata[19], \sa_snapshot_ia_wdata.f.lower [19]);
tran (sa_snapshot_ia_wdata[18], \sa_snapshot_ia_wdata.r.part0 [18]);
tran (sa_snapshot_ia_wdata[18], \sa_snapshot_ia_wdata.f.lower [18]);
tran (sa_snapshot_ia_wdata[17], \sa_snapshot_ia_wdata.r.part0 [17]);
tran (sa_snapshot_ia_wdata[17], \sa_snapshot_ia_wdata.f.lower [17]);
tran (sa_snapshot_ia_wdata[16], \sa_snapshot_ia_wdata.r.part0 [16]);
tran (sa_snapshot_ia_wdata[16], \sa_snapshot_ia_wdata.f.lower [16]);
tran (sa_snapshot_ia_wdata[15], \sa_snapshot_ia_wdata.r.part0 [15]);
tran (sa_snapshot_ia_wdata[15], \sa_snapshot_ia_wdata.f.lower [15]);
tran (sa_snapshot_ia_wdata[14], \sa_snapshot_ia_wdata.r.part0 [14]);
tran (sa_snapshot_ia_wdata[14], \sa_snapshot_ia_wdata.f.lower [14]);
tran (sa_snapshot_ia_wdata[13], \sa_snapshot_ia_wdata.r.part0 [13]);
tran (sa_snapshot_ia_wdata[13], \sa_snapshot_ia_wdata.f.lower [13]);
tran (sa_snapshot_ia_wdata[12], \sa_snapshot_ia_wdata.r.part0 [12]);
tran (sa_snapshot_ia_wdata[12], \sa_snapshot_ia_wdata.f.lower [12]);
tran (sa_snapshot_ia_wdata[11], \sa_snapshot_ia_wdata.r.part0 [11]);
tran (sa_snapshot_ia_wdata[11], \sa_snapshot_ia_wdata.f.lower [11]);
tran (sa_snapshot_ia_wdata[10], \sa_snapshot_ia_wdata.r.part0 [10]);
tran (sa_snapshot_ia_wdata[10], \sa_snapshot_ia_wdata.f.lower [10]);
tran (sa_snapshot_ia_wdata[9], \sa_snapshot_ia_wdata.r.part0 [9]);
tran (sa_snapshot_ia_wdata[9], \sa_snapshot_ia_wdata.f.lower [9]);
tran (sa_snapshot_ia_wdata[8], \sa_snapshot_ia_wdata.r.part0 [8]);
tran (sa_snapshot_ia_wdata[8], \sa_snapshot_ia_wdata.f.lower [8]);
tran (sa_snapshot_ia_wdata[7], \sa_snapshot_ia_wdata.r.part0 [7]);
tran (sa_snapshot_ia_wdata[7], \sa_snapshot_ia_wdata.f.lower [7]);
tran (sa_snapshot_ia_wdata[6], \sa_snapshot_ia_wdata.r.part0 [6]);
tran (sa_snapshot_ia_wdata[6], \sa_snapshot_ia_wdata.f.lower [6]);
tran (sa_snapshot_ia_wdata[5], \sa_snapshot_ia_wdata.r.part0 [5]);
tran (sa_snapshot_ia_wdata[5], \sa_snapshot_ia_wdata.f.lower [5]);
tran (sa_snapshot_ia_wdata[4], \sa_snapshot_ia_wdata.r.part0 [4]);
tran (sa_snapshot_ia_wdata[4], \sa_snapshot_ia_wdata.f.lower [4]);
tran (sa_snapshot_ia_wdata[3], \sa_snapshot_ia_wdata.r.part0 [3]);
tran (sa_snapshot_ia_wdata[3], \sa_snapshot_ia_wdata.f.lower [3]);
tran (sa_snapshot_ia_wdata[2], \sa_snapshot_ia_wdata.r.part0 [2]);
tran (sa_snapshot_ia_wdata[2], \sa_snapshot_ia_wdata.f.lower [2]);
tran (sa_snapshot_ia_wdata[1], \sa_snapshot_ia_wdata.r.part0 [1]);
tran (sa_snapshot_ia_wdata[1], \sa_snapshot_ia_wdata.f.lower [1]);
tran (sa_snapshot_ia_wdata[0], \sa_snapshot_ia_wdata.r.part0 [0]);
tran (sa_snapshot_ia_wdata[0], \sa_snapshot_ia_wdata.f.lower [0]);
tran (sa_snapshot_ia_wdata[63], \sa_snapshot_ia_wdata.r.part1 [31]);
tran (sa_snapshot_ia_wdata[63], \sa_snapshot_ia_wdata.f.unused [13]);
tran (sa_snapshot_ia_wdata[62], \sa_snapshot_ia_wdata.r.part1 [30]);
tran (sa_snapshot_ia_wdata[62], \sa_snapshot_ia_wdata.f.unused [12]);
tran (sa_snapshot_ia_wdata[61], \sa_snapshot_ia_wdata.r.part1 [29]);
tran (sa_snapshot_ia_wdata[61], \sa_snapshot_ia_wdata.f.unused [11]);
tran (sa_snapshot_ia_wdata[60], \sa_snapshot_ia_wdata.r.part1 [28]);
tran (sa_snapshot_ia_wdata[60], \sa_snapshot_ia_wdata.f.unused [10]);
tran (sa_snapshot_ia_wdata[59], \sa_snapshot_ia_wdata.r.part1 [27]);
tran (sa_snapshot_ia_wdata[59], \sa_snapshot_ia_wdata.f.unused [9]);
tran (sa_snapshot_ia_wdata[58], \sa_snapshot_ia_wdata.r.part1 [26]);
tran (sa_snapshot_ia_wdata[58], \sa_snapshot_ia_wdata.f.unused [8]);
tran (sa_snapshot_ia_wdata[57], \sa_snapshot_ia_wdata.r.part1 [25]);
tran (sa_snapshot_ia_wdata[57], \sa_snapshot_ia_wdata.f.unused [7]);
tran (sa_snapshot_ia_wdata[56], \sa_snapshot_ia_wdata.r.part1 [24]);
tran (sa_snapshot_ia_wdata[56], \sa_snapshot_ia_wdata.f.unused [6]);
tran (sa_snapshot_ia_wdata[55], \sa_snapshot_ia_wdata.r.part1 [23]);
tran (sa_snapshot_ia_wdata[55], \sa_snapshot_ia_wdata.f.unused [5]);
tran (sa_snapshot_ia_wdata[54], \sa_snapshot_ia_wdata.r.part1 [22]);
tran (sa_snapshot_ia_wdata[54], \sa_snapshot_ia_wdata.f.unused [4]);
tran (sa_snapshot_ia_wdata[53], \sa_snapshot_ia_wdata.r.part1 [21]);
tran (sa_snapshot_ia_wdata[53], \sa_snapshot_ia_wdata.f.unused [3]);
tran (sa_snapshot_ia_wdata[52], \sa_snapshot_ia_wdata.r.part1 [20]);
tran (sa_snapshot_ia_wdata[52], \sa_snapshot_ia_wdata.f.unused [2]);
tran (sa_snapshot_ia_wdata[51], \sa_snapshot_ia_wdata.r.part1 [19]);
tran (sa_snapshot_ia_wdata[51], \sa_snapshot_ia_wdata.f.unused [1]);
tran (sa_snapshot_ia_wdata[50], \sa_snapshot_ia_wdata.r.part1 [18]);
tran (sa_snapshot_ia_wdata[50], \sa_snapshot_ia_wdata.f.unused [0]);
tran (sa_snapshot_ia_wdata[49], \sa_snapshot_ia_wdata.r.part1 [17]);
tran (sa_snapshot_ia_wdata[49], \sa_snapshot_ia_wdata.f.upper [17]);
tran (sa_snapshot_ia_wdata[48], \sa_snapshot_ia_wdata.r.part1 [16]);
tran (sa_snapshot_ia_wdata[48], \sa_snapshot_ia_wdata.f.upper [16]);
tran (sa_snapshot_ia_wdata[47], \sa_snapshot_ia_wdata.r.part1 [15]);
tran (sa_snapshot_ia_wdata[47], \sa_snapshot_ia_wdata.f.upper [15]);
tran (sa_snapshot_ia_wdata[46], \sa_snapshot_ia_wdata.r.part1 [14]);
tran (sa_snapshot_ia_wdata[46], \sa_snapshot_ia_wdata.f.upper [14]);
tran (sa_snapshot_ia_wdata[45], \sa_snapshot_ia_wdata.r.part1 [13]);
tran (sa_snapshot_ia_wdata[45], \sa_snapshot_ia_wdata.f.upper [13]);
tran (sa_snapshot_ia_wdata[44], \sa_snapshot_ia_wdata.r.part1 [12]);
tran (sa_snapshot_ia_wdata[44], \sa_snapshot_ia_wdata.f.upper [12]);
tran (sa_snapshot_ia_wdata[43], \sa_snapshot_ia_wdata.r.part1 [11]);
tran (sa_snapshot_ia_wdata[43], \sa_snapshot_ia_wdata.f.upper [11]);
tran (sa_snapshot_ia_wdata[42], \sa_snapshot_ia_wdata.r.part1 [10]);
tran (sa_snapshot_ia_wdata[42], \sa_snapshot_ia_wdata.f.upper [10]);
tran (sa_snapshot_ia_wdata[41], \sa_snapshot_ia_wdata.r.part1 [9]);
tran (sa_snapshot_ia_wdata[41], \sa_snapshot_ia_wdata.f.upper [9]);
tran (sa_snapshot_ia_wdata[40], \sa_snapshot_ia_wdata.r.part1 [8]);
tran (sa_snapshot_ia_wdata[40], \sa_snapshot_ia_wdata.f.upper [8]);
tran (sa_snapshot_ia_wdata[39], \sa_snapshot_ia_wdata.r.part1 [7]);
tran (sa_snapshot_ia_wdata[39], \sa_snapshot_ia_wdata.f.upper [7]);
tran (sa_snapshot_ia_wdata[38], \sa_snapshot_ia_wdata.r.part1 [6]);
tran (sa_snapshot_ia_wdata[38], \sa_snapshot_ia_wdata.f.upper [6]);
tran (sa_snapshot_ia_wdata[37], \sa_snapshot_ia_wdata.r.part1 [5]);
tran (sa_snapshot_ia_wdata[37], \sa_snapshot_ia_wdata.f.upper [5]);
tran (sa_snapshot_ia_wdata[36], \sa_snapshot_ia_wdata.r.part1 [4]);
tran (sa_snapshot_ia_wdata[36], \sa_snapshot_ia_wdata.f.upper [4]);
tran (sa_snapshot_ia_wdata[35], \sa_snapshot_ia_wdata.r.part1 [3]);
tran (sa_snapshot_ia_wdata[35], \sa_snapshot_ia_wdata.f.upper [3]);
tran (sa_snapshot_ia_wdata[34], \sa_snapshot_ia_wdata.r.part1 [2]);
tran (sa_snapshot_ia_wdata[34], \sa_snapshot_ia_wdata.f.upper [2]);
tran (sa_snapshot_ia_wdata[33], \sa_snapshot_ia_wdata.r.part1 [1]);
tran (sa_snapshot_ia_wdata[33], \sa_snapshot_ia_wdata.f.upper [1]);
tran (sa_snapshot_ia_wdata[32], \sa_snapshot_ia_wdata.r.part1 [0]);
tran (sa_snapshot_ia_wdata[32], \sa_snapshot_ia_wdata.f.upper [0]);
tran (sa_snapshot_ia_config[8], \sa_snapshot_ia_config.r.part0 [8]);
tran (sa_snapshot_ia_config[8], \sa_snapshot_ia_config.f.op [3]);
tran (sa_snapshot_ia_config[7], \sa_snapshot_ia_config.r.part0 [7]);
tran (sa_snapshot_ia_config[7], \sa_snapshot_ia_config.f.op [2]);
tran (sa_snapshot_ia_config[6], \sa_snapshot_ia_config.r.part0 [6]);
tran (sa_snapshot_ia_config[6], \sa_snapshot_ia_config.f.op [1]);
tran (sa_snapshot_ia_config[5], \sa_snapshot_ia_config.r.part0 [5]);
tran (sa_snapshot_ia_config[5], \sa_snapshot_ia_config.f.op [0]);
tran (sa_snapshot_ia_config[4], \sa_snapshot_ia_config.r.part0 [4]);
tran (sa_snapshot_ia_config[4], \sa_snapshot_ia_config.f.addr [4]);
tran (sa_snapshot_ia_config[3], \sa_snapshot_ia_config.r.part0 [3]);
tran (sa_snapshot_ia_config[3], \sa_snapshot_ia_config.f.addr [3]);
tran (sa_snapshot_ia_config[2], \sa_snapshot_ia_config.r.part0 [2]);
tran (sa_snapshot_ia_config[2], \sa_snapshot_ia_config.f.addr [2]);
tran (sa_snapshot_ia_config[1], \sa_snapshot_ia_config.r.part0 [1]);
tran (sa_snapshot_ia_config[1], \sa_snapshot_ia_config.f.addr [1]);
tran (sa_snapshot_ia_config[0], \sa_snapshot_ia_config.r.part0 [0]);
tran (sa_snapshot_ia_config[0], \sa_snapshot_ia_config.f.addr [0]);
tran (sa_count_ia_wdata[31], \sa_count_ia_wdata.r.part0 [31]);
tran (sa_count_ia_wdata[31], \sa_count_ia_wdata.f.lower [31]);
tran (sa_count_ia_wdata[30], \sa_count_ia_wdata.r.part0 [30]);
tran (sa_count_ia_wdata[30], \sa_count_ia_wdata.f.lower [30]);
tran (sa_count_ia_wdata[29], \sa_count_ia_wdata.r.part0 [29]);
tran (sa_count_ia_wdata[29], \sa_count_ia_wdata.f.lower [29]);
tran (sa_count_ia_wdata[28], \sa_count_ia_wdata.r.part0 [28]);
tran (sa_count_ia_wdata[28], \sa_count_ia_wdata.f.lower [28]);
tran (sa_count_ia_wdata[27], \sa_count_ia_wdata.r.part0 [27]);
tran (sa_count_ia_wdata[27], \sa_count_ia_wdata.f.lower [27]);
tran (sa_count_ia_wdata[26], \sa_count_ia_wdata.r.part0 [26]);
tran (sa_count_ia_wdata[26], \sa_count_ia_wdata.f.lower [26]);
tran (sa_count_ia_wdata[25], \sa_count_ia_wdata.r.part0 [25]);
tran (sa_count_ia_wdata[25], \sa_count_ia_wdata.f.lower [25]);
tran (sa_count_ia_wdata[24], \sa_count_ia_wdata.r.part0 [24]);
tran (sa_count_ia_wdata[24], \sa_count_ia_wdata.f.lower [24]);
tran (sa_count_ia_wdata[23], \sa_count_ia_wdata.r.part0 [23]);
tran (sa_count_ia_wdata[23], \sa_count_ia_wdata.f.lower [23]);
tran (sa_count_ia_wdata[22], \sa_count_ia_wdata.r.part0 [22]);
tran (sa_count_ia_wdata[22], \sa_count_ia_wdata.f.lower [22]);
tran (sa_count_ia_wdata[21], \sa_count_ia_wdata.r.part0 [21]);
tran (sa_count_ia_wdata[21], \sa_count_ia_wdata.f.lower [21]);
tran (sa_count_ia_wdata[20], \sa_count_ia_wdata.r.part0 [20]);
tran (sa_count_ia_wdata[20], \sa_count_ia_wdata.f.lower [20]);
tran (sa_count_ia_wdata[19], \sa_count_ia_wdata.r.part0 [19]);
tran (sa_count_ia_wdata[19], \sa_count_ia_wdata.f.lower [19]);
tran (sa_count_ia_wdata[18], \sa_count_ia_wdata.r.part0 [18]);
tran (sa_count_ia_wdata[18], \sa_count_ia_wdata.f.lower [18]);
tran (sa_count_ia_wdata[17], \sa_count_ia_wdata.r.part0 [17]);
tran (sa_count_ia_wdata[17], \sa_count_ia_wdata.f.lower [17]);
tran (sa_count_ia_wdata[16], \sa_count_ia_wdata.r.part0 [16]);
tran (sa_count_ia_wdata[16], \sa_count_ia_wdata.f.lower [16]);
tran (sa_count_ia_wdata[15], \sa_count_ia_wdata.r.part0 [15]);
tran (sa_count_ia_wdata[15], \sa_count_ia_wdata.f.lower [15]);
tran (sa_count_ia_wdata[14], \sa_count_ia_wdata.r.part0 [14]);
tran (sa_count_ia_wdata[14], \sa_count_ia_wdata.f.lower [14]);
tran (sa_count_ia_wdata[13], \sa_count_ia_wdata.r.part0 [13]);
tran (sa_count_ia_wdata[13], \sa_count_ia_wdata.f.lower [13]);
tran (sa_count_ia_wdata[12], \sa_count_ia_wdata.r.part0 [12]);
tran (sa_count_ia_wdata[12], \sa_count_ia_wdata.f.lower [12]);
tran (sa_count_ia_wdata[11], \sa_count_ia_wdata.r.part0 [11]);
tran (sa_count_ia_wdata[11], \sa_count_ia_wdata.f.lower [11]);
tran (sa_count_ia_wdata[10], \sa_count_ia_wdata.r.part0 [10]);
tran (sa_count_ia_wdata[10], \sa_count_ia_wdata.f.lower [10]);
tran (sa_count_ia_wdata[9], \sa_count_ia_wdata.r.part0 [9]);
tran (sa_count_ia_wdata[9], \sa_count_ia_wdata.f.lower [9]);
tran (sa_count_ia_wdata[8], \sa_count_ia_wdata.r.part0 [8]);
tran (sa_count_ia_wdata[8], \sa_count_ia_wdata.f.lower [8]);
tran (sa_count_ia_wdata[7], \sa_count_ia_wdata.r.part0 [7]);
tran (sa_count_ia_wdata[7], \sa_count_ia_wdata.f.lower [7]);
tran (sa_count_ia_wdata[6], \sa_count_ia_wdata.r.part0 [6]);
tran (sa_count_ia_wdata[6], \sa_count_ia_wdata.f.lower [6]);
tran (sa_count_ia_wdata[5], \sa_count_ia_wdata.r.part0 [5]);
tran (sa_count_ia_wdata[5], \sa_count_ia_wdata.f.lower [5]);
tran (sa_count_ia_wdata[4], \sa_count_ia_wdata.r.part0 [4]);
tran (sa_count_ia_wdata[4], \sa_count_ia_wdata.f.lower [4]);
tran (sa_count_ia_wdata[3], \sa_count_ia_wdata.r.part0 [3]);
tran (sa_count_ia_wdata[3], \sa_count_ia_wdata.f.lower [3]);
tran (sa_count_ia_wdata[2], \sa_count_ia_wdata.r.part0 [2]);
tran (sa_count_ia_wdata[2], \sa_count_ia_wdata.f.lower [2]);
tran (sa_count_ia_wdata[1], \sa_count_ia_wdata.r.part0 [1]);
tran (sa_count_ia_wdata[1], \sa_count_ia_wdata.f.lower [1]);
tran (sa_count_ia_wdata[0], \sa_count_ia_wdata.r.part0 [0]);
tran (sa_count_ia_wdata[0], \sa_count_ia_wdata.f.lower [0]);
tran (sa_count_ia_wdata[63], \sa_count_ia_wdata.r.part1 [31]);
tran (sa_count_ia_wdata[63], \sa_count_ia_wdata.f.unused [13]);
tran (sa_count_ia_wdata[62], \sa_count_ia_wdata.r.part1 [30]);
tran (sa_count_ia_wdata[62], \sa_count_ia_wdata.f.unused [12]);
tran (sa_count_ia_wdata[61], \sa_count_ia_wdata.r.part1 [29]);
tran (sa_count_ia_wdata[61], \sa_count_ia_wdata.f.unused [11]);
tran (sa_count_ia_wdata[60], \sa_count_ia_wdata.r.part1 [28]);
tran (sa_count_ia_wdata[60], \sa_count_ia_wdata.f.unused [10]);
tran (sa_count_ia_wdata[59], \sa_count_ia_wdata.r.part1 [27]);
tran (sa_count_ia_wdata[59], \sa_count_ia_wdata.f.unused [9]);
tran (sa_count_ia_wdata[58], \sa_count_ia_wdata.r.part1 [26]);
tran (sa_count_ia_wdata[58], \sa_count_ia_wdata.f.unused [8]);
tran (sa_count_ia_wdata[57], \sa_count_ia_wdata.r.part1 [25]);
tran (sa_count_ia_wdata[57], \sa_count_ia_wdata.f.unused [7]);
tran (sa_count_ia_wdata[56], \sa_count_ia_wdata.r.part1 [24]);
tran (sa_count_ia_wdata[56], \sa_count_ia_wdata.f.unused [6]);
tran (sa_count_ia_wdata[55], \sa_count_ia_wdata.r.part1 [23]);
tran (sa_count_ia_wdata[55], \sa_count_ia_wdata.f.unused [5]);
tran (sa_count_ia_wdata[54], \sa_count_ia_wdata.r.part1 [22]);
tran (sa_count_ia_wdata[54], \sa_count_ia_wdata.f.unused [4]);
tran (sa_count_ia_wdata[53], \sa_count_ia_wdata.r.part1 [21]);
tran (sa_count_ia_wdata[53], \sa_count_ia_wdata.f.unused [3]);
tran (sa_count_ia_wdata[52], \sa_count_ia_wdata.r.part1 [20]);
tran (sa_count_ia_wdata[52], \sa_count_ia_wdata.f.unused [2]);
tran (sa_count_ia_wdata[51], \sa_count_ia_wdata.r.part1 [19]);
tran (sa_count_ia_wdata[51], \sa_count_ia_wdata.f.unused [1]);
tran (sa_count_ia_wdata[50], \sa_count_ia_wdata.r.part1 [18]);
tran (sa_count_ia_wdata[50], \sa_count_ia_wdata.f.unused [0]);
tran (sa_count_ia_wdata[49], \sa_count_ia_wdata.r.part1 [17]);
tran (sa_count_ia_wdata[49], \sa_count_ia_wdata.f.upper [17]);
tran (sa_count_ia_wdata[48], \sa_count_ia_wdata.r.part1 [16]);
tran (sa_count_ia_wdata[48], \sa_count_ia_wdata.f.upper [16]);
tran (sa_count_ia_wdata[47], \sa_count_ia_wdata.r.part1 [15]);
tran (sa_count_ia_wdata[47], \sa_count_ia_wdata.f.upper [15]);
tran (sa_count_ia_wdata[46], \sa_count_ia_wdata.r.part1 [14]);
tran (sa_count_ia_wdata[46], \sa_count_ia_wdata.f.upper [14]);
tran (sa_count_ia_wdata[45], \sa_count_ia_wdata.r.part1 [13]);
tran (sa_count_ia_wdata[45], \sa_count_ia_wdata.f.upper [13]);
tran (sa_count_ia_wdata[44], \sa_count_ia_wdata.r.part1 [12]);
tran (sa_count_ia_wdata[44], \sa_count_ia_wdata.f.upper [12]);
tran (sa_count_ia_wdata[43], \sa_count_ia_wdata.r.part1 [11]);
tran (sa_count_ia_wdata[43], \sa_count_ia_wdata.f.upper [11]);
tran (sa_count_ia_wdata[42], \sa_count_ia_wdata.r.part1 [10]);
tran (sa_count_ia_wdata[42], \sa_count_ia_wdata.f.upper [10]);
tran (sa_count_ia_wdata[41], \sa_count_ia_wdata.r.part1 [9]);
tran (sa_count_ia_wdata[41], \sa_count_ia_wdata.f.upper [9]);
tran (sa_count_ia_wdata[40], \sa_count_ia_wdata.r.part1 [8]);
tran (sa_count_ia_wdata[40], \sa_count_ia_wdata.f.upper [8]);
tran (sa_count_ia_wdata[39], \sa_count_ia_wdata.r.part1 [7]);
tran (sa_count_ia_wdata[39], \sa_count_ia_wdata.f.upper [7]);
tran (sa_count_ia_wdata[38], \sa_count_ia_wdata.r.part1 [6]);
tran (sa_count_ia_wdata[38], \sa_count_ia_wdata.f.upper [6]);
tran (sa_count_ia_wdata[37], \sa_count_ia_wdata.r.part1 [5]);
tran (sa_count_ia_wdata[37], \sa_count_ia_wdata.f.upper [5]);
tran (sa_count_ia_wdata[36], \sa_count_ia_wdata.r.part1 [4]);
tran (sa_count_ia_wdata[36], \sa_count_ia_wdata.f.upper [4]);
tran (sa_count_ia_wdata[35], \sa_count_ia_wdata.r.part1 [3]);
tran (sa_count_ia_wdata[35], \sa_count_ia_wdata.f.upper [3]);
tran (sa_count_ia_wdata[34], \sa_count_ia_wdata.r.part1 [2]);
tran (sa_count_ia_wdata[34], \sa_count_ia_wdata.f.upper [2]);
tran (sa_count_ia_wdata[33], \sa_count_ia_wdata.r.part1 [1]);
tran (sa_count_ia_wdata[33], \sa_count_ia_wdata.f.upper [1]);
tran (sa_count_ia_wdata[32], \sa_count_ia_wdata.r.part1 [0]);
tran (sa_count_ia_wdata[32], \sa_count_ia_wdata.f.upper [0]);
tran (sa_count_ia_config[8], \sa_count_ia_config.r.part0 [8]);
tran (sa_count_ia_config[8], \sa_count_ia_config.f.op [3]);
tran (sa_count_ia_config[7], \sa_count_ia_config.r.part0 [7]);
tran (sa_count_ia_config[7], \sa_count_ia_config.f.op [2]);
tran (sa_count_ia_config[6], \sa_count_ia_config.r.part0 [6]);
tran (sa_count_ia_config[6], \sa_count_ia_config.f.op [1]);
tran (sa_count_ia_config[5], \sa_count_ia_config.r.part0 [5]);
tran (sa_count_ia_config[5], \sa_count_ia_config.f.op [0]);
tran (sa_count_ia_config[4], \sa_count_ia_config.r.part0 [4]);
tran (sa_count_ia_config[4], \sa_count_ia_config.f.addr [4]);
tran (sa_count_ia_config[3], \sa_count_ia_config.r.part0 [3]);
tran (sa_count_ia_config[3], \sa_count_ia_config.f.addr [3]);
tran (sa_count_ia_config[2], \sa_count_ia_config.r.part0 [2]);
tran (sa_count_ia_config[2], \sa_count_ia_config.f.addr [2]);
tran (sa_count_ia_config[1], \sa_count_ia_config.r.part0 [1]);
tran (sa_count_ia_config[1], \sa_count_ia_config.f.addr [1]);
tran (sa_count_ia_config[0], \sa_count_ia_config.r.part0 [0]);
tran (sa_count_ia_config[0], \sa_count_ia_config.f.addr [0]);
tran (sa_ctrl_ia_wdata[31], \sa_ctrl_ia_wdata.r.part0 [31]);
tran (sa_ctrl_ia_wdata[31], \sa_ctrl_ia_wdata.f.spare [26]);
tran (sa_ctrl_ia_wdata[30], \sa_ctrl_ia_wdata.r.part0 [30]);
tran (sa_ctrl_ia_wdata[30], \sa_ctrl_ia_wdata.f.spare [25]);
tran (sa_ctrl_ia_wdata[29], \sa_ctrl_ia_wdata.r.part0 [29]);
tran (sa_ctrl_ia_wdata[29], \sa_ctrl_ia_wdata.f.spare [24]);
tran (sa_ctrl_ia_wdata[28], \sa_ctrl_ia_wdata.r.part0 [28]);
tran (sa_ctrl_ia_wdata[28], \sa_ctrl_ia_wdata.f.spare [23]);
tran (sa_ctrl_ia_wdata[27], \sa_ctrl_ia_wdata.r.part0 [27]);
tran (sa_ctrl_ia_wdata[27], \sa_ctrl_ia_wdata.f.spare [22]);
tran (sa_ctrl_ia_wdata[26], \sa_ctrl_ia_wdata.r.part0 [26]);
tran (sa_ctrl_ia_wdata[26], \sa_ctrl_ia_wdata.f.spare [21]);
tran (sa_ctrl_ia_wdata[25], \sa_ctrl_ia_wdata.r.part0 [25]);
tran (sa_ctrl_ia_wdata[25], \sa_ctrl_ia_wdata.f.spare [20]);
tran (sa_ctrl_ia_wdata[24], \sa_ctrl_ia_wdata.r.part0 [24]);
tran (sa_ctrl_ia_wdata[24], \sa_ctrl_ia_wdata.f.spare [19]);
tran (sa_ctrl_ia_wdata[23], \sa_ctrl_ia_wdata.r.part0 [23]);
tran (sa_ctrl_ia_wdata[23], \sa_ctrl_ia_wdata.f.spare [18]);
tran (sa_ctrl_ia_wdata[22], \sa_ctrl_ia_wdata.r.part0 [22]);
tran (sa_ctrl_ia_wdata[22], \sa_ctrl_ia_wdata.f.spare [17]);
tran (sa_ctrl_ia_wdata[21], \sa_ctrl_ia_wdata.r.part0 [21]);
tran (sa_ctrl_ia_wdata[21], \sa_ctrl_ia_wdata.f.spare [16]);
tran (sa_ctrl_ia_wdata[20], \sa_ctrl_ia_wdata.r.part0 [20]);
tran (sa_ctrl_ia_wdata[20], \sa_ctrl_ia_wdata.f.spare [15]);
tran (sa_ctrl_ia_wdata[19], \sa_ctrl_ia_wdata.r.part0 [19]);
tran (sa_ctrl_ia_wdata[19], \sa_ctrl_ia_wdata.f.spare [14]);
tran (sa_ctrl_ia_wdata[18], \sa_ctrl_ia_wdata.r.part0 [18]);
tran (sa_ctrl_ia_wdata[18], \sa_ctrl_ia_wdata.f.spare [13]);
tran (sa_ctrl_ia_wdata[17], \sa_ctrl_ia_wdata.r.part0 [17]);
tran (sa_ctrl_ia_wdata[17], \sa_ctrl_ia_wdata.f.spare [12]);
tran (sa_ctrl_ia_wdata[16], \sa_ctrl_ia_wdata.r.part0 [16]);
tran (sa_ctrl_ia_wdata[16], \sa_ctrl_ia_wdata.f.spare [11]);
tran (sa_ctrl_ia_wdata[15], \sa_ctrl_ia_wdata.r.part0 [15]);
tran (sa_ctrl_ia_wdata[15], \sa_ctrl_ia_wdata.f.spare [10]);
tran (sa_ctrl_ia_wdata[14], \sa_ctrl_ia_wdata.r.part0 [14]);
tran (sa_ctrl_ia_wdata[14], \sa_ctrl_ia_wdata.f.spare [9]);
tran (sa_ctrl_ia_wdata[13], \sa_ctrl_ia_wdata.r.part0 [13]);
tran (sa_ctrl_ia_wdata[13], \sa_ctrl_ia_wdata.f.spare [8]);
tran (sa_ctrl_ia_wdata[12], \sa_ctrl_ia_wdata.r.part0 [12]);
tran (sa_ctrl_ia_wdata[12], \sa_ctrl_ia_wdata.f.spare [7]);
tran (sa_ctrl_ia_wdata[11], \sa_ctrl_ia_wdata.r.part0 [11]);
tran (sa_ctrl_ia_wdata[11], \sa_ctrl_ia_wdata.f.spare [6]);
tran (sa_ctrl_ia_wdata[10], \sa_ctrl_ia_wdata.r.part0 [10]);
tran (sa_ctrl_ia_wdata[10], \sa_ctrl_ia_wdata.f.spare [5]);
tran (sa_ctrl_ia_wdata[9], \sa_ctrl_ia_wdata.r.part0 [9]);
tran (sa_ctrl_ia_wdata[9], \sa_ctrl_ia_wdata.f.spare [4]);
tran (sa_ctrl_ia_wdata[8], \sa_ctrl_ia_wdata.r.part0 [8]);
tran (sa_ctrl_ia_wdata[8], \sa_ctrl_ia_wdata.f.spare [3]);
tran (sa_ctrl_ia_wdata[7], \sa_ctrl_ia_wdata.r.part0 [7]);
tran (sa_ctrl_ia_wdata[7], \sa_ctrl_ia_wdata.f.spare [2]);
tran (sa_ctrl_ia_wdata[6], \sa_ctrl_ia_wdata.r.part0 [6]);
tran (sa_ctrl_ia_wdata[6], \sa_ctrl_ia_wdata.f.spare [1]);
tran (sa_ctrl_ia_wdata[5], \sa_ctrl_ia_wdata.r.part0 [5]);
tran (sa_ctrl_ia_wdata[5], \sa_ctrl_ia_wdata.f.spare [0]);
tran (sa_ctrl_ia_wdata[4], \sa_ctrl_ia_wdata.r.part0 [4]);
tran (sa_ctrl_ia_wdata[4], \sa_ctrl_ia_wdata.f.sa_event_sel [4]);
tran (sa_ctrl_ia_wdata[3], \sa_ctrl_ia_wdata.r.part0 [3]);
tran (sa_ctrl_ia_wdata[3], \sa_ctrl_ia_wdata.f.sa_event_sel [3]);
tran (sa_ctrl_ia_wdata[2], \sa_ctrl_ia_wdata.r.part0 [2]);
tran (sa_ctrl_ia_wdata[2], \sa_ctrl_ia_wdata.f.sa_event_sel [2]);
tran (sa_ctrl_ia_wdata[1], \sa_ctrl_ia_wdata.r.part0 [1]);
tran (sa_ctrl_ia_wdata[1], \sa_ctrl_ia_wdata.f.sa_event_sel [1]);
tran (sa_ctrl_ia_wdata[0], \sa_ctrl_ia_wdata.r.part0 [0]);
tran (sa_ctrl_ia_wdata[0], \sa_ctrl_ia_wdata.f.sa_event_sel [0]);
tran (sa_ctrl_ia_config[8], \sa_ctrl_ia_config.r.part0 [8]);
tran (sa_ctrl_ia_config[8], \sa_ctrl_ia_config.f.op [3]);
tran (sa_ctrl_ia_config[7], \sa_ctrl_ia_config.r.part0 [7]);
tran (sa_ctrl_ia_config[7], \sa_ctrl_ia_config.f.op [2]);
tran (sa_ctrl_ia_config[6], \sa_ctrl_ia_config.r.part0 [6]);
tran (sa_ctrl_ia_config[6], \sa_ctrl_ia_config.f.op [1]);
tran (sa_ctrl_ia_config[5], \sa_ctrl_ia_config.r.part0 [5]);
tran (sa_ctrl_ia_config[5], \sa_ctrl_ia_config.f.op [0]);
tran (sa_ctrl_ia_config[4], \sa_ctrl_ia_config.r.part0 [4]);
tran (sa_ctrl_ia_config[4], \sa_ctrl_ia_config.f.addr [4]);
tran (sa_ctrl_ia_config[3], \sa_ctrl_ia_config.r.part0 [3]);
tran (sa_ctrl_ia_config[3], \sa_ctrl_ia_config.f.addr [3]);
tran (sa_ctrl_ia_config[2], \sa_ctrl_ia_config.r.part0 [2]);
tran (sa_ctrl_ia_config[2], \sa_ctrl_ia_config.f.addr [2]);
tran (sa_ctrl_ia_config[1], \sa_ctrl_ia_config.r.part0 [1]);
tran (sa_ctrl_ia_config[1], \sa_ctrl_ia_config.f.addr [1]);
tran (sa_ctrl_ia_config[0], \sa_ctrl_ia_config.r.part0 [0]);
tran (sa_ctrl_ia_config[0], \sa_ctrl_ia_config.f.addr [0]);
tran (kme_cceip0_ob_out_post[82], \kme_cceip0_ob_out_post.tvalid );
tran (kme_cceip0_ob_out_post[81], \kme_cceip0_ob_out_post.tlast );
tran (kme_cceip0_ob_out_post[80], \kme_cceip0_ob_out_post.tid [0]);
tran (kme_cceip0_ob_out_post[79], \kme_cceip0_ob_out_post.tstrb [7]);
tran (kme_cceip0_ob_out_post[78], \kme_cceip0_ob_out_post.tstrb [6]);
tran (kme_cceip0_ob_out_post[77], \kme_cceip0_ob_out_post.tstrb [5]);
tran (kme_cceip0_ob_out_post[76], \kme_cceip0_ob_out_post.tstrb [4]);
tran (kme_cceip0_ob_out_post[75], \kme_cceip0_ob_out_post.tstrb [3]);
tran (kme_cceip0_ob_out_post[74], \kme_cceip0_ob_out_post.tstrb [2]);
tran (kme_cceip0_ob_out_post[73], \kme_cceip0_ob_out_post.tstrb [1]);
tran (kme_cceip0_ob_out_post[72], \kme_cceip0_ob_out_post.tstrb [0]);
tran (kme_cceip0_ob_out_post[71], \kme_cceip0_ob_out_post.tuser [7]);
tran (kme_cceip0_ob_out_post[70], \kme_cceip0_ob_out_post.tuser [6]);
tran (kme_cceip0_ob_out_post[69], \kme_cceip0_ob_out_post.tuser [5]);
tran (kme_cceip0_ob_out_post[68], \kme_cceip0_ob_out_post.tuser [4]);
tran (kme_cceip0_ob_out_post[67], \kme_cceip0_ob_out_post.tuser [3]);
tran (kme_cceip0_ob_out_post[66], \kme_cceip0_ob_out_post.tuser [2]);
tran (kme_cceip0_ob_out_post[65], \kme_cceip0_ob_out_post.tuser [1]);
tran (kme_cceip0_ob_out_post[64], \kme_cceip0_ob_out_post.tuser [0]);
tran (kme_cceip0_ob_out_post[63], \kme_cceip0_ob_out_post.tdata [63]);
tran (kme_cceip0_ob_out_post[62], \kme_cceip0_ob_out_post.tdata [62]);
tran (kme_cceip0_ob_out_post[61], \kme_cceip0_ob_out_post.tdata [61]);
tran (kme_cceip0_ob_out_post[60], \kme_cceip0_ob_out_post.tdata [60]);
tran (kme_cceip0_ob_out_post[59], \kme_cceip0_ob_out_post.tdata [59]);
tran (kme_cceip0_ob_out_post[58], \kme_cceip0_ob_out_post.tdata [58]);
tran (kme_cceip0_ob_out_post[57], \kme_cceip0_ob_out_post.tdata [57]);
tran (kme_cceip0_ob_out_post[56], \kme_cceip0_ob_out_post.tdata [56]);
tran (kme_cceip0_ob_out_post[55], \kme_cceip0_ob_out_post.tdata [55]);
tran (kme_cceip0_ob_out_post[54], \kme_cceip0_ob_out_post.tdata [54]);
tran (kme_cceip0_ob_out_post[53], \kme_cceip0_ob_out_post.tdata [53]);
tran (kme_cceip0_ob_out_post[52], \kme_cceip0_ob_out_post.tdata [52]);
tran (kme_cceip0_ob_out_post[51], \kme_cceip0_ob_out_post.tdata [51]);
tran (kme_cceip0_ob_out_post[50], \kme_cceip0_ob_out_post.tdata [50]);
tran (kme_cceip0_ob_out_post[49], \kme_cceip0_ob_out_post.tdata [49]);
tran (kme_cceip0_ob_out_post[48], \kme_cceip0_ob_out_post.tdata [48]);
tran (kme_cceip0_ob_out_post[47], \kme_cceip0_ob_out_post.tdata [47]);
tran (kme_cceip0_ob_out_post[46], \kme_cceip0_ob_out_post.tdata [46]);
tran (kme_cceip0_ob_out_post[45], \kme_cceip0_ob_out_post.tdata [45]);
tran (kme_cceip0_ob_out_post[44], \kme_cceip0_ob_out_post.tdata [44]);
tran (kme_cceip0_ob_out_post[43], \kme_cceip0_ob_out_post.tdata [43]);
tran (kme_cceip0_ob_out_post[42], \kme_cceip0_ob_out_post.tdata [42]);
tran (kme_cceip0_ob_out_post[41], \kme_cceip0_ob_out_post.tdata [41]);
tran (kme_cceip0_ob_out_post[40], \kme_cceip0_ob_out_post.tdata [40]);
tran (kme_cceip0_ob_out_post[39], \kme_cceip0_ob_out_post.tdata [39]);
tran (kme_cceip0_ob_out_post[38], \kme_cceip0_ob_out_post.tdata [38]);
tran (kme_cceip0_ob_out_post[37], \kme_cceip0_ob_out_post.tdata [37]);
tran (kme_cceip0_ob_out_post[36], \kme_cceip0_ob_out_post.tdata [36]);
tran (kme_cceip0_ob_out_post[35], \kme_cceip0_ob_out_post.tdata [35]);
tran (kme_cceip0_ob_out_post[34], \kme_cceip0_ob_out_post.tdata [34]);
tran (kme_cceip0_ob_out_post[33], \kme_cceip0_ob_out_post.tdata [33]);
tran (kme_cceip0_ob_out_post[32], \kme_cceip0_ob_out_post.tdata [32]);
tran (kme_cceip0_ob_out_post[31], \kme_cceip0_ob_out_post.tdata [31]);
tran (kme_cceip0_ob_out_post[30], \kme_cceip0_ob_out_post.tdata [30]);
tran (kme_cceip0_ob_out_post[29], \kme_cceip0_ob_out_post.tdata [29]);
tran (kme_cceip0_ob_out_post[28], \kme_cceip0_ob_out_post.tdata [28]);
tran (kme_cceip0_ob_out_post[27], \kme_cceip0_ob_out_post.tdata [27]);
tran (kme_cceip0_ob_out_post[26], \kme_cceip0_ob_out_post.tdata [26]);
tran (kme_cceip0_ob_out_post[25], \kme_cceip0_ob_out_post.tdata [25]);
tran (kme_cceip0_ob_out_post[24], \kme_cceip0_ob_out_post.tdata [24]);
tran (kme_cceip0_ob_out_post[23], \kme_cceip0_ob_out_post.tdata [23]);
tran (kme_cceip0_ob_out_post[22], \kme_cceip0_ob_out_post.tdata [22]);
tran (kme_cceip0_ob_out_post[21], \kme_cceip0_ob_out_post.tdata [21]);
tran (kme_cceip0_ob_out_post[20], \kme_cceip0_ob_out_post.tdata [20]);
tran (kme_cceip0_ob_out_post[19], \kme_cceip0_ob_out_post.tdata [19]);
tran (kme_cceip0_ob_out_post[18], \kme_cceip0_ob_out_post.tdata [18]);
tran (kme_cceip0_ob_out_post[17], \kme_cceip0_ob_out_post.tdata [17]);
tran (kme_cceip0_ob_out_post[16], \kme_cceip0_ob_out_post.tdata [16]);
tran (kme_cceip0_ob_out_post[15], \kme_cceip0_ob_out_post.tdata [15]);
tran (kme_cceip0_ob_out_post[14], \kme_cceip0_ob_out_post.tdata [14]);
tran (kme_cceip0_ob_out_post[13], \kme_cceip0_ob_out_post.tdata [13]);
tran (kme_cceip0_ob_out_post[12], \kme_cceip0_ob_out_post.tdata [12]);
tran (kme_cceip0_ob_out_post[11], \kme_cceip0_ob_out_post.tdata [11]);
tran (kme_cceip0_ob_out_post[10], \kme_cceip0_ob_out_post.tdata [10]);
tran (kme_cceip0_ob_out_post[9], \kme_cceip0_ob_out_post.tdata [9]);
tran (kme_cceip0_ob_out_post[8], \kme_cceip0_ob_out_post.tdata [8]);
tran (kme_cceip0_ob_out_post[7], \kme_cceip0_ob_out_post.tdata [7]);
tran (kme_cceip0_ob_out_post[6], \kme_cceip0_ob_out_post.tdata [6]);
tran (kme_cceip0_ob_out_post[5], \kme_cceip0_ob_out_post.tdata [5]);
tran (kme_cceip0_ob_out_post[4], \kme_cceip0_ob_out_post.tdata [4]);
tran (kme_cceip0_ob_out_post[3], \kme_cceip0_ob_out_post.tdata [3]);
tran (kme_cceip0_ob_out_post[2], \kme_cceip0_ob_out_post.tdata [2]);
tran (kme_cceip0_ob_out_post[1], \kme_cceip0_ob_out_post.tdata [1]);
tran (kme_cceip0_ob_out_post[0], \kme_cceip0_ob_out_post.tdata [0]);
tran (kme_cceip1_ob_out_post[82], \kme_cceip1_ob_out_post.tvalid );
tran (kme_cceip1_ob_out_post[81], \kme_cceip1_ob_out_post.tlast );
tran (kme_cceip1_ob_out_post[80], \kme_cceip1_ob_out_post.tid [0]);
tran (kme_cceip1_ob_out_post[79], \kme_cceip1_ob_out_post.tstrb [7]);
tran (kme_cceip1_ob_out_post[78], \kme_cceip1_ob_out_post.tstrb [6]);
tran (kme_cceip1_ob_out_post[77], \kme_cceip1_ob_out_post.tstrb [5]);
tran (kme_cceip1_ob_out_post[76], \kme_cceip1_ob_out_post.tstrb [4]);
tran (kme_cceip1_ob_out_post[75], \kme_cceip1_ob_out_post.tstrb [3]);
tran (kme_cceip1_ob_out_post[74], \kme_cceip1_ob_out_post.tstrb [2]);
tran (kme_cceip1_ob_out_post[73], \kme_cceip1_ob_out_post.tstrb [1]);
tran (kme_cceip1_ob_out_post[72], \kme_cceip1_ob_out_post.tstrb [0]);
tran (kme_cceip1_ob_out_post[71], \kme_cceip1_ob_out_post.tuser [7]);
tran (kme_cceip1_ob_out_post[70], \kme_cceip1_ob_out_post.tuser [6]);
tran (kme_cceip1_ob_out_post[69], \kme_cceip1_ob_out_post.tuser [5]);
tran (kme_cceip1_ob_out_post[68], \kme_cceip1_ob_out_post.tuser [4]);
tran (kme_cceip1_ob_out_post[67], \kme_cceip1_ob_out_post.tuser [3]);
tran (kme_cceip1_ob_out_post[66], \kme_cceip1_ob_out_post.tuser [2]);
tran (kme_cceip1_ob_out_post[65], \kme_cceip1_ob_out_post.tuser [1]);
tran (kme_cceip1_ob_out_post[64], \kme_cceip1_ob_out_post.tuser [0]);
tran (kme_cceip1_ob_out_post[63], \kme_cceip1_ob_out_post.tdata [63]);
tran (kme_cceip1_ob_out_post[62], \kme_cceip1_ob_out_post.tdata [62]);
tran (kme_cceip1_ob_out_post[61], \kme_cceip1_ob_out_post.tdata [61]);
tran (kme_cceip1_ob_out_post[60], \kme_cceip1_ob_out_post.tdata [60]);
tran (kme_cceip1_ob_out_post[59], \kme_cceip1_ob_out_post.tdata [59]);
tran (kme_cceip1_ob_out_post[58], \kme_cceip1_ob_out_post.tdata [58]);
tran (kme_cceip1_ob_out_post[57], \kme_cceip1_ob_out_post.tdata [57]);
tran (kme_cceip1_ob_out_post[56], \kme_cceip1_ob_out_post.tdata [56]);
tran (kme_cceip1_ob_out_post[55], \kme_cceip1_ob_out_post.tdata [55]);
tran (kme_cceip1_ob_out_post[54], \kme_cceip1_ob_out_post.tdata [54]);
tran (kme_cceip1_ob_out_post[53], \kme_cceip1_ob_out_post.tdata [53]);
tran (kme_cceip1_ob_out_post[52], \kme_cceip1_ob_out_post.tdata [52]);
tran (kme_cceip1_ob_out_post[51], \kme_cceip1_ob_out_post.tdata [51]);
tran (kme_cceip1_ob_out_post[50], \kme_cceip1_ob_out_post.tdata [50]);
tran (kme_cceip1_ob_out_post[49], \kme_cceip1_ob_out_post.tdata [49]);
tran (kme_cceip1_ob_out_post[48], \kme_cceip1_ob_out_post.tdata [48]);
tran (kme_cceip1_ob_out_post[47], \kme_cceip1_ob_out_post.tdata [47]);
tran (kme_cceip1_ob_out_post[46], \kme_cceip1_ob_out_post.tdata [46]);
tran (kme_cceip1_ob_out_post[45], \kme_cceip1_ob_out_post.tdata [45]);
tran (kme_cceip1_ob_out_post[44], \kme_cceip1_ob_out_post.tdata [44]);
tran (kme_cceip1_ob_out_post[43], \kme_cceip1_ob_out_post.tdata [43]);
tran (kme_cceip1_ob_out_post[42], \kme_cceip1_ob_out_post.tdata [42]);
tran (kme_cceip1_ob_out_post[41], \kme_cceip1_ob_out_post.tdata [41]);
tran (kme_cceip1_ob_out_post[40], \kme_cceip1_ob_out_post.tdata [40]);
tran (kme_cceip1_ob_out_post[39], \kme_cceip1_ob_out_post.tdata [39]);
tran (kme_cceip1_ob_out_post[38], \kme_cceip1_ob_out_post.tdata [38]);
tran (kme_cceip1_ob_out_post[37], \kme_cceip1_ob_out_post.tdata [37]);
tran (kme_cceip1_ob_out_post[36], \kme_cceip1_ob_out_post.tdata [36]);
tran (kme_cceip1_ob_out_post[35], \kme_cceip1_ob_out_post.tdata [35]);
tran (kme_cceip1_ob_out_post[34], \kme_cceip1_ob_out_post.tdata [34]);
tran (kme_cceip1_ob_out_post[33], \kme_cceip1_ob_out_post.tdata [33]);
tran (kme_cceip1_ob_out_post[32], \kme_cceip1_ob_out_post.tdata [32]);
tran (kme_cceip1_ob_out_post[31], \kme_cceip1_ob_out_post.tdata [31]);
tran (kme_cceip1_ob_out_post[30], \kme_cceip1_ob_out_post.tdata [30]);
tran (kme_cceip1_ob_out_post[29], \kme_cceip1_ob_out_post.tdata [29]);
tran (kme_cceip1_ob_out_post[28], \kme_cceip1_ob_out_post.tdata [28]);
tran (kme_cceip1_ob_out_post[27], \kme_cceip1_ob_out_post.tdata [27]);
tran (kme_cceip1_ob_out_post[26], \kme_cceip1_ob_out_post.tdata [26]);
tran (kme_cceip1_ob_out_post[25], \kme_cceip1_ob_out_post.tdata [25]);
tran (kme_cceip1_ob_out_post[24], \kme_cceip1_ob_out_post.tdata [24]);
tran (kme_cceip1_ob_out_post[23], \kme_cceip1_ob_out_post.tdata [23]);
tran (kme_cceip1_ob_out_post[22], \kme_cceip1_ob_out_post.tdata [22]);
tran (kme_cceip1_ob_out_post[21], \kme_cceip1_ob_out_post.tdata [21]);
tran (kme_cceip1_ob_out_post[20], \kme_cceip1_ob_out_post.tdata [20]);
tran (kme_cceip1_ob_out_post[19], \kme_cceip1_ob_out_post.tdata [19]);
tran (kme_cceip1_ob_out_post[18], \kme_cceip1_ob_out_post.tdata [18]);
tran (kme_cceip1_ob_out_post[17], \kme_cceip1_ob_out_post.tdata [17]);
tran (kme_cceip1_ob_out_post[16], \kme_cceip1_ob_out_post.tdata [16]);
tran (kme_cceip1_ob_out_post[15], \kme_cceip1_ob_out_post.tdata [15]);
tran (kme_cceip1_ob_out_post[14], \kme_cceip1_ob_out_post.tdata [14]);
tran (kme_cceip1_ob_out_post[13], \kme_cceip1_ob_out_post.tdata [13]);
tran (kme_cceip1_ob_out_post[12], \kme_cceip1_ob_out_post.tdata [12]);
tran (kme_cceip1_ob_out_post[11], \kme_cceip1_ob_out_post.tdata [11]);
tran (kme_cceip1_ob_out_post[10], \kme_cceip1_ob_out_post.tdata [10]);
tran (kme_cceip1_ob_out_post[9], \kme_cceip1_ob_out_post.tdata [9]);
tran (kme_cceip1_ob_out_post[8], \kme_cceip1_ob_out_post.tdata [8]);
tran (kme_cceip1_ob_out_post[7], \kme_cceip1_ob_out_post.tdata [7]);
tran (kme_cceip1_ob_out_post[6], \kme_cceip1_ob_out_post.tdata [6]);
tran (kme_cceip1_ob_out_post[5], \kme_cceip1_ob_out_post.tdata [5]);
tran (kme_cceip1_ob_out_post[4], \kme_cceip1_ob_out_post.tdata [4]);
tran (kme_cceip1_ob_out_post[3], \kme_cceip1_ob_out_post.tdata [3]);
tran (kme_cceip1_ob_out_post[2], \kme_cceip1_ob_out_post.tdata [2]);
tran (kme_cceip1_ob_out_post[1], \kme_cceip1_ob_out_post.tdata [1]);
tran (kme_cceip1_ob_out_post[0], \kme_cceip1_ob_out_post.tdata [0]);
tran (kme_cceip2_ob_out_post[82], \kme_cceip2_ob_out_post.tvalid );
tran (kme_cceip2_ob_out_post[81], \kme_cceip2_ob_out_post.tlast );
tran (kme_cceip2_ob_out_post[80], \kme_cceip2_ob_out_post.tid [0]);
tran (kme_cceip2_ob_out_post[79], \kme_cceip2_ob_out_post.tstrb [7]);
tran (kme_cceip2_ob_out_post[78], \kme_cceip2_ob_out_post.tstrb [6]);
tran (kme_cceip2_ob_out_post[77], \kme_cceip2_ob_out_post.tstrb [5]);
tran (kme_cceip2_ob_out_post[76], \kme_cceip2_ob_out_post.tstrb [4]);
tran (kme_cceip2_ob_out_post[75], \kme_cceip2_ob_out_post.tstrb [3]);
tran (kme_cceip2_ob_out_post[74], \kme_cceip2_ob_out_post.tstrb [2]);
tran (kme_cceip2_ob_out_post[73], \kme_cceip2_ob_out_post.tstrb [1]);
tran (kme_cceip2_ob_out_post[72], \kme_cceip2_ob_out_post.tstrb [0]);
tran (kme_cceip2_ob_out_post[71], \kme_cceip2_ob_out_post.tuser [7]);
tran (kme_cceip2_ob_out_post[70], \kme_cceip2_ob_out_post.tuser [6]);
tran (kme_cceip2_ob_out_post[69], \kme_cceip2_ob_out_post.tuser [5]);
tran (kme_cceip2_ob_out_post[68], \kme_cceip2_ob_out_post.tuser [4]);
tran (kme_cceip2_ob_out_post[67], \kme_cceip2_ob_out_post.tuser [3]);
tran (kme_cceip2_ob_out_post[66], \kme_cceip2_ob_out_post.tuser [2]);
tran (kme_cceip2_ob_out_post[65], \kme_cceip2_ob_out_post.tuser [1]);
tran (kme_cceip2_ob_out_post[64], \kme_cceip2_ob_out_post.tuser [0]);
tran (kme_cceip2_ob_out_post[63], \kme_cceip2_ob_out_post.tdata [63]);
tran (kme_cceip2_ob_out_post[62], \kme_cceip2_ob_out_post.tdata [62]);
tran (kme_cceip2_ob_out_post[61], \kme_cceip2_ob_out_post.tdata [61]);
tran (kme_cceip2_ob_out_post[60], \kme_cceip2_ob_out_post.tdata [60]);
tran (kme_cceip2_ob_out_post[59], \kme_cceip2_ob_out_post.tdata [59]);
tran (kme_cceip2_ob_out_post[58], \kme_cceip2_ob_out_post.tdata [58]);
tran (kme_cceip2_ob_out_post[57], \kme_cceip2_ob_out_post.tdata [57]);
tran (kme_cceip2_ob_out_post[56], \kme_cceip2_ob_out_post.tdata [56]);
tran (kme_cceip2_ob_out_post[55], \kme_cceip2_ob_out_post.tdata [55]);
tran (kme_cceip2_ob_out_post[54], \kme_cceip2_ob_out_post.tdata [54]);
tran (kme_cceip2_ob_out_post[53], \kme_cceip2_ob_out_post.tdata [53]);
tran (kme_cceip2_ob_out_post[52], \kme_cceip2_ob_out_post.tdata [52]);
tran (kme_cceip2_ob_out_post[51], \kme_cceip2_ob_out_post.tdata [51]);
tran (kme_cceip2_ob_out_post[50], \kme_cceip2_ob_out_post.tdata [50]);
tran (kme_cceip2_ob_out_post[49], \kme_cceip2_ob_out_post.tdata [49]);
tran (kme_cceip2_ob_out_post[48], \kme_cceip2_ob_out_post.tdata [48]);
tran (kme_cceip2_ob_out_post[47], \kme_cceip2_ob_out_post.tdata [47]);
tran (kme_cceip2_ob_out_post[46], \kme_cceip2_ob_out_post.tdata [46]);
tran (kme_cceip2_ob_out_post[45], \kme_cceip2_ob_out_post.tdata [45]);
tran (kme_cceip2_ob_out_post[44], \kme_cceip2_ob_out_post.tdata [44]);
tran (kme_cceip2_ob_out_post[43], \kme_cceip2_ob_out_post.tdata [43]);
tran (kme_cceip2_ob_out_post[42], \kme_cceip2_ob_out_post.tdata [42]);
tran (kme_cceip2_ob_out_post[41], \kme_cceip2_ob_out_post.tdata [41]);
tran (kme_cceip2_ob_out_post[40], \kme_cceip2_ob_out_post.tdata [40]);
tran (kme_cceip2_ob_out_post[39], \kme_cceip2_ob_out_post.tdata [39]);
tran (kme_cceip2_ob_out_post[38], \kme_cceip2_ob_out_post.tdata [38]);
tran (kme_cceip2_ob_out_post[37], \kme_cceip2_ob_out_post.tdata [37]);
tran (kme_cceip2_ob_out_post[36], \kme_cceip2_ob_out_post.tdata [36]);
tran (kme_cceip2_ob_out_post[35], \kme_cceip2_ob_out_post.tdata [35]);
tran (kme_cceip2_ob_out_post[34], \kme_cceip2_ob_out_post.tdata [34]);
tran (kme_cceip2_ob_out_post[33], \kme_cceip2_ob_out_post.tdata [33]);
tran (kme_cceip2_ob_out_post[32], \kme_cceip2_ob_out_post.tdata [32]);
tran (kme_cceip2_ob_out_post[31], \kme_cceip2_ob_out_post.tdata [31]);
tran (kme_cceip2_ob_out_post[30], \kme_cceip2_ob_out_post.tdata [30]);
tran (kme_cceip2_ob_out_post[29], \kme_cceip2_ob_out_post.tdata [29]);
tran (kme_cceip2_ob_out_post[28], \kme_cceip2_ob_out_post.tdata [28]);
tran (kme_cceip2_ob_out_post[27], \kme_cceip2_ob_out_post.tdata [27]);
tran (kme_cceip2_ob_out_post[26], \kme_cceip2_ob_out_post.tdata [26]);
tran (kme_cceip2_ob_out_post[25], \kme_cceip2_ob_out_post.tdata [25]);
tran (kme_cceip2_ob_out_post[24], \kme_cceip2_ob_out_post.tdata [24]);
tran (kme_cceip2_ob_out_post[23], \kme_cceip2_ob_out_post.tdata [23]);
tran (kme_cceip2_ob_out_post[22], \kme_cceip2_ob_out_post.tdata [22]);
tran (kme_cceip2_ob_out_post[21], \kme_cceip2_ob_out_post.tdata [21]);
tran (kme_cceip2_ob_out_post[20], \kme_cceip2_ob_out_post.tdata [20]);
tran (kme_cceip2_ob_out_post[19], \kme_cceip2_ob_out_post.tdata [19]);
tran (kme_cceip2_ob_out_post[18], \kme_cceip2_ob_out_post.tdata [18]);
tran (kme_cceip2_ob_out_post[17], \kme_cceip2_ob_out_post.tdata [17]);
tran (kme_cceip2_ob_out_post[16], \kme_cceip2_ob_out_post.tdata [16]);
tran (kme_cceip2_ob_out_post[15], \kme_cceip2_ob_out_post.tdata [15]);
tran (kme_cceip2_ob_out_post[14], \kme_cceip2_ob_out_post.tdata [14]);
tran (kme_cceip2_ob_out_post[13], \kme_cceip2_ob_out_post.tdata [13]);
tran (kme_cceip2_ob_out_post[12], \kme_cceip2_ob_out_post.tdata [12]);
tran (kme_cceip2_ob_out_post[11], \kme_cceip2_ob_out_post.tdata [11]);
tran (kme_cceip2_ob_out_post[10], \kme_cceip2_ob_out_post.tdata [10]);
tran (kme_cceip2_ob_out_post[9], \kme_cceip2_ob_out_post.tdata [9]);
tran (kme_cceip2_ob_out_post[8], \kme_cceip2_ob_out_post.tdata [8]);
tran (kme_cceip2_ob_out_post[7], \kme_cceip2_ob_out_post.tdata [7]);
tran (kme_cceip2_ob_out_post[6], \kme_cceip2_ob_out_post.tdata [6]);
tran (kme_cceip2_ob_out_post[5], \kme_cceip2_ob_out_post.tdata [5]);
tran (kme_cceip2_ob_out_post[4], \kme_cceip2_ob_out_post.tdata [4]);
tran (kme_cceip2_ob_out_post[3], \kme_cceip2_ob_out_post.tdata [3]);
tran (kme_cceip2_ob_out_post[2], \kme_cceip2_ob_out_post.tdata [2]);
tran (kme_cceip2_ob_out_post[1], \kme_cceip2_ob_out_post.tdata [1]);
tran (kme_cceip2_ob_out_post[0], \kme_cceip2_ob_out_post.tdata [0]);
tran (kme_cceip3_ob_out_post[82], \kme_cceip3_ob_out_post.tvalid );
tran (kme_cceip3_ob_out_post[81], \kme_cceip3_ob_out_post.tlast );
tran (kme_cceip3_ob_out_post[80], \kme_cceip3_ob_out_post.tid [0]);
tran (kme_cceip3_ob_out_post[79], \kme_cceip3_ob_out_post.tstrb [7]);
tran (kme_cceip3_ob_out_post[78], \kme_cceip3_ob_out_post.tstrb [6]);
tran (kme_cceip3_ob_out_post[77], \kme_cceip3_ob_out_post.tstrb [5]);
tran (kme_cceip3_ob_out_post[76], \kme_cceip3_ob_out_post.tstrb [4]);
tran (kme_cceip3_ob_out_post[75], \kme_cceip3_ob_out_post.tstrb [3]);
tran (kme_cceip3_ob_out_post[74], \kme_cceip3_ob_out_post.tstrb [2]);
tran (kme_cceip3_ob_out_post[73], \kme_cceip3_ob_out_post.tstrb [1]);
tran (kme_cceip3_ob_out_post[72], \kme_cceip3_ob_out_post.tstrb [0]);
tran (kme_cceip3_ob_out_post[71], \kme_cceip3_ob_out_post.tuser [7]);
tran (kme_cceip3_ob_out_post[70], \kme_cceip3_ob_out_post.tuser [6]);
tran (kme_cceip3_ob_out_post[69], \kme_cceip3_ob_out_post.tuser [5]);
tran (kme_cceip3_ob_out_post[68], \kme_cceip3_ob_out_post.tuser [4]);
tran (kme_cceip3_ob_out_post[67], \kme_cceip3_ob_out_post.tuser [3]);
tran (kme_cceip3_ob_out_post[66], \kme_cceip3_ob_out_post.tuser [2]);
tran (kme_cceip3_ob_out_post[65], \kme_cceip3_ob_out_post.tuser [1]);
tran (kme_cceip3_ob_out_post[64], \kme_cceip3_ob_out_post.tuser [0]);
tran (kme_cceip3_ob_out_post[63], \kme_cceip3_ob_out_post.tdata [63]);
tran (kme_cceip3_ob_out_post[62], \kme_cceip3_ob_out_post.tdata [62]);
tran (kme_cceip3_ob_out_post[61], \kme_cceip3_ob_out_post.tdata [61]);
tran (kme_cceip3_ob_out_post[60], \kme_cceip3_ob_out_post.tdata [60]);
tran (kme_cceip3_ob_out_post[59], \kme_cceip3_ob_out_post.tdata [59]);
tran (kme_cceip3_ob_out_post[58], \kme_cceip3_ob_out_post.tdata [58]);
tran (kme_cceip3_ob_out_post[57], \kme_cceip3_ob_out_post.tdata [57]);
tran (kme_cceip3_ob_out_post[56], \kme_cceip3_ob_out_post.tdata [56]);
tran (kme_cceip3_ob_out_post[55], \kme_cceip3_ob_out_post.tdata [55]);
tran (kme_cceip3_ob_out_post[54], \kme_cceip3_ob_out_post.tdata [54]);
tran (kme_cceip3_ob_out_post[53], \kme_cceip3_ob_out_post.tdata [53]);
tran (kme_cceip3_ob_out_post[52], \kme_cceip3_ob_out_post.tdata [52]);
tran (kme_cceip3_ob_out_post[51], \kme_cceip3_ob_out_post.tdata [51]);
tran (kme_cceip3_ob_out_post[50], \kme_cceip3_ob_out_post.tdata [50]);
tran (kme_cceip3_ob_out_post[49], \kme_cceip3_ob_out_post.tdata [49]);
tran (kme_cceip3_ob_out_post[48], \kme_cceip3_ob_out_post.tdata [48]);
tran (kme_cceip3_ob_out_post[47], \kme_cceip3_ob_out_post.tdata [47]);
tran (kme_cceip3_ob_out_post[46], \kme_cceip3_ob_out_post.tdata [46]);
tran (kme_cceip3_ob_out_post[45], \kme_cceip3_ob_out_post.tdata [45]);
tran (kme_cceip3_ob_out_post[44], \kme_cceip3_ob_out_post.tdata [44]);
tran (kme_cceip3_ob_out_post[43], \kme_cceip3_ob_out_post.tdata [43]);
tran (kme_cceip3_ob_out_post[42], \kme_cceip3_ob_out_post.tdata [42]);
tran (kme_cceip3_ob_out_post[41], \kme_cceip3_ob_out_post.tdata [41]);
tran (kme_cceip3_ob_out_post[40], \kme_cceip3_ob_out_post.tdata [40]);
tran (kme_cceip3_ob_out_post[39], \kme_cceip3_ob_out_post.tdata [39]);
tran (kme_cceip3_ob_out_post[38], \kme_cceip3_ob_out_post.tdata [38]);
tran (kme_cceip3_ob_out_post[37], \kme_cceip3_ob_out_post.tdata [37]);
tran (kme_cceip3_ob_out_post[36], \kme_cceip3_ob_out_post.tdata [36]);
tran (kme_cceip3_ob_out_post[35], \kme_cceip3_ob_out_post.tdata [35]);
tran (kme_cceip3_ob_out_post[34], \kme_cceip3_ob_out_post.tdata [34]);
tran (kme_cceip3_ob_out_post[33], \kme_cceip3_ob_out_post.tdata [33]);
tran (kme_cceip3_ob_out_post[32], \kme_cceip3_ob_out_post.tdata [32]);
tran (kme_cceip3_ob_out_post[31], \kme_cceip3_ob_out_post.tdata [31]);
tran (kme_cceip3_ob_out_post[30], \kme_cceip3_ob_out_post.tdata [30]);
tran (kme_cceip3_ob_out_post[29], \kme_cceip3_ob_out_post.tdata [29]);
tran (kme_cceip3_ob_out_post[28], \kme_cceip3_ob_out_post.tdata [28]);
tran (kme_cceip3_ob_out_post[27], \kme_cceip3_ob_out_post.tdata [27]);
tran (kme_cceip3_ob_out_post[26], \kme_cceip3_ob_out_post.tdata [26]);
tran (kme_cceip3_ob_out_post[25], \kme_cceip3_ob_out_post.tdata [25]);
tran (kme_cceip3_ob_out_post[24], \kme_cceip3_ob_out_post.tdata [24]);
tran (kme_cceip3_ob_out_post[23], \kme_cceip3_ob_out_post.tdata [23]);
tran (kme_cceip3_ob_out_post[22], \kme_cceip3_ob_out_post.tdata [22]);
tran (kme_cceip3_ob_out_post[21], \kme_cceip3_ob_out_post.tdata [21]);
tran (kme_cceip3_ob_out_post[20], \kme_cceip3_ob_out_post.tdata [20]);
tran (kme_cceip3_ob_out_post[19], \kme_cceip3_ob_out_post.tdata [19]);
tran (kme_cceip3_ob_out_post[18], \kme_cceip3_ob_out_post.tdata [18]);
tran (kme_cceip3_ob_out_post[17], \kme_cceip3_ob_out_post.tdata [17]);
tran (kme_cceip3_ob_out_post[16], \kme_cceip3_ob_out_post.tdata [16]);
tran (kme_cceip3_ob_out_post[15], \kme_cceip3_ob_out_post.tdata [15]);
tran (kme_cceip3_ob_out_post[14], \kme_cceip3_ob_out_post.tdata [14]);
tran (kme_cceip3_ob_out_post[13], \kme_cceip3_ob_out_post.tdata [13]);
tran (kme_cceip3_ob_out_post[12], \kme_cceip3_ob_out_post.tdata [12]);
tran (kme_cceip3_ob_out_post[11], \kme_cceip3_ob_out_post.tdata [11]);
tran (kme_cceip3_ob_out_post[10], \kme_cceip3_ob_out_post.tdata [10]);
tran (kme_cceip3_ob_out_post[9], \kme_cceip3_ob_out_post.tdata [9]);
tran (kme_cceip3_ob_out_post[8], \kme_cceip3_ob_out_post.tdata [8]);
tran (kme_cceip3_ob_out_post[7], \kme_cceip3_ob_out_post.tdata [7]);
tran (kme_cceip3_ob_out_post[6], \kme_cceip3_ob_out_post.tdata [6]);
tran (kme_cceip3_ob_out_post[5], \kme_cceip3_ob_out_post.tdata [5]);
tran (kme_cceip3_ob_out_post[4], \kme_cceip3_ob_out_post.tdata [4]);
tran (kme_cceip3_ob_out_post[3], \kme_cceip3_ob_out_post.tdata [3]);
tran (kme_cceip3_ob_out_post[2], \kme_cceip3_ob_out_post.tdata [2]);
tran (kme_cceip3_ob_out_post[1], \kme_cceip3_ob_out_post.tdata [1]);
tran (kme_cceip3_ob_out_post[0], \kme_cceip3_ob_out_post.tdata [0]);
tran (kme_cddip0_ob_out_post[82], \kme_cddip0_ob_out_post.tvalid );
tran (kme_cddip0_ob_out_post[81], \kme_cddip0_ob_out_post.tlast );
tran (kme_cddip0_ob_out_post[80], \kme_cddip0_ob_out_post.tid [0]);
tran (kme_cddip0_ob_out_post[79], \kme_cddip0_ob_out_post.tstrb [7]);
tran (kme_cddip0_ob_out_post[78], \kme_cddip0_ob_out_post.tstrb [6]);
tran (kme_cddip0_ob_out_post[77], \kme_cddip0_ob_out_post.tstrb [5]);
tran (kme_cddip0_ob_out_post[76], \kme_cddip0_ob_out_post.tstrb [4]);
tran (kme_cddip0_ob_out_post[75], \kme_cddip0_ob_out_post.tstrb [3]);
tran (kme_cddip0_ob_out_post[74], \kme_cddip0_ob_out_post.tstrb [2]);
tran (kme_cddip0_ob_out_post[73], \kme_cddip0_ob_out_post.tstrb [1]);
tran (kme_cddip0_ob_out_post[72], \kme_cddip0_ob_out_post.tstrb [0]);
tran (kme_cddip0_ob_out_post[71], \kme_cddip0_ob_out_post.tuser [7]);
tran (kme_cddip0_ob_out_post[70], \kme_cddip0_ob_out_post.tuser [6]);
tran (kme_cddip0_ob_out_post[69], \kme_cddip0_ob_out_post.tuser [5]);
tran (kme_cddip0_ob_out_post[68], \kme_cddip0_ob_out_post.tuser [4]);
tran (kme_cddip0_ob_out_post[67], \kme_cddip0_ob_out_post.tuser [3]);
tran (kme_cddip0_ob_out_post[66], \kme_cddip0_ob_out_post.tuser [2]);
tran (kme_cddip0_ob_out_post[65], \kme_cddip0_ob_out_post.tuser [1]);
tran (kme_cddip0_ob_out_post[64], \kme_cddip0_ob_out_post.tuser [0]);
tran (kme_cddip0_ob_out_post[63], \kme_cddip0_ob_out_post.tdata [63]);
tran (kme_cddip0_ob_out_post[62], \kme_cddip0_ob_out_post.tdata [62]);
tran (kme_cddip0_ob_out_post[61], \kme_cddip0_ob_out_post.tdata [61]);
tran (kme_cddip0_ob_out_post[60], \kme_cddip0_ob_out_post.tdata [60]);
tran (kme_cddip0_ob_out_post[59], \kme_cddip0_ob_out_post.tdata [59]);
tran (kme_cddip0_ob_out_post[58], \kme_cddip0_ob_out_post.tdata [58]);
tran (kme_cddip0_ob_out_post[57], \kme_cddip0_ob_out_post.tdata [57]);
tran (kme_cddip0_ob_out_post[56], \kme_cddip0_ob_out_post.tdata [56]);
tran (kme_cddip0_ob_out_post[55], \kme_cddip0_ob_out_post.tdata [55]);
tran (kme_cddip0_ob_out_post[54], \kme_cddip0_ob_out_post.tdata [54]);
tran (kme_cddip0_ob_out_post[53], \kme_cddip0_ob_out_post.tdata [53]);
tran (kme_cddip0_ob_out_post[52], \kme_cddip0_ob_out_post.tdata [52]);
tran (kme_cddip0_ob_out_post[51], \kme_cddip0_ob_out_post.tdata [51]);
tran (kme_cddip0_ob_out_post[50], \kme_cddip0_ob_out_post.tdata [50]);
tran (kme_cddip0_ob_out_post[49], \kme_cddip0_ob_out_post.tdata [49]);
tran (kme_cddip0_ob_out_post[48], \kme_cddip0_ob_out_post.tdata [48]);
tran (kme_cddip0_ob_out_post[47], \kme_cddip0_ob_out_post.tdata [47]);
tran (kme_cddip0_ob_out_post[46], \kme_cddip0_ob_out_post.tdata [46]);
tran (kme_cddip0_ob_out_post[45], \kme_cddip0_ob_out_post.tdata [45]);
tran (kme_cddip0_ob_out_post[44], \kme_cddip0_ob_out_post.tdata [44]);
tran (kme_cddip0_ob_out_post[43], \kme_cddip0_ob_out_post.tdata [43]);
tran (kme_cddip0_ob_out_post[42], \kme_cddip0_ob_out_post.tdata [42]);
tran (kme_cddip0_ob_out_post[41], \kme_cddip0_ob_out_post.tdata [41]);
tran (kme_cddip0_ob_out_post[40], \kme_cddip0_ob_out_post.tdata [40]);
tran (kme_cddip0_ob_out_post[39], \kme_cddip0_ob_out_post.tdata [39]);
tran (kme_cddip0_ob_out_post[38], \kme_cddip0_ob_out_post.tdata [38]);
tran (kme_cddip0_ob_out_post[37], \kme_cddip0_ob_out_post.tdata [37]);
tran (kme_cddip0_ob_out_post[36], \kme_cddip0_ob_out_post.tdata [36]);
tran (kme_cddip0_ob_out_post[35], \kme_cddip0_ob_out_post.tdata [35]);
tran (kme_cddip0_ob_out_post[34], \kme_cddip0_ob_out_post.tdata [34]);
tran (kme_cddip0_ob_out_post[33], \kme_cddip0_ob_out_post.tdata [33]);
tran (kme_cddip0_ob_out_post[32], \kme_cddip0_ob_out_post.tdata [32]);
tran (kme_cddip0_ob_out_post[31], \kme_cddip0_ob_out_post.tdata [31]);
tran (kme_cddip0_ob_out_post[30], \kme_cddip0_ob_out_post.tdata [30]);
tran (kme_cddip0_ob_out_post[29], \kme_cddip0_ob_out_post.tdata [29]);
tran (kme_cddip0_ob_out_post[28], \kme_cddip0_ob_out_post.tdata [28]);
tran (kme_cddip0_ob_out_post[27], \kme_cddip0_ob_out_post.tdata [27]);
tran (kme_cddip0_ob_out_post[26], \kme_cddip0_ob_out_post.tdata [26]);
tran (kme_cddip0_ob_out_post[25], \kme_cddip0_ob_out_post.tdata [25]);
tran (kme_cddip0_ob_out_post[24], \kme_cddip0_ob_out_post.tdata [24]);
tran (kme_cddip0_ob_out_post[23], \kme_cddip0_ob_out_post.tdata [23]);
tran (kme_cddip0_ob_out_post[22], \kme_cddip0_ob_out_post.tdata [22]);
tran (kme_cddip0_ob_out_post[21], \kme_cddip0_ob_out_post.tdata [21]);
tran (kme_cddip0_ob_out_post[20], \kme_cddip0_ob_out_post.tdata [20]);
tran (kme_cddip0_ob_out_post[19], \kme_cddip0_ob_out_post.tdata [19]);
tran (kme_cddip0_ob_out_post[18], \kme_cddip0_ob_out_post.tdata [18]);
tran (kme_cddip0_ob_out_post[17], \kme_cddip0_ob_out_post.tdata [17]);
tran (kme_cddip0_ob_out_post[16], \kme_cddip0_ob_out_post.tdata [16]);
tran (kme_cddip0_ob_out_post[15], \kme_cddip0_ob_out_post.tdata [15]);
tran (kme_cddip0_ob_out_post[14], \kme_cddip0_ob_out_post.tdata [14]);
tran (kme_cddip0_ob_out_post[13], \kme_cddip0_ob_out_post.tdata [13]);
tran (kme_cddip0_ob_out_post[12], \kme_cddip0_ob_out_post.tdata [12]);
tran (kme_cddip0_ob_out_post[11], \kme_cddip0_ob_out_post.tdata [11]);
tran (kme_cddip0_ob_out_post[10], \kme_cddip0_ob_out_post.tdata [10]);
tran (kme_cddip0_ob_out_post[9], \kme_cddip0_ob_out_post.tdata [9]);
tran (kme_cddip0_ob_out_post[8], \kme_cddip0_ob_out_post.tdata [8]);
tran (kme_cddip0_ob_out_post[7], \kme_cddip0_ob_out_post.tdata [7]);
tran (kme_cddip0_ob_out_post[6], \kme_cddip0_ob_out_post.tdata [6]);
tran (kme_cddip0_ob_out_post[5], \kme_cddip0_ob_out_post.tdata [5]);
tran (kme_cddip0_ob_out_post[4], \kme_cddip0_ob_out_post.tdata [4]);
tran (kme_cddip0_ob_out_post[3], \kme_cddip0_ob_out_post.tdata [3]);
tran (kme_cddip0_ob_out_post[2], \kme_cddip0_ob_out_post.tdata [2]);
tran (kme_cddip0_ob_out_post[1], \kme_cddip0_ob_out_post.tdata [1]);
tran (kme_cddip0_ob_out_post[0], \kme_cddip0_ob_out_post.tdata [0]);
tran (kme_cddip1_ob_out_post[82], \kme_cddip1_ob_out_post.tvalid );
tran (kme_cddip1_ob_out_post[81], \kme_cddip1_ob_out_post.tlast );
tran (kme_cddip1_ob_out_post[80], \kme_cddip1_ob_out_post.tid [0]);
tran (kme_cddip1_ob_out_post[79], \kme_cddip1_ob_out_post.tstrb [7]);
tran (kme_cddip1_ob_out_post[78], \kme_cddip1_ob_out_post.tstrb [6]);
tran (kme_cddip1_ob_out_post[77], \kme_cddip1_ob_out_post.tstrb [5]);
tran (kme_cddip1_ob_out_post[76], \kme_cddip1_ob_out_post.tstrb [4]);
tran (kme_cddip1_ob_out_post[75], \kme_cddip1_ob_out_post.tstrb [3]);
tran (kme_cddip1_ob_out_post[74], \kme_cddip1_ob_out_post.tstrb [2]);
tran (kme_cddip1_ob_out_post[73], \kme_cddip1_ob_out_post.tstrb [1]);
tran (kme_cddip1_ob_out_post[72], \kme_cddip1_ob_out_post.tstrb [0]);
tran (kme_cddip1_ob_out_post[71], \kme_cddip1_ob_out_post.tuser [7]);
tran (kme_cddip1_ob_out_post[70], \kme_cddip1_ob_out_post.tuser [6]);
tran (kme_cddip1_ob_out_post[69], \kme_cddip1_ob_out_post.tuser [5]);
tran (kme_cddip1_ob_out_post[68], \kme_cddip1_ob_out_post.tuser [4]);
tran (kme_cddip1_ob_out_post[67], \kme_cddip1_ob_out_post.tuser [3]);
tran (kme_cddip1_ob_out_post[66], \kme_cddip1_ob_out_post.tuser [2]);
tran (kme_cddip1_ob_out_post[65], \kme_cddip1_ob_out_post.tuser [1]);
tran (kme_cddip1_ob_out_post[64], \kme_cddip1_ob_out_post.tuser [0]);
tran (kme_cddip1_ob_out_post[63], \kme_cddip1_ob_out_post.tdata [63]);
tran (kme_cddip1_ob_out_post[62], \kme_cddip1_ob_out_post.tdata [62]);
tran (kme_cddip1_ob_out_post[61], \kme_cddip1_ob_out_post.tdata [61]);
tran (kme_cddip1_ob_out_post[60], \kme_cddip1_ob_out_post.tdata [60]);
tran (kme_cddip1_ob_out_post[59], \kme_cddip1_ob_out_post.tdata [59]);
tran (kme_cddip1_ob_out_post[58], \kme_cddip1_ob_out_post.tdata [58]);
tran (kme_cddip1_ob_out_post[57], \kme_cddip1_ob_out_post.tdata [57]);
tran (kme_cddip1_ob_out_post[56], \kme_cddip1_ob_out_post.tdata [56]);
tran (kme_cddip1_ob_out_post[55], \kme_cddip1_ob_out_post.tdata [55]);
tran (kme_cddip1_ob_out_post[54], \kme_cddip1_ob_out_post.tdata [54]);
tran (kme_cddip1_ob_out_post[53], \kme_cddip1_ob_out_post.tdata [53]);
tran (kme_cddip1_ob_out_post[52], \kme_cddip1_ob_out_post.tdata [52]);
tran (kme_cddip1_ob_out_post[51], \kme_cddip1_ob_out_post.tdata [51]);
tran (kme_cddip1_ob_out_post[50], \kme_cddip1_ob_out_post.tdata [50]);
tran (kme_cddip1_ob_out_post[49], \kme_cddip1_ob_out_post.tdata [49]);
tran (kme_cddip1_ob_out_post[48], \kme_cddip1_ob_out_post.tdata [48]);
tran (kme_cddip1_ob_out_post[47], \kme_cddip1_ob_out_post.tdata [47]);
tran (kme_cddip1_ob_out_post[46], \kme_cddip1_ob_out_post.tdata [46]);
tran (kme_cddip1_ob_out_post[45], \kme_cddip1_ob_out_post.tdata [45]);
tran (kme_cddip1_ob_out_post[44], \kme_cddip1_ob_out_post.tdata [44]);
tran (kme_cddip1_ob_out_post[43], \kme_cddip1_ob_out_post.tdata [43]);
tran (kme_cddip1_ob_out_post[42], \kme_cddip1_ob_out_post.tdata [42]);
tran (kme_cddip1_ob_out_post[41], \kme_cddip1_ob_out_post.tdata [41]);
tran (kme_cddip1_ob_out_post[40], \kme_cddip1_ob_out_post.tdata [40]);
tran (kme_cddip1_ob_out_post[39], \kme_cddip1_ob_out_post.tdata [39]);
tran (kme_cddip1_ob_out_post[38], \kme_cddip1_ob_out_post.tdata [38]);
tran (kme_cddip1_ob_out_post[37], \kme_cddip1_ob_out_post.tdata [37]);
tran (kme_cddip1_ob_out_post[36], \kme_cddip1_ob_out_post.tdata [36]);
tran (kme_cddip1_ob_out_post[35], \kme_cddip1_ob_out_post.tdata [35]);
tran (kme_cddip1_ob_out_post[34], \kme_cddip1_ob_out_post.tdata [34]);
tran (kme_cddip1_ob_out_post[33], \kme_cddip1_ob_out_post.tdata [33]);
tran (kme_cddip1_ob_out_post[32], \kme_cddip1_ob_out_post.tdata [32]);
tran (kme_cddip1_ob_out_post[31], \kme_cddip1_ob_out_post.tdata [31]);
tran (kme_cddip1_ob_out_post[30], \kme_cddip1_ob_out_post.tdata [30]);
tran (kme_cddip1_ob_out_post[29], \kme_cddip1_ob_out_post.tdata [29]);
tran (kme_cddip1_ob_out_post[28], \kme_cddip1_ob_out_post.tdata [28]);
tran (kme_cddip1_ob_out_post[27], \kme_cddip1_ob_out_post.tdata [27]);
tran (kme_cddip1_ob_out_post[26], \kme_cddip1_ob_out_post.tdata [26]);
tran (kme_cddip1_ob_out_post[25], \kme_cddip1_ob_out_post.tdata [25]);
tran (kme_cddip1_ob_out_post[24], \kme_cddip1_ob_out_post.tdata [24]);
tran (kme_cddip1_ob_out_post[23], \kme_cddip1_ob_out_post.tdata [23]);
tran (kme_cddip1_ob_out_post[22], \kme_cddip1_ob_out_post.tdata [22]);
tran (kme_cddip1_ob_out_post[21], \kme_cddip1_ob_out_post.tdata [21]);
tran (kme_cddip1_ob_out_post[20], \kme_cddip1_ob_out_post.tdata [20]);
tran (kme_cddip1_ob_out_post[19], \kme_cddip1_ob_out_post.tdata [19]);
tran (kme_cddip1_ob_out_post[18], \kme_cddip1_ob_out_post.tdata [18]);
tran (kme_cddip1_ob_out_post[17], \kme_cddip1_ob_out_post.tdata [17]);
tran (kme_cddip1_ob_out_post[16], \kme_cddip1_ob_out_post.tdata [16]);
tran (kme_cddip1_ob_out_post[15], \kme_cddip1_ob_out_post.tdata [15]);
tran (kme_cddip1_ob_out_post[14], \kme_cddip1_ob_out_post.tdata [14]);
tran (kme_cddip1_ob_out_post[13], \kme_cddip1_ob_out_post.tdata [13]);
tran (kme_cddip1_ob_out_post[12], \kme_cddip1_ob_out_post.tdata [12]);
tran (kme_cddip1_ob_out_post[11], \kme_cddip1_ob_out_post.tdata [11]);
tran (kme_cddip1_ob_out_post[10], \kme_cddip1_ob_out_post.tdata [10]);
tran (kme_cddip1_ob_out_post[9], \kme_cddip1_ob_out_post.tdata [9]);
tran (kme_cddip1_ob_out_post[8], \kme_cddip1_ob_out_post.tdata [8]);
tran (kme_cddip1_ob_out_post[7], \kme_cddip1_ob_out_post.tdata [7]);
tran (kme_cddip1_ob_out_post[6], \kme_cddip1_ob_out_post.tdata [6]);
tran (kme_cddip1_ob_out_post[5], \kme_cddip1_ob_out_post.tdata [5]);
tran (kme_cddip1_ob_out_post[4], \kme_cddip1_ob_out_post.tdata [4]);
tran (kme_cddip1_ob_out_post[3], \kme_cddip1_ob_out_post.tdata [3]);
tran (kme_cddip1_ob_out_post[2], \kme_cddip1_ob_out_post.tdata [2]);
tran (kme_cddip1_ob_out_post[1], \kme_cddip1_ob_out_post.tdata [1]);
tran (kme_cddip1_ob_out_post[0], \kme_cddip1_ob_out_post.tdata [0]);
tran (kme_cddip2_ob_out_post[82], \kme_cddip2_ob_out_post.tvalid );
tran (kme_cddip2_ob_out_post[81], \kme_cddip2_ob_out_post.tlast );
tran (kme_cddip2_ob_out_post[80], \kme_cddip2_ob_out_post.tid [0]);
tran (kme_cddip2_ob_out_post[79], \kme_cddip2_ob_out_post.tstrb [7]);
tran (kme_cddip2_ob_out_post[78], \kme_cddip2_ob_out_post.tstrb [6]);
tran (kme_cddip2_ob_out_post[77], \kme_cddip2_ob_out_post.tstrb [5]);
tran (kme_cddip2_ob_out_post[76], \kme_cddip2_ob_out_post.tstrb [4]);
tran (kme_cddip2_ob_out_post[75], \kme_cddip2_ob_out_post.tstrb [3]);
tran (kme_cddip2_ob_out_post[74], \kme_cddip2_ob_out_post.tstrb [2]);
tran (kme_cddip2_ob_out_post[73], \kme_cddip2_ob_out_post.tstrb [1]);
tran (kme_cddip2_ob_out_post[72], \kme_cddip2_ob_out_post.tstrb [0]);
tran (kme_cddip2_ob_out_post[71], \kme_cddip2_ob_out_post.tuser [7]);
tran (kme_cddip2_ob_out_post[70], \kme_cddip2_ob_out_post.tuser [6]);
tran (kme_cddip2_ob_out_post[69], \kme_cddip2_ob_out_post.tuser [5]);
tran (kme_cddip2_ob_out_post[68], \kme_cddip2_ob_out_post.tuser [4]);
tran (kme_cddip2_ob_out_post[67], \kme_cddip2_ob_out_post.tuser [3]);
tran (kme_cddip2_ob_out_post[66], \kme_cddip2_ob_out_post.tuser [2]);
tran (kme_cddip2_ob_out_post[65], \kme_cddip2_ob_out_post.tuser [1]);
tran (kme_cddip2_ob_out_post[64], \kme_cddip2_ob_out_post.tuser [0]);
tran (kme_cddip2_ob_out_post[63], \kme_cddip2_ob_out_post.tdata [63]);
tran (kme_cddip2_ob_out_post[62], \kme_cddip2_ob_out_post.tdata [62]);
tran (kme_cddip2_ob_out_post[61], \kme_cddip2_ob_out_post.tdata [61]);
tran (kme_cddip2_ob_out_post[60], \kme_cddip2_ob_out_post.tdata [60]);
tran (kme_cddip2_ob_out_post[59], \kme_cddip2_ob_out_post.tdata [59]);
tran (kme_cddip2_ob_out_post[58], \kme_cddip2_ob_out_post.tdata [58]);
tran (kme_cddip2_ob_out_post[57], \kme_cddip2_ob_out_post.tdata [57]);
tran (kme_cddip2_ob_out_post[56], \kme_cddip2_ob_out_post.tdata [56]);
tran (kme_cddip2_ob_out_post[55], \kme_cddip2_ob_out_post.tdata [55]);
tran (kme_cddip2_ob_out_post[54], \kme_cddip2_ob_out_post.tdata [54]);
tran (kme_cddip2_ob_out_post[53], \kme_cddip2_ob_out_post.tdata [53]);
tran (kme_cddip2_ob_out_post[52], \kme_cddip2_ob_out_post.tdata [52]);
tran (kme_cddip2_ob_out_post[51], \kme_cddip2_ob_out_post.tdata [51]);
tran (kme_cddip2_ob_out_post[50], \kme_cddip2_ob_out_post.tdata [50]);
tran (kme_cddip2_ob_out_post[49], \kme_cddip2_ob_out_post.tdata [49]);
tran (kme_cddip2_ob_out_post[48], \kme_cddip2_ob_out_post.tdata [48]);
tran (kme_cddip2_ob_out_post[47], \kme_cddip2_ob_out_post.tdata [47]);
tran (kme_cddip2_ob_out_post[46], \kme_cddip2_ob_out_post.tdata [46]);
tran (kme_cddip2_ob_out_post[45], \kme_cddip2_ob_out_post.tdata [45]);
tran (kme_cddip2_ob_out_post[44], \kme_cddip2_ob_out_post.tdata [44]);
tran (kme_cddip2_ob_out_post[43], \kme_cddip2_ob_out_post.tdata [43]);
tran (kme_cddip2_ob_out_post[42], \kme_cddip2_ob_out_post.tdata [42]);
tran (kme_cddip2_ob_out_post[41], \kme_cddip2_ob_out_post.tdata [41]);
tran (kme_cddip2_ob_out_post[40], \kme_cddip2_ob_out_post.tdata [40]);
tran (kme_cddip2_ob_out_post[39], \kme_cddip2_ob_out_post.tdata [39]);
tran (kme_cddip2_ob_out_post[38], \kme_cddip2_ob_out_post.tdata [38]);
tran (kme_cddip2_ob_out_post[37], \kme_cddip2_ob_out_post.tdata [37]);
tran (kme_cddip2_ob_out_post[36], \kme_cddip2_ob_out_post.tdata [36]);
tran (kme_cddip2_ob_out_post[35], \kme_cddip2_ob_out_post.tdata [35]);
tran (kme_cddip2_ob_out_post[34], \kme_cddip2_ob_out_post.tdata [34]);
tran (kme_cddip2_ob_out_post[33], \kme_cddip2_ob_out_post.tdata [33]);
tran (kme_cddip2_ob_out_post[32], \kme_cddip2_ob_out_post.tdata [32]);
tran (kme_cddip2_ob_out_post[31], \kme_cddip2_ob_out_post.tdata [31]);
tran (kme_cddip2_ob_out_post[30], \kme_cddip2_ob_out_post.tdata [30]);
tran (kme_cddip2_ob_out_post[29], \kme_cddip2_ob_out_post.tdata [29]);
tran (kme_cddip2_ob_out_post[28], \kme_cddip2_ob_out_post.tdata [28]);
tran (kme_cddip2_ob_out_post[27], \kme_cddip2_ob_out_post.tdata [27]);
tran (kme_cddip2_ob_out_post[26], \kme_cddip2_ob_out_post.tdata [26]);
tran (kme_cddip2_ob_out_post[25], \kme_cddip2_ob_out_post.tdata [25]);
tran (kme_cddip2_ob_out_post[24], \kme_cddip2_ob_out_post.tdata [24]);
tran (kme_cddip2_ob_out_post[23], \kme_cddip2_ob_out_post.tdata [23]);
tran (kme_cddip2_ob_out_post[22], \kme_cddip2_ob_out_post.tdata [22]);
tran (kme_cddip2_ob_out_post[21], \kme_cddip2_ob_out_post.tdata [21]);
tran (kme_cddip2_ob_out_post[20], \kme_cddip2_ob_out_post.tdata [20]);
tran (kme_cddip2_ob_out_post[19], \kme_cddip2_ob_out_post.tdata [19]);
tran (kme_cddip2_ob_out_post[18], \kme_cddip2_ob_out_post.tdata [18]);
tran (kme_cddip2_ob_out_post[17], \kme_cddip2_ob_out_post.tdata [17]);
tran (kme_cddip2_ob_out_post[16], \kme_cddip2_ob_out_post.tdata [16]);
tran (kme_cddip2_ob_out_post[15], \kme_cddip2_ob_out_post.tdata [15]);
tran (kme_cddip2_ob_out_post[14], \kme_cddip2_ob_out_post.tdata [14]);
tran (kme_cddip2_ob_out_post[13], \kme_cddip2_ob_out_post.tdata [13]);
tran (kme_cddip2_ob_out_post[12], \kme_cddip2_ob_out_post.tdata [12]);
tran (kme_cddip2_ob_out_post[11], \kme_cddip2_ob_out_post.tdata [11]);
tran (kme_cddip2_ob_out_post[10], \kme_cddip2_ob_out_post.tdata [10]);
tran (kme_cddip2_ob_out_post[9], \kme_cddip2_ob_out_post.tdata [9]);
tran (kme_cddip2_ob_out_post[8], \kme_cddip2_ob_out_post.tdata [8]);
tran (kme_cddip2_ob_out_post[7], \kme_cddip2_ob_out_post.tdata [7]);
tran (kme_cddip2_ob_out_post[6], \kme_cddip2_ob_out_post.tdata [6]);
tran (kme_cddip2_ob_out_post[5], \kme_cddip2_ob_out_post.tdata [5]);
tran (kme_cddip2_ob_out_post[4], \kme_cddip2_ob_out_post.tdata [4]);
tran (kme_cddip2_ob_out_post[3], \kme_cddip2_ob_out_post.tdata [3]);
tran (kme_cddip2_ob_out_post[2], \kme_cddip2_ob_out_post.tdata [2]);
tran (kme_cddip2_ob_out_post[1], \kme_cddip2_ob_out_post.tdata [1]);
tran (kme_cddip2_ob_out_post[0], \kme_cddip2_ob_out_post.tdata [0]);
tran (kme_cddip3_ob_out_post[82], \kme_cddip3_ob_out_post.tvalid );
tran (kme_cddip3_ob_out_post[81], \kme_cddip3_ob_out_post.tlast );
tran (kme_cddip3_ob_out_post[80], \kme_cddip3_ob_out_post.tid [0]);
tran (kme_cddip3_ob_out_post[79], \kme_cddip3_ob_out_post.tstrb [7]);
tran (kme_cddip3_ob_out_post[78], \kme_cddip3_ob_out_post.tstrb [6]);
tran (kme_cddip3_ob_out_post[77], \kme_cddip3_ob_out_post.tstrb [5]);
tran (kme_cddip3_ob_out_post[76], \kme_cddip3_ob_out_post.tstrb [4]);
tran (kme_cddip3_ob_out_post[75], \kme_cddip3_ob_out_post.tstrb [3]);
tran (kme_cddip3_ob_out_post[74], \kme_cddip3_ob_out_post.tstrb [2]);
tran (kme_cddip3_ob_out_post[73], \kme_cddip3_ob_out_post.tstrb [1]);
tran (kme_cddip3_ob_out_post[72], \kme_cddip3_ob_out_post.tstrb [0]);
tran (kme_cddip3_ob_out_post[71], \kme_cddip3_ob_out_post.tuser [7]);
tran (kme_cddip3_ob_out_post[70], \kme_cddip3_ob_out_post.tuser [6]);
tran (kme_cddip3_ob_out_post[69], \kme_cddip3_ob_out_post.tuser [5]);
tran (kme_cddip3_ob_out_post[68], \kme_cddip3_ob_out_post.tuser [4]);
tran (kme_cddip3_ob_out_post[67], \kme_cddip3_ob_out_post.tuser [3]);
tran (kme_cddip3_ob_out_post[66], \kme_cddip3_ob_out_post.tuser [2]);
tran (kme_cddip3_ob_out_post[65], \kme_cddip3_ob_out_post.tuser [1]);
tran (kme_cddip3_ob_out_post[64], \kme_cddip3_ob_out_post.tuser [0]);
tran (kme_cddip3_ob_out_post[63], \kme_cddip3_ob_out_post.tdata [63]);
tran (kme_cddip3_ob_out_post[62], \kme_cddip3_ob_out_post.tdata [62]);
tran (kme_cddip3_ob_out_post[61], \kme_cddip3_ob_out_post.tdata [61]);
tran (kme_cddip3_ob_out_post[60], \kme_cddip3_ob_out_post.tdata [60]);
tran (kme_cddip3_ob_out_post[59], \kme_cddip3_ob_out_post.tdata [59]);
tran (kme_cddip3_ob_out_post[58], \kme_cddip3_ob_out_post.tdata [58]);
tran (kme_cddip3_ob_out_post[57], \kme_cddip3_ob_out_post.tdata [57]);
tran (kme_cddip3_ob_out_post[56], \kme_cddip3_ob_out_post.tdata [56]);
tran (kme_cddip3_ob_out_post[55], \kme_cddip3_ob_out_post.tdata [55]);
tran (kme_cddip3_ob_out_post[54], \kme_cddip3_ob_out_post.tdata [54]);
tran (kme_cddip3_ob_out_post[53], \kme_cddip3_ob_out_post.tdata [53]);
tran (kme_cddip3_ob_out_post[52], \kme_cddip3_ob_out_post.tdata [52]);
tran (kme_cddip3_ob_out_post[51], \kme_cddip3_ob_out_post.tdata [51]);
tran (kme_cddip3_ob_out_post[50], \kme_cddip3_ob_out_post.tdata [50]);
tran (kme_cddip3_ob_out_post[49], \kme_cddip3_ob_out_post.tdata [49]);
tran (kme_cddip3_ob_out_post[48], \kme_cddip3_ob_out_post.tdata [48]);
tran (kme_cddip3_ob_out_post[47], \kme_cddip3_ob_out_post.tdata [47]);
tran (kme_cddip3_ob_out_post[46], \kme_cddip3_ob_out_post.tdata [46]);
tran (kme_cddip3_ob_out_post[45], \kme_cddip3_ob_out_post.tdata [45]);
tran (kme_cddip3_ob_out_post[44], \kme_cddip3_ob_out_post.tdata [44]);
tran (kme_cddip3_ob_out_post[43], \kme_cddip3_ob_out_post.tdata [43]);
tran (kme_cddip3_ob_out_post[42], \kme_cddip3_ob_out_post.tdata [42]);
tran (kme_cddip3_ob_out_post[41], \kme_cddip3_ob_out_post.tdata [41]);
tran (kme_cddip3_ob_out_post[40], \kme_cddip3_ob_out_post.tdata [40]);
tran (kme_cddip3_ob_out_post[39], \kme_cddip3_ob_out_post.tdata [39]);
tran (kme_cddip3_ob_out_post[38], \kme_cddip3_ob_out_post.tdata [38]);
tran (kme_cddip3_ob_out_post[37], \kme_cddip3_ob_out_post.tdata [37]);
tran (kme_cddip3_ob_out_post[36], \kme_cddip3_ob_out_post.tdata [36]);
tran (kme_cddip3_ob_out_post[35], \kme_cddip3_ob_out_post.tdata [35]);
tran (kme_cddip3_ob_out_post[34], \kme_cddip3_ob_out_post.tdata [34]);
tran (kme_cddip3_ob_out_post[33], \kme_cddip3_ob_out_post.tdata [33]);
tran (kme_cddip3_ob_out_post[32], \kme_cddip3_ob_out_post.tdata [32]);
tran (kme_cddip3_ob_out_post[31], \kme_cddip3_ob_out_post.tdata [31]);
tran (kme_cddip3_ob_out_post[30], \kme_cddip3_ob_out_post.tdata [30]);
tran (kme_cddip3_ob_out_post[29], \kme_cddip3_ob_out_post.tdata [29]);
tran (kme_cddip3_ob_out_post[28], \kme_cddip3_ob_out_post.tdata [28]);
tran (kme_cddip3_ob_out_post[27], \kme_cddip3_ob_out_post.tdata [27]);
tran (kme_cddip3_ob_out_post[26], \kme_cddip3_ob_out_post.tdata [26]);
tran (kme_cddip3_ob_out_post[25], \kme_cddip3_ob_out_post.tdata [25]);
tran (kme_cddip3_ob_out_post[24], \kme_cddip3_ob_out_post.tdata [24]);
tran (kme_cddip3_ob_out_post[23], \kme_cddip3_ob_out_post.tdata [23]);
tran (kme_cddip3_ob_out_post[22], \kme_cddip3_ob_out_post.tdata [22]);
tran (kme_cddip3_ob_out_post[21], \kme_cddip3_ob_out_post.tdata [21]);
tran (kme_cddip3_ob_out_post[20], \kme_cddip3_ob_out_post.tdata [20]);
tran (kme_cddip3_ob_out_post[19], \kme_cddip3_ob_out_post.tdata [19]);
tran (kme_cddip3_ob_out_post[18], \kme_cddip3_ob_out_post.tdata [18]);
tran (kme_cddip3_ob_out_post[17], \kme_cddip3_ob_out_post.tdata [17]);
tran (kme_cddip3_ob_out_post[16], \kme_cddip3_ob_out_post.tdata [16]);
tran (kme_cddip3_ob_out_post[15], \kme_cddip3_ob_out_post.tdata [15]);
tran (kme_cddip3_ob_out_post[14], \kme_cddip3_ob_out_post.tdata [14]);
tran (kme_cddip3_ob_out_post[13], \kme_cddip3_ob_out_post.tdata [13]);
tran (kme_cddip3_ob_out_post[12], \kme_cddip3_ob_out_post.tdata [12]);
tran (kme_cddip3_ob_out_post[11], \kme_cddip3_ob_out_post.tdata [11]);
tran (kme_cddip3_ob_out_post[10], \kme_cddip3_ob_out_post.tdata [10]);
tran (kme_cddip3_ob_out_post[9], \kme_cddip3_ob_out_post.tdata [9]);
tran (kme_cddip3_ob_out_post[8], \kme_cddip3_ob_out_post.tdata [8]);
tran (kme_cddip3_ob_out_post[7], \kme_cddip3_ob_out_post.tdata [7]);
tran (kme_cddip3_ob_out_post[6], \kme_cddip3_ob_out_post.tdata [6]);
tran (kme_cddip3_ob_out_post[5], \kme_cddip3_ob_out_post.tdata [5]);
tran (kme_cddip3_ob_out_post[4], \kme_cddip3_ob_out_post.tdata [4]);
tran (kme_cddip3_ob_out_post[3], \kme_cddip3_ob_out_post.tdata [3]);
tran (kme_cddip3_ob_out_post[2], \kme_cddip3_ob_out_post.tdata [2]);
tran (kme_cddip3_ob_out_post[1], \kme_cddip3_ob_out_post.tdata [1]);
tran (kme_cddip3_ob_out_post[0], \kme_cddip3_ob_out_post.tdata [0]);
tran (cceip0_out_ia_status[16], \cceip0_out_ia_status.r.part0 [16]);
tran (cceip0_out_ia_status[16], \cceip0_out_ia_status.f.code [2]);
tran (cceip0_out_ia_status[15], \cceip0_out_ia_status.r.part0 [15]);
tran (cceip0_out_ia_status[15], \cceip0_out_ia_status.f.code [1]);
tran (cceip0_out_ia_status[14], \cceip0_out_ia_status.r.part0 [14]);
tran (cceip0_out_ia_status[14], \cceip0_out_ia_status.f.code [0]);
tran (cceip0_out_ia_status[13], \cceip0_out_ia_status.r.part0 [13]);
tran (cceip0_out_ia_status[13], \cceip0_out_ia_status.f.datawords [4]);
tran (cceip0_out_ia_status[12], \cceip0_out_ia_status.r.part0 [12]);
tran (cceip0_out_ia_status[12], \cceip0_out_ia_status.f.datawords [3]);
tran (cceip0_out_ia_status[11], \cceip0_out_ia_status.r.part0 [11]);
tran (cceip0_out_ia_status[11], \cceip0_out_ia_status.f.datawords [2]);
tran (cceip0_out_ia_status[10], \cceip0_out_ia_status.r.part0 [10]);
tran (cceip0_out_ia_status[10], \cceip0_out_ia_status.f.datawords [1]);
tran (cceip0_out_ia_status[9], \cceip0_out_ia_status.r.part0 [9]);
tran (cceip0_out_ia_status[9], \cceip0_out_ia_status.f.datawords [0]);
tran (cceip0_out_ia_status[8], \cceip0_out_ia_status.r.part0 [8]);
tran (cceip0_out_ia_status[8], \cceip0_out_ia_status.f.addr [8]);
tran (cceip0_out_ia_status[7], \cceip0_out_ia_status.r.part0 [7]);
tran (cceip0_out_ia_status[7], \cceip0_out_ia_status.f.addr [7]);
tran (cceip0_out_ia_status[6], \cceip0_out_ia_status.r.part0 [6]);
tran (cceip0_out_ia_status[6], \cceip0_out_ia_status.f.addr [6]);
tran (cceip0_out_ia_status[5], \cceip0_out_ia_status.r.part0 [5]);
tran (cceip0_out_ia_status[5], \cceip0_out_ia_status.f.addr [5]);
tran (cceip0_out_ia_status[4], \cceip0_out_ia_status.r.part0 [4]);
tran (cceip0_out_ia_status[4], \cceip0_out_ia_status.f.addr [4]);
tran (cceip0_out_ia_status[3], \cceip0_out_ia_status.r.part0 [3]);
tran (cceip0_out_ia_status[3], \cceip0_out_ia_status.f.addr [3]);
tran (cceip0_out_ia_status[2], \cceip0_out_ia_status.r.part0 [2]);
tran (cceip0_out_ia_status[2], \cceip0_out_ia_status.f.addr [2]);
tran (cceip0_out_ia_status[1], \cceip0_out_ia_status.r.part0 [1]);
tran (cceip0_out_ia_status[1], \cceip0_out_ia_status.f.addr [1]);
tran (cceip0_out_ia_status[0], \cceip0_out_ia_status.r.part0 [0]);
tran (cceip0_out_ia_status[0], \cceip0_out_ia_status.f.addr [0]);
tran (cceip0_out_ia_capability[15], \cceip0_out_ia_capability.r.part0 [15]);
tran (cceip0_out_ia_capability[15], \cceip0_out_ia_capability.f.ack_error );
tran (cceip0_out_ia_capability[14], \cceip0_out_ia_capability.r.part0 [14]);
tran (cceip0_out_ia_capability[14], \cceip0_out_ia_capability.f.sim_tmo );
tran (cceip0_out_ia_capability[13], \cceip0_out_ia_capability.r.part0 [13]);
tran (cceip0_out_ia_capability[13], \cceip0_out_ia_capability.f.reserved_op [3]);
tran (cceip0_out_ia_capability[12], \cceip0_out_ia_capability.r.part0 [12]);
tran (cceip0_out_ia_capability[12], \cceip0_out_ia_capability.f.reserved_op [2]);
tran (cceip0_out_ia_capability[11], \cceip0_out_ia_capability.r.part0 [11]);
tran (cceip0_out_ia_capability[11], \cceip0_out_ia_capability.f.reserved_op [1]);
tran (cceip0_out_ia_capability[10], \cceip0_out_ia_capability.r.part0 [10]);
tran (cceip0_out_ia_capability[10], \cceip0_out_ia_capability.f.reserved_op [0]);
tran (cceip0_out_ia_capability[9], \cceip0_out_ia_capability.r.part0 [9]);
tran (cceip0_out_ia_capability[9], \cceip0_out_ia_capability.f.compare );
tran (cceip0_out_ia_capability[8], \cceip0_out_ia_capability.r.part0 [8]);
tran (cceip0_out_ia_capability[8], \cceip0_out_ia_capability.f.set_init_start );
tran (cceip0_out_ia_capability[7], \cceip0_out_ia_capability.r.part0 [7]);
tran (cceip0_out_ia_capability[7], \cceip0_out_ia_capability.f.initialize_inc );
tran (cceip0_out_ia_capability[6], \cceip0_out_ia_capability.r.part0 [6]);
tran (cceip0_out_ia_capability[6], \cceip0_out_ia_capability.f.initialize );
tran (cceip0_out_ia_capability[5], \cceip0_out_ia_capability.r.part0 [5]);
tran (cceip0_out_ia_capability[5], \cceip0_out_ia_capability.f.reset );
tran (cceip0_out_ia_capability[4], \cceip0_out_ia_capability.r.part0 [4]);
tran (cceip0_out_ia_capability[4], \cceip0_out_ia_capability.f.disabled );
tran (cceip0_out_ia_capability[3], \cceip0_out_ia_capability.r.part0 [3]);
tran (cceip0_out_ia_capability[3], \cceip0_out_ia_capability.f.enable );
tran (cceip0_out_ia_capability[2], \cceip0_out_ia_capability.r.part0 [2]);
tran (cceip0_out_ia_capability[2], \cceip0_out_ia_capability.f.write );
tran (cceip0_out_ia_capability[1], \cceip0_out_ia_capability.r.part0 [1]);
tran (cceip0_out_ia_capability[1], \cceip0_out_ia_capability.f.read );
tran (cceip0_out_ia_capability[0], \cceip0_out_ia_capability.r.part0 [0]);
tran (cceip0_out_ia_capability[0], \cceip0_out_ia_capability.f.nop );
tran (cceip0_out_ia_capability[19], \cceip0_out_ia_capability.r.part0 [19]);
tran (cceip0_out_ia_capability[19], \cceip0_out_ia_capability.f.mem_type [3]);
tran (cceip0_out_ia_capability[18], \cceip0_out_ia_capability.r.part0 [18]);
tran (cceip0_out_ia_capability[18], \cceip0_out_ia_capability.f.mem_type [2]);
tran (cceip0_out_ia_capability[17], \cceip0_out_ia_capability.r.part0 [17]);
tran (cceip0_out_ia_capability[17], \cceip0_out_ia_capability.f.mem_type [1]);
tran (cceip0_out_ia_capability[16], \cceip0_out_ia_capability.r.part0 [16]);
tran (cceip0_out_ia_capability[16], \cceip0_out_ia_capability.f.mem_type [0]);
tran (cceip0_out_ia_rdata[95], \cceip0_out_ia_rdata.r.part2 [31]);
tran (cceip0_out_ia_rdata[95], \cceip0_out_ia_rdata.f.tdata_hi [31]);
tran (cceip0_out_ia_rdata[94], \cceip0_out_ia_rdata.r.part2 [30]);
tran (cceip0_out_ia_rdata[94], \cceip0_out_ia_rdata.f.tdata_hi [30]);
tran (cceip0_out_ia_rdata[93], \cceip0_out_ia_rdata.r.part2 [29]);
tran (cceip0_out_ia_rdata[93], \cceip0_out_ia_rdata.f.tdata_hi [29]);
tran (cceip0_out_ia_rdata[92], \cceip0_out_ia_rdata.r.part2 [28]);
tran (cceip0_out_ia_rdata[92], \cceip0_out_ia_rdata.f.tdata_hi [28]);
tran (cceip0_out_ia_rdata[91], \cceip0_out_ia_rdata.r.part2 [27]);
tran (cceip0_out_ia_rdata[91], \cceip0_out_ia_rdata.f.tdata_hi [27]);
tran (cceip0_out_ia_rdata[90], \cceip0_out_ia_rdata.r.part2 [26]);
tran (cceip0_out_ia_rdata[90], \cceip0_out_ia_rdata.f.tdata_hi [26]);
tran (cceip0_out_ia_rdata[89], \cceip0_out_ia_rdata.r.part2 [25]);
tran (cceip0_out_ia_rdata[89], \cceip0_out_ia_rdata.f.tdata_hi [25]);
tran (cceip0_out_ia_rdata[88], \cceip0_out_ia_rdata.r.part2 [24]);
tran (cceip0_out_ia_rdata[88], \cceip0_out_ia_rdata.f.tdata_hi [24]);
tran (cceip0_out_ia_rdata[87], \cceip0_out_ia_rdata.r.part2 [23]);
tran (cceip0_out_ia_rdata[87], \cceip0_out_ia_rdata.f.tdata_hi [23]);
tran (cceip0_out_ia_rdata[86], \cceip0_out_ia_rdata.r.part2 [22]);
tran (cceip0_out_ia_rdata[86], \cceip0_out_ia_rdata.f.tdata_hi [22]);
tran (cceip0_out_ia_rdata[85], \cceip0_out_ia_rdata.r.part2 [21]);
tran (cceip0_out_ia_rdata[85], \cceip0_out_ia_rdata.f.tdata_hi [21]);
tran (cceip0_out_ia_rdata[84], \cceip0_out_ia_rdata.r.part2 [20]);
tran (cceip0_out_ia_rdata[84], \cceip0_out_ia_rdata.f.tdata_hi [20]);
tran (cceip0_out_ia_rdata[83], \cceip0_out_ia_rdata.r.part2 [19]);
tran (cceip0_out_ia_rdata[83], \cceip0_out_ia_rdata.f.tdata_hi [19]);
tran (cceip0_out_ia_rdata[82], \cceip0_out_ia_rdata.r.part2 [18]);
tran (cceip0_out_ia_rdata[82], \cceip0_out_ia_rdata.f.tdata_hi [18]);
tran (cceip0_out_ia_rdata[81], \cceip0_out_ia_rdata.r.part2 [17]);
tran (cceip0_out_ia_rdata[81], \cceip0_out_ia_rdata.f.tdata_hi [17]);
tran (cceip0_out_ia_rdata[80], \cceip0_out_ia_rdata.r.part2 [16]);
tran (cceip0_out_ia_rdata[80], \cceip0_out_ia_rdata.f.tdata_hi [16]);
tran (cceip0_out_ia_rdata[79], \cceip0_out_ia_rdata.r.part2 [15]);
tran (cceip0_out_ia_rdata[79], \cceip0_out_ia_rdata.f.tdata_hi [15]);
tran (cceip0_out_ia_rdata[78], \cceip0_out_ia_rdata.r.part2 [14]);
tran (cceip0_out_ia_rdata[78], \cceip0_out_ia_rdata.f.tdata_hi [14]);
tran (cceip0_out_ia_rdata[77], \cceip0_out_ia_rdata.r.part2 [13]);
tran (cceip0_out_ia_rdata[77], \cceip0_out_ia_rdata.f.tdata_hi [13]);
tran (cceip0_out_ia_rdata[76], \cceip0_out_ia_rdata.r.part2 [12]);
tran (cceip0_out_ia_rdata[76], \cceip0_out_ia_rdata.f.tdata_hi [12]);
tran (cceip0_out_ia_rdata[75], \cceip0_out_ia_rdata.r.part2 [11]);
tran (cceip0_out_ia_rdata[75], \cceip0_out_ia_rdata.f.tdata_hi [11]);
tran (cceip0_out_ia_rdata[74], \cceip0_out_ia_rdata.r.part2 [10]);
tran (cceip0_out_ia_rdata[74], \cceip0_out_ia_rdata.f.tdata_hi [10]);
tran (cceip0_out_ia_rdata[73], \cceip0_out_ia_rdata.r.part2 [9]);
tran (cceip0_out_ia_rdata[73], \cceip0_out_ia_rdata.f.tdata_hi [9]);
tran (cceip0_out_ia_rdata[72], \cceip0_out_ia_rdata.r.part2 [8]);
tran (cceip0_out_ia_rdata[72], \cceip0_out_ia_rdata.f.tdata_hi [8]);
tran (cceip0_out_ia_rdata[71], \cceip0_out_ia_rdata.r.part2 [7]);
tran (cceip0_out_ia_rdata[71], \cceip0_out_ia_rdata.f.tdata_hi [7]);
tran (cceip0_out_ia_rdata[70], \cceip0_out_ia_rdata.r.part2 [6]);
tran (cceip0_out_ia_rdata[70], \cceip0_out_ia_rdata.f.tdata_hi [6]);
tran (cceip0_out_ia_rdata[69], \cceip0_out_ia_rdata.r.part2 [5]);
tran (cceip0_out_ia_rdata[69], \cceip0_out_ia_rdata.f.tdata_hi [5]);
tran (cceip0_out_ia_rdata[68], \cceip0_out_ia_rdata.r.part2 [4]);
tran (cceip0_out_ia_rdata[68], \cceip0_out_ia_rdata.f.tdata_hi [4]);
tran (cceip0_out_ia_rdata[67], \cceip0_out_ia_rdata.r.part2 [3]);
tran (cceip0_out_ia_rdata[67], \cceip0_out_ia_rdata.f.tdata_hi [3]);
tran (cceip0_out_ia_rdata[66], \cceip0_out_ia_rdata.r.part2 [2]);
tran (cceip0_out_ia_rdata[66], \cceip0_out_ia_rdata.f.tdata_hi [2]);
tran (cceip0_out_ia_rdata[65], \cceip0_out_ia_rdata.r.part2 [1]);
tran (cceip0_out_ia_rdata[65], \cceip0_out_ia_rdata.f.tdata_hi [1]);
tran (cceip0_out_ia_rdata[64], \cceip0_out_ia_rdata.r.part2 [0]);
tran (cceip0_out_ia_rdata[64], \cceip0_out_ia_rdata.f.tdata_hi [0]);
tran (cceip0_out_ia_rdata[63], \cceip0_out_ia_rdata.r.part1 [31]);
tran (cceip0_out_ia_rdata[63], \cceip0_out_ia_rdata.f.tdata_lo [31]);
tran (cceip0_out_ia_rdata[62], \cceip0_out_ia_rdata.r.part1 [30]);
tran (cceip0_out_ia_rdata[62], \cceip0_out_ia_rdata.f.tdata_lo [30]);
tran (cceip0_out_ia_rdata[61], \cceip0_out_ia_rdata.r.part1 [29]);
tran (cceip0_out_ia_rdata[61], \cceip0_out_ia_rdata.f.tdata_lo [29]);
tran (cceip0_out_ia_rdata[60], \cceip0_out_ia_rdata.r.part1 [28]);
tran (cceip0_out_ia_rdata[60], \cceip0_out_ia_rdata.f.tdata_lo [28]);
tran (cceip0_out_ia_rdata[59], \cceip0_out_ia_rdata.r.part1 [27]);
tran (cceip0_out_ia_rdata[59], \cceip0_out_ia_rdata.f.tdata_lo [27]);
tran (cceip0_out_ia_rdata[58], \cceip0_out_ia_rdata.r.part1 [26]);
tran (cceip0_out_ia_rdata[58], \cceip0_out_ia_rdata.f.tdata_lo [26]);
tran (cceip0_out_ia_rdata[57], \cceip0_out_ia_rdata.r.part1 [25]);
tran (cceip0_out_ia_rdata[57], \cceip0_out_ia_rdata.f.tdata_lo [25]);
tran (cceip0_out_ia_rdata[56], \cceip0_out_ia_rdata.r.part1 [24]);
tran (cceip0_out_ia_rdata[56], \cceip0_out_ia_rdata.f.tdata_lo [24]);
tran (cceip0_out_ia_rdata[55], \cceip0_out_ia_rdata.r.part1 [23]);
tran (cceip0_out_ia_rdata[55], \cceip0_out_ia_rdata.f.tdata_lo [23]);
tran (cceip0_out_ia_rdata[54], \cceip0_out_ia_rdata.r.part1 [22]);
tran (cceip0_out_ia_rdata[54], \cceip0_out_ia_rdata.f.tdata_lo [22]);
tran (cceip0_out_ia_rdata[53], \cceip0_out_ia_rdata.r.part1 [21]);
tran (cceip0_out_ia_rdata[53], \cceip0_out_ia_rdata.f.tdata_lo [21]);
tran (cceip0_out_ia_rdata[52], \cceip0_out_ia_rdata.r.part1 [20]);
tran (cceip0_out_ia_rdata[52], \cceip0_out_ia_rdata.f.tdata_lo [20]);
tran (cceip0_out_ia_rdata[51], \cceip0_out_ia_rdata.r.part1 [19]);
tran (cceip0_out_ia_rdata[51], \cceip0_out_ia_rdata.f.tdata_lo [19]);
tran (cceip0_out_ia_rdata[50], \cceip0_out_ia_rdata.r.part1 [18]);
tran (cceip0_out_ia_rdata[50], \cceip0_out_ia_rdata.f.tdata_lo [18]);
tran (cceip0_out_ia_rdata[49], \cceip0_out_ia_rdata.r.part1 [17]);
tran (cceip0_out_ia_rdata[49], \cceip0_out_ia_rdata.f.tdata_lo [17]);
tran (cceip0_out_ia_rdata[48], \cceip0_out_ia_rdata.r.part1 [16]);
tran (cceip0_out_ia_rdata[48], \cceip0_out_ia_rdata.f.tdata_lo [16]);
tran (cceip0_out_ia_rdata[47], \cceip0_out_ia_rdata.r.part1 [15]);
tran (cceip0_out_ia_rdata[47], \cceip0_out_ia_rdata.f.tdata_lo [15]);
tran (cceip0_out_ia_rdata[46], \cceip0_out_ia_rdata.r.part1 [14]);
tran (cceip0_out_ia_rdata[46], \cceip0_out_ia_rdata.f.tdata_lo [14]);
tran (cceip0_out_ia_rdata[45], \cceip0_out_ia_rdata.r.part1 [13]);
tran (cceip0_out_ia_rdata[45], \cceip0_out_ia_rdata.f.tdata_lo [13]);
tran (cceip0_out_ia_rdata[44], \cceip0_out_ia_rdata.r.part1 [12]);
tran (cceip0_out_ia_rdata[44], \cceip0_out_ia_rdata.f.tdata_lo [12]);
tran (cceip0_out_ia_rdata[43], \cceip0_out_ia_rdata.r.part1 [11]);
tran (cceip0_out_ia_rdata[43], \cceip0_out_ia_rdata.f.tdata_lo [11]);
tran (cceip0_out_ia_rdata[42], \cceip0_out_ia_rdata.r.part1 [10]);
tran (cceip0_out_ia_rdata[42], \cceip0_out_ia_rdata.f.tdata_lo [10]);
tran (cceip0_out_ia_rdata[41], \cceip0_out_ia_rdata.r.part1 [9]);
tran (cceip0_out_ia_rdata[41], \cceip0_out_ia_rdata.f.tdata_lo [9]);
tran (cceip0_out_ia_rdata[40], \cceip0_out_ia_rdata.r.part1 [8]);
tran (cceip0_out_ia_rdata[40], \cceip0_out_ia_rdata.f.tdata_lo [8]);
tran (cceip0_out_ia_rdata[39], \cceip0_out_ia_rdata.r.part1 [7]);
tran (cceip0_out_ia_rdata[39], \cceip0_out_ia_rdata.f.tdata_lo [7]);
tran (cceip0_out_ia_rdata[38], \cceip0_out_ia_rdata.r.part1 [6]);
tran (cceip0_out_ia_rdata[38], \cceip0_out_ia_rdata.f.tdata_lo [6]);
tran (cceip0_out_ia_rdata[37], \cceip0_out_ia_rdata.r.part1 [5]);
tran (cceip0_out_ia_rdata[37], \cceip0_out_ia_rdata.f.tdata_lo [5]);
tran (cceip0_out_ia_rdata[36], \cceip0_out_ia_rdata.r.part1 [4]);
tran (cceip0_out_ia_rdata[36], \cceip0_out_ia_rdata.f.tdata_lo [4]);
tran (cceip0_out_ia_rdata[35], \cceip0_out_ia_rdata.r.part1 [3]);
tran (cceip0_out_ia_rdata[35], \cceip0_out_ia_rdata.f.tdata_lo [3]);
tran (cceip0_out_ia_rdata[34], \cceip0_out_ia_rdata.r.part1 [2]);
tran (cceip0_out_ia_rdata[34], \cceip0_out_ia_rdata.f.tdata_lo [2]);
tran (cceip0_out_ia_rdata[33], \cceip0_out_ia_rdata.r.part1 [1]);
tran (cceip0_out_ia_rdata[33], \cceip0_out_ia_rdata.f.tdata_lo [1]);
tran (cceip0_out_ia_rdata[32], \cceip0_out_ia_rdata.r.part1 [0]);
tran (cceip0_out_ia_rdata[32], \cceip0_out_ia_rdata.f.tdata_lo [0]);
tran (cceip0_out_ia_rdata[31], \cceip0_out_ia_rdata.r.part0 [31]);
tran (cceip0_out_ia_rdata[31], \cceip0_out_ia_rdata.f.eob );
tran (cceip0_out_ia_rdata[30], \cceip0_out_ia_rdata.r.part0 [30]);
tran (cceip0_out_ia_rdata[30], \cceip0_out_ia_rdata.f.bytes_vld [7]);
tran (cceip0_out_ia_rdata[29], \cceip0_out_ia_rdata.r.part0 [29]);
tran (cceip0_out_ia_rdata[29], \cceip0_out_ia_rdata.f.bytes_vld [6]);
tran (cceip0_out_ia_rdata[28], \cceip0_out_ia_rdata.r.part0 [28]);
tran (cceip0_out_ia_rdata[28], \cceip0_out_ia_rdata.f.bytes_vld [5]);
tran (cceip0_out_ia_rdata[27], \cceip0_out_ia_rdata.r.part0 [27]);
tran (cceip0_out_ia_rdata[27], \cceip0_out_ia_rdata.f.bytes_vld [4]);
tran (cceip0_out_ia_rdata[26], \cceip0_out_ia_rdata.r.part0 [26]);
tran (cceip0_out_ia_rdata[26], \cceip0_out_ia_rdata.f.bytes_vld [3]);
tran (cceip0_out_ia_rdata[25], \cceip0_out_ia_rdata.r.part0 [25]);
tran (cceip0_out_ia_rdata[25], \cceip0_out_ia_rdata.f.bytes_vld [2]);
tran (cceip0_out_ia_rdata[24], \cceip0_out_ia_rdata.r.part0 [24]);
tran (cceip0_out_ia_rdata[24], \cceip0_out_ia_rdata.f.bytes_vld [1]);
tran (cceip0_out_ia_rdata[23], \cceip0_out_ia_rdata.r.part0 [23]);
tran (cceip0_out_ia_rdata[23], \cceip0_out_ia_rdata.f.bytes_vld [0]);
tran (cceip0_out_ia_rdata[22], \cceip0_out_ia_rdata.r.part0 [22]);
tran (cceip0_out_ia_rdata[22], \cceip0_out_ia_rdata.f.unused1 [7]);
tran (cceip0_out_ia_rdata[21], \cceip0_out_ia_rdata.r.part0 [21]);
tran (cceip0_out_ia_rdata[21], \cceip0_out_ia_rdata.f.unused1 [6]);
tran (cceip0_out_ia_rdata[20], \cceip0_out_ia_rdata.r.part0 [20]);
tran (cceip0_out_ia_rdata[20], \cceip0_out_ia_rdata.f.unused1 [5]);
tran (cceip0_out_ia_rdata[19], \cceip0_out_ia_rdata.r.part0 [19]);
tran (cceip0_out_ia_rdata[19], \cceip0_out_ia_rdata.f.unused1 [4]);
tran (cceip0_out_ia_rdata[18], \cceip0_out_ia_rdata.r.part0 [18]);
tran (cceip0_out_ia_rdata[18], \cceip0_out_ia_rdata.f.unused1 [3]);
tran (cceip0_out_ia_rdata[17], \cceip0_out_ia_rdata.r.part0 [17]);
tran (cceip0_out_ia_rdata[17], \cceip0_out_ia_rdata.f.unused1 [2]);
tran (cceip0_out_ia_rdata[16], \cceip0_out_ia_rdata.r.part0 [16]);
tran (cceip0_out_ia_rdata[16], \cceip0_out_ia_rdata.f.unused1 [1]);
tran (cceip0_out_ia_rdata[15], \cceip0_out_ia_rdata.r.part0 [15]);
tran (cceip0_out_ia_rdata[15], \cceip0_out_ia_rdata.f.unused1 [0]);
tran (cceip0_out_ia_rdata[14], \cceip0_out_ia_rdata.r.part0 [14]);
tran (cceip0_out_ia_rdata[14], \cceip0_out_ia_rdata.f.tid );
tran (cceip0_out_ia_rdata[13], \cceip0_out_ia_rdata.r.part0 [13]);
tran (cceip0_out_ia_rdata[13], \cceip0_out_ia_rdata.f.tuser [7]);
tran (cceip0_out_ia_rdata[12], \cceip0_out_ia_rdata.r.part0 [12]);
tran (cceip0_out_ia_rdata[12], \cceip0_out_ia_rdata.f.tuser [6]);
tran (cceip0_out_ia_rdata[11], \cceip0_out_ia_rdata.r.part0 [11]);
tran (cceip0_out_ia_rdata[11], \cceip0_out_ia_rdata.f.tuser [5]);
tran (cceip0_out_ia_rdata[10], \cceip0_out_ia_rdata.r.part0 [10]);
tran (cceip0_out_ia_rdata[10], \cceip0_out_ia_rdata.f.tuser [4]);
tran (cceip0_out_ia_rdata[9], \cceip0_out_ia_rdata.r.part0 [9]);
tran (cceip0_out_ia_rdata[9], \cceip0_out_ia_rdata.f.tuser [3]);
tran (cceip0_out_ia_rdata[8], \cceip0_out_ia_rdata.r.part0 [8]);
tran (cceip0_out_ia_rdata[8], \cceip0_out_ia_rdata.f.tuser [2]);
tran (cceip0_out_ia_rdata[7], \cceip0_out_ia_rdata.r.part0 [7]);
tran (cceip0_out_ia_rdata[7], \cceip0_out_ia_rdata.f.tuser [1]);
tran (cceip0_out_ia_rdata[6], \cceip0_out_ia_rdata.r.part0 [6]);
tran (cceip0_out_ia_rdata[6], \cceip0_out_ia_rdata.f.tuser [0]);
tran (cceip0_out_ia_rdata[5], \cceip0_out_ia_rdata.r.part0 [5]);
tran (cceip0_out_ia_rdata[5], \cceip0_out_ia_rdata.f.unused0 [5]);
tran (cceip0_out_ia_rdata[4], \cceip0_out_ia_rdata.r.part0 [4]);
tran (cceip0_out_ia_rdata[4], \cceip0_out_ia_rdata.f.unused0 [4]);
tran (cceip0_out_ia_rdata[3], \cceip0_out_ia_rdata.r.part0 [3]);
tran (cceip0_out_ia_rdata[3], \cceip0_out_ia_rdata.f.unused0 [3]);
tran (cceip0_out_ia_rdata[2], \cceip0_out_ia_rdata.r.part0 [2]);
tran (cceip0_out_ia_rdata[2], \cceip0_out_ia_rdata.f.unused0 [2]);
tran (cceip0_out_ia_rdata[1], \cceip0_out_ia_rdata.r.part0 [1]);
tran (cceip0_out_ia_rdata[1], \cceip0_out_ia_rdata.f.unused0 [1]);
tran (cceip0_out_ia_rdata[0], \cceip0_out_ia_rdata.r.part0 [0]);
tran (cceip0_out_ia_rdata[0], \cceip0_out_ia_rdata.f.unused0 [0]);
tran (cceip0_out_im_status[11], \cceip0_out_im_status.r.part0 [11]);
tran (cceip0_out_im_status[11], \cceip0_out_im_status.f.bank_hi );
tran (cceip0_out_im_status[10], \cceip0_out_im_status.r.part0 [10]);
tran (cceip0_out_im_status[10], \cceip0_out_im_status.f.bank_lo );
tran (cceip0_out_im_status[9], \cceip0_out_im_status.r.part0 [9]);
tran (cceip0_out_im_status[9], \cceip0_out_im_status.f.overflow );
tran (cceip0_out_im_status[8], \cceip0_out_im_status.r.part0 [8]);
tran (cceip0_out_im_status[8], \cceip0_out_im_status.f.wr_pointer [8]);
tran (cceip0_out_im_status[7], \cceip0_out_im_status.r.part0 [7]);
tran (cceip0_out_im_status[7], \cceip0_out_im_status.f.wr_pointer [7]);
tran (cceip0_out_im_status[6], \cceip0_out_im_status.r.part0 [6]);
tran (cceip0_out_im_status[6], \cceip0_out_im_status.f.wr_pointer [6]);
tran (cceip0_out_im_status[5], \cceip0_out_im_status.r.part0 [5]);
tran (cceip0_out_im_status[5], \cceip0_out_im_status.f.wr_pointer [5]);
tran (cceip0_out_im_status[4], \cceip0_out_im_status.r.part0 [4]);
tran (cceip0_out_im_status[4], \cceip0_out_im_status.f.wr_pointer [4]);
tran (cceip0_out_im_status[3], \cceip0_out_im_status.r.part0 [3]);
tran (cceip0_out_im_status[3], \cceip0_out_im_status.f.wr_pointer [3]);
tran (cceip0_out_im_status[2], \cceip0_out_im_status.r.part0 [2]);
tran (cceip0_out_im_status[2], \cceip0_out_im_status.f.wr_pointer [2]);
tran (cceip0_out_im_status[1], \cceip0_out_im_status.r.part0 [1]);
tran (cceip0_out_im_status[1], \cceip0_out_im_status.f.wr_pointer [1]);
tran (cceip0_out_im_status[0], \cceip0_out_im_status.r.part0 [0]);
tran (cceip0_out_im_status[0], \cceip0_out_im_status.f.wr_pointer [0]);
tran (cceip1_out_ia_status[16], \cceip1_out_ia_status.r.part0 [16]);
tran (cceip1_out_ia_status[16], \cceip1_out_ia_status.f.code [2]);
tran (cceip1_out_ia_status[15], \cceip1_out_ia_status.r.part0 [15]);
tran (cceip1_out_ia_status[15], \cceip1_out_ia_status.f.code [1]);
tran (cceip1_out_ia_status[14], \cceip1_out_ia_status.r.part0 [14]);
tran (cceip1_out_ia_status[14], \cceip1_out_ia_status.f.code [0]);
tran (cceip1_out_ia_status[13], \cceip1_out_ia_status.r.part0 [13]);
tran (cceip1_out_ia_status[13], \cceip1_out_ia_status.f.datawords [4]);
tran (cceip1_out_ia_status[12], \cceip1_out_ia_status.r.part0 [12]);
tran (cceip1_out_ia_status[12], \cceip1_out_ia_status.f.datawords [3]);
tran (cceip1_out_ia_status[11], \cceip1_out_ia_status.r.part0 [11]);
tran (cceip1_out_ia_status[11], \cceip1_out_ia_status.f.datawords [2]);
tran (cceip1_out_ia_status[10], \cceip1_out_ia_status.r.part0 [10]);
tran (cceip1_out_ia_status[10], \cceip1_out_ia_status.f.datawords [1]);
tran (cceip1_out_ia_status[9], \cceip1_out_ia_status.r.part0 [9]);
tran (cceip1_out_ia_status[9], \cceip1_out_ia_status.f.datawords [0]);
tran (cceip1_out_ia_status[8], \cceip1_out_ia_status.r.part0 [8]);
tran (cceip1_out_ia_status[8], \cceip1_out_ia_status.f.addr [8]);
tran (cceip1_out_ia_status[7], \cceip1_out_ia_status.r.part0 [7]);
tran (cceip1_out_ia_status[7], \cceip1_out_ia_status.f.addr [7]);
tran (cceip1_out_ia_status[6], \cceip1_out_ia_status.r.part0 [6]);
tran (cceip1_out_ia_status[6], \cceip1_out_ia_status.f.addr [6]);
tran (cceip1_out_ia_status[5], \cceip1_out_ia_status.r.part0 [5]);
tran (cceip1_out_ia_status[5], \cceip1_out_ia_status.f.addr [5]);
tran (cceip1_out_ia_status[4], \cceip1_out_ia_status.r.part0 [4]);
tran (cceip1_out_ia_status[4], \cceip1_out_ia_status.f.addr [4]);
tran (cceip1_out_ia_status[3], \cceip1_out_ia_status.r.part0 [3]);
tran (cceip1_out_ia_status[3], \cceip1_out_ia_status.f.addr [3]);
tran (cceip1_out_ia_status[2], \cceip1_out_ia_status.r.part0 [2]);
tran (cceip1_out_ia_status[2], \cceip1_out_ia_status.f.addr [2]);
tran (cceip1_out_ia_status[1], \cceip1_out_ia_status.r.part0 [1]);
tran (cceip1_out_ia_status[1], \cceip1_out_ia_status.f.addr [1]);
tran (cceip1_out_ia_status[0], \cceip1_out_ia_status.r.part0 [0]);
tran (cceip1_out_ia_status[0], \cceip1_out_ia_status.f.addr [0]);
tran (cceip1_out_ia_capability[15], \cceip1_out_ia_capability.r.part0 [15]);
tran (cceip1_out_ia_capability[15], \cceip1_out_ia_capability.f.ack_error );
tran (cceip1_out_ia_capability[14], \cceip1_out_ia_capability.r.part0 [14]);
tran (cceip1_out_ia_capability[14], \cceip1_out_ia_capability.f.sim_tmo );
tran (cceip1_out_ia_capability[13], \cceip1_out_ia_capability.r.part0 [13]);
tran (cceip1_out_ia_capability[13], \cceip1_out_ia_capability.f.reserved_op [3]);
tran (cceip1_out_ia_capability[12], \cceip1_out_ia_capability.r.part0 [12]);
tran (cceip1_out_ia_capability[12], \cceip1_out_ia_capability.f.reserved_op [2]);
tran (cceip1_out_ia_capability[11], \cceip1_out_ia_capability.r.part0 [11]);
tran (cceip1_out_ia_capability[11], \cceip1_out_ia_capability.f.reserved_op [1]);
tran (cceip1_out_ia_capability[10], \cceip1_out_ia_capability.r.part0 [10]);
tran (cceip1_out_ia_capability[10], \cceip1_out_ia_capability.f.reserved_op [0]);
tran (cceip1_out_ia_capability[9], \cceip1_out_ia_capability.r.part0 [9]);
tran (cceip1_out_ia_capability[9], \cceip1_out_ia_capability.f.compare );
tran (cceip1_out_ia_capability[8], \cceip1_out_ia_capability.r.part0 [8]);
tran (cceip1_out_ia_capability[8], \cceip1_out_ia_capability.f.set_init_start );
tran (cceip1_out_ia_capability[7], \cceip1_out_ia_capability.r.part0 [7]);
tran (cceip1_out_ia_capability[7], \cceip1_out_ia_capability.f.initialize_inc );
tran (cceip1_out_ia_capability[6], \cceip1_out_ia_capability.r.part0 [6]);
tran (cceip1_out_ia_capability[6], \cceip1_out_ia_capability.f.initialize );
tran (cceip1_out_ia_capability[5], \cceip1_out_ia_capability.r.part0 [5]);
tran (cceip1_out_ia_capability[5], \cceip1_out_ia_capability.f.reset );
tran (cceip1_out_ia_capability[4], \cceip1_out_ia_capability.r.part0 [4]);
tran (cceip1_out_ia_capability[4], \cceip1_out_ia_capability.f.disabled );
tran (cceip1_out_ia_capability[3], \cceip1_out_ia_capability.r.part0 [3]);
tran (cceip1_out_ia_capability[3], \cceip1_out_ia_capability.f.enable );
tran (cceip1_out_ia_capability[2], \cceip1_out_ia_capability.r.part0 [2]);
tran (cceip1_out_ia_capability[2], \cceip1_out_ia_capability.f.write );
tran (cceip1_out_ia_capability[1], \cceip1_out_ia_capability.r.part0 [1]);
tran (cceip1_out_ia_capability[1], \cceip1_out_ia_capability.f.read );
tran (cceip1_out_ia_capability[0], \cceip1_out_ia_capability.r.part0 [0]);
tran (cceip1_out_ia_capability[0], \cceip1_out_ia_capability.f.nop );
tran (cceip1_out_ia_capability[19], \cceip1_out_ia_capability.r.part0 [19]);
tran (cceip1_out_ia_capability[19], \cceip1_out_ia_capability.f.mem_type [3]);
tran (cceip1_out_ia_capability[18], \cceip1_out_ia_capability.r.part0 [18]);
tran (cceip1_out_ia_capability[18], \cceip1_out_ia_capability.f.mem_type [2]);
tran (cceip1_out_ia_capability[17], \cceip1_out_ia_capability.r.part0 [17]);
tran (cceip1_out_ia_capability[17], \cceip1_out_ia_capability.f.mem_type [1]);
tran (cceip1_out_ia_capability[16], \cceip1_out_ia_capability.r.part0 [16]);
tran (cceip1_out_ia_capability[16], \cceip1_out_ia_capability.f.mem_type [0]);
tran (cceip1_out_ia_rdata[95], \cceip1_out_ia_rdata.r.part2 [31]);
tran (cceip1_out_ia_rdata[95], \cceip1_out_ia_rdata.f.tdata_hi [31]);
tran (cceip1_out_ia_rdata[94], \cceip1_out_ia_rdata.r.part2 [30]);
tran (cceip1_out_ia_rdata[94], \cceip1_out_ia_rdata.f.tdata_hi [30]);
tran (cceip1_out_ia_rdata[93], \cceip1_out_ia_rdata.r.part2 [29]);
tran (cceip1_out_ia_rdata[93], \cceip1_out_ia_rdata.f.tdata_hi [29]);
tran (cceip1_out_ia_rdata[92], \cceip1_out_ia_rdata.r.part2 [28]);
tran (cceip1_out_ia_rdata[92], \cceip1_out_ia_rdata.f.tdata_hi [28]);
tran (cceip1_out_ia_rdata[91], \cceip1_out_ia_rdata.r.part2 [27]);
tran (cceip1_out_ia_rdata[91], \cceip1_out_ia_rdata.f.tdata_hi [27]);
tran (cceip1_out_ia_rdata[90], \cceip1_out_ia_rdata.r.part2 [26]);
tran (cceip1_out_ia_rdata[90], \cceip1_out_ia_rdata.f.tdata_hi [26]);
tran (cceip1_out_ia_rdata[89], \cceip1_out_ia_rdata.r.part2 [25]);
tran (cceip1_out_ia_rdata[89], \cceip1_out_ia_rdata.f.tdata_hi [25]);
tran (cceip1_out_ia_rdata[88], \cceip1_out_ia_rdata.r.part2 [24]);
tran (cceip1_out_ia_rdata[88], \cceip1_out_ia_rdata.f.tdata_hi [24]);
tran (cceip1_out_ia_rdata[87], \cceip1_out_ia_rdata.r.part2 [23]);
tran (cceip1_out_ia_rdata[87], \cceip1_out_ia_rdata.f.tdata_hi [23]);
tran (cceip1_out_ia_rdata[86], \cceip1_out_ia_rdata.r.part2 [22]);
tran (cceip1_out_ia_rdata[86], \cceip1_out_ia_rdata.f.tdata_hi [22]);
tran (cceip1_out_ia_rdata[85], \cceip1_out_ia_rdata.r.part2 [21]);
tran (cceip1_out_ia_rdata[85], \cceip1_out_ia_rdata.f.tdata_hi [21]);
tran (cceip1_out_ia_rdata[84], \cceip1_out_ia_rdata.r.part2 [20]);
tran (cceip1_out_ia_rdata[84], \cceip1_out_ia_rdata.f.tdata_hi [20]);
tran (cceip1_out_ia_rdata[83], \cceip1_out_ia_rdata.r.part2 [19]);
tran (cceip1_out_ia_rdata[83], \cceip1_out_ia_rdata.f.tdata_hi [19]);
tran (cceip1_out_ia_rdata[82], \cceip1_out_ia_rdata.r.part2 [18]);
tran (cceip1_out_ia_rdata[82], \cceip1_out_ia_rdata.f.tdata_hi [18]);
tran (cceip1_out_ia_rdata[81], \cceip1_out_ia_rdata.r.part2 [17]);
tran (cceip1_out_ia_rdata[81], \cceip1_out_ia_rdata.f.tdata_hi [17]);
tran (cceip1_out_ia_rdata[80], \cceip1_out_ia_rdata.r.part2 [16]);
tran (cceip1_out_ia_rdata[80], \cceip1_out_ia_rdata.f.tdata_hi [16]);
tran (cceip1_out_ia_rdata[79], \cceip1_out_ia_rdata.r.part2 [15]);
tran (cceip1_out_ia_rdata[79], \cceip1_out_ia_rdata.f.tdata_hi [15]);
tran (cceip1_out_ia_rdata[78], \cceip1_out_ia_rdata.r.part2 [14]);
tran (cceip1_out_ia_rdata[78], \cceip1_out_ia_rdata.f.tdata_hi [14]);
tran (cceip1_out_ia_rdata[77], \cceip1_out_ia_rdata.r.part2 [13]);
tran (cceip1_out_ia_rdata[77], \cceip1_out_ia_rdata.f.tdata_hi [13]);
tran (cceip1_out_ia_rdata[76], \cceip1_out_ia_rdata.r.part2 [12]);
tran (cceip1_out_ia_rdata[76], \cceip1_out_ia_rdata.f.tdata_hi [12]);
tran (cceip1_out_ia_rdata[75], \cceip1_out_ia_rdata.r.part2 [11]);
tran (cceip1_out_ia_rdata[75], \cceip1_out_ia_rdata.f.tdata_hi [11]);
tran (cceip1_out_ia_rdata[74], \cceip1_out_ia_rdata.r.part2 [10]);
tran (cceip1_out_ia_rdata[74], \cceip1_out_ia_rdata.f.tdata_hi [10]);
tran (cceip1_out_ia_rdata[73], \cceip1_out_ia_rdata.r.part2 [9]);
tran (cceip1_out_ia_rdata[73], \cceip1_out_ia_rdata.f.tdata_hi [9]);
tran (cceip1_out_ia_rdata[72], \cceip1_out_ia_rdata.r.part2 [8]);
tran (cceip1_out_ia_rdata[72], \cceip1_out_ia_rdata.f.tdata_hi [8]);
tran (cceip1_out_ia_rdata[71], \cceip1_out_ia_rdata.r.part2 [7]);
tran (cceip1_out_ia_rdata[71], \cceip1_out_ia_rdata.f.tdata_hi [7]);
tran (cceip1_out_ia_rdata[70], \cceip1_out_ia_rdata.r.part2 [6]);
tran (cceip1_out_ia_rdata[70], \cceip1_out_ia_rdata.f.tdata_hi [6]);
tran (cceip1_out_ia_rdata[69], \cceip1_out_ia_rdata.r.part2 [5]);
tran (cceip1_out_ia_rdata[69], \cceip1_out_ia_rdata.f.tdata_hi [5]);
tran (cceip1_out_ia_rdata[68], \cceip1_out_ia_rdata.r.part2 [4]);
tran (cceip1_out_ia_rdata[68], \cceip1_out_ia_rdata.f.tdata_hi [4]);
tran (cceip1_out_ia_rdata[67], \cceip1_out_ia_rdata.r.part2 [3]);
tran (cceip1_out_ia_rdata[67], \cceip1_out_ia_rdata.f.tdata_hi [3]);
tran (cceip1_out_ia_rdata[66], \cceip1_out_ia_rdata.r.part2 [2]);
tran (cceip1_out_ia_rdata[66], \cceip1_out_ia_rdata.f.tdata_hi [2]);
tran (cceip1_out_ia_rdata[65], \cceip1_out_ia_rdata.r.part2 [1]);
tran (cceip1_out_ia_rdata[65], \cceip1_out_ia_rdata.f.tdata_hi [1]);
tran (cceip1_out_ia_rdata[64], \cceip1_out_ia_rdata.r.part2 [0]);
tran (cceip1_out_ia_rdata[64], \cceip1_out_ia_rdata.f.tdata_hi [0]);
tran (cceip1_out_ia_rdata[63], \cceip1_out_ia_rdata.r.part1 [31]);
tran (cceip1_out_ia_rdata[63], \cceip1_out_ia_rdata.f.tdata_lo [31]);
tran (cceip1_out_ia_rdata[62], \cceip1_out_ia_rdata.r.part1 [30]);
tran (cceip1_out_ia_rdata[62], \cceip1_out_ia_rdata.f.tdata_lo [30]);
tran (cceip1_out_ia_rdata[61], \cceip1_out_ia_rdata.r.part1 [29]);
tran (cceip1_out_ia_rdata[61], \cceip1_out_ia_rdata.f.tdata_lo [29]);
tran (cceip1_out_ia_rdata[60], \cceip1_out_ia_rdata.r.part1 [28]);
tran (cceip1_out_ia_rdata[60], \cceip1_out_ia_rdata.f.tdata_lo [28]);
tran (cceip1_out_ia_rdata[59], \cceip1_out_ia_rdata.r.part1 [27]);
tran (cceip1_out_ia_rdata[59], \cceip1_out_ia_rdata.f.tdata_lo [27]);
tran (cceip1_out_ia_rdata[58], \cceip1_out_ia_rdata.r.part1 [26]);
tran (cceip1_out_ia_rdata[58], \cceip1_out_ia_rdata.f.tdata_lo [26]);
tran (cceip1_out_ia_rdata[57], \cceip1_out_ia_rdata.r.part1 [25]);
tran (cceip1_out_ia_rdata[57], \cceip1_out_ia_rdata.f.tdata_lo [25]);
tran (cceip1_out_ia_rdata[56], \cceip1_out_ia_rdata.r.part1 [24]);
tran (cceip1_out_ia_rdata[56], \cceip1_out_ia_rdata.f.tdata_lo [24]);
tran (cceip1_out_ia_rdata[55], \cceip1_out_ia_rdata.r.part1 [23]);
tran (cceip1_out_ia_rdata[55], \cceip1_out_ia_rdata.f.tdata_lo [23]);
tran (cceip1_out_ia_rdata[54], \cceip1_out_ia_rdata.r.part1 [22]);
tran (cceip1_out_ia_rdata[54], \cceip1_out_ia_rdata.f.tdata_lo [22]);
tran (cceip1_out_ia_rdata[53], \cceip1_out_ia_rdata.r.part1 [21]);
tran (cceip1_out_ia_rdata[53], \cceip1_out_ia_rdata.f.tdata_lo [21]);
tran (cceip1_out_ia_rdata[52], \cceip1_out_ia_rdata.r.part1 [20]);
tran (cceip1_out_ia_rdata[52], \cceip1_out_ia_rdata.f.tdata_lo [20]);
tran (cceip1_out_ia_rdata[51], \cceip1_out_ia_rdata.r.part1 [19]);
tran (cceip1_out_ia_rdata[51], \cceip1_out_ia_rdata.f.tdata_lo [19]);
tran (cceip1_out_ia_rdata[50], \cceip1_out_ia_rdata.r.part1 [18]);
tran (cceip1_out_ia_rdata[50], \cceip1_out_ia_rdata.f.tdata_lo [18]);
tran (cceip1_out_ia_rdata[49], \cceip1_out_ia_rdata.r.part1 [17]);
tran (cceip1_out_ia_rdata[49], \cceip1_out_ia_rdata.f.tdata_lo [17]);
tran (cceip1_out_ia_rdata[48], \cceip1_out_ia_rdata.r.part1 [16]);
tran (cceip1_out_ia_rdata[48], \cceip1_out_ia_rdata.f.tdata_lo [16]);
tran (cceip1_out_ia_rdata[47], \cceip1_out_ia_rdata.r.part1 [15]);
tran (cceip1_out_ia_rdata[47], \cceip1_out_ia_rdata.f.tdata_lo [15]);
tran (cceip1_out_ia_rdata[46], \cceip1_out_ia_rdata.r.part1 [14]);
tran (cceip1_out_ia_rdata[46], \cceip1_out_ia_rdata.f.tdata_lo [14]);
tran (cceip1_out_ia_rdata[45], \cceip1_out_ia_rdata.r.part1 [13]);
tran (cceip1_out_ia_rdata[45], \cceip1_out_ia_rdata.f.tdata_lo [13]);
tran (cceip1_out_ia_rdata[44], \cceip1_out_ia_rdata.r.part1 [12]);
tran (cceip1_out_ia_rdata[44], \cceip1_out_ia_rdata.f.tdata_lo [12]);
tran (cceip1_out_ia_rdata[43], \cceip1_out_ia_rdata.r.part1 [11]);
tran (cceip1_out_ia_rdata[43], \cceip1_out_ia_rdata.f.tdata_lo [11]);
tran (cceip1_out_ia_rdata[42], \cceip1_out_ia_rdata.r.part1 [10]);
tran (cceip1_out_ia_rdata[42], \cceip1_out_ia_rdata.f.tdata_lo [10]);
tran (cceip1_out_ia_rdata[41], \cceip1_out_ia_rdata.r.part1 [9]);
tran (cceip1_out_ia_rdata[41], \cceip1_out_ia_rdata.f.tdata_lo [9]);
tran (cceip1_out_ia_rdata[40], \cceip1_out_ia_rdata.r.part1 [8]);
tran (cceip1_out_ia_rdata[40], \cceip1_out_ia_rdata.f.tdata_lo [8]);
tran (cceip1_out_ia_rdata[39], \cceip1_out_ia_rdata.r.part1 [7]);
tran (cceip1_out_ia_rdata[39], \cceip1_out_ia_rdata.f.tdata_lo [7]);
tran (cceip1_out_ia_rdata[38], \cceip1_out_ia_rdata.r.part1 [6]);
tran (cceip1_out_ia_rdata[38], \cceip1_out_ia_rdata.f.tdata_lo [6]);
tran (cceip1_out_ia_rdata[37], \cceip1_out_ia_rdata.r.part1 [5]);
tran (cceip1_out_ia_rdata[37], \cceip1_out_ia_rdata.f.tdata_lo [5]);
tran (cceip1_out_ia_rdata[36], \cceip1_out_ia_rdata.r.part1 [4]);
tran (cceip1_out_ia_rdata[36], \cceip1_out_ia_rdata.f.tdata_lo [4]);
tran (cceip1_out_ia_rdata[35], \cceip1_out_ia_rdata.r.part1 [3]);
tran (cceip1_out_ia_rdata[35], \cceip1_out_ia_rdata.f.tdata_lo [3]);
tran (cceip1_out_ia_rdata[34], \cceip1_out_ia_rdata.r.part1 [2]);
tran (cceip1_out_ia_rdata[34], \cceip1_out_ia_rdata.f.tdata_lo [2]);
tran (cceip1_out_ia_rdata[33], \cceip1_out_ia_rdata.r.part1 [1]);
tran (cceip1_out_ia_rdata[33], \cceip1_out_ia_rdata.f.tdata_lo [1]);
tran (cceip1_out_ia_rdata[32], \cceip1_out_ia_rdata.r.part1 [0]);
tran (cceip1_out_ia_rdata[32], \cceip1_out_ia_rdata.f.tdata_lo [0]);
tran (cceip1_out_ia_rdata[31], \cceip1_out_ia_rdata.r.part0 [31]);
tran (cceip1_out_ia_rdata[31], \cceip1_out_ia_rdata.f.eob );
tran (cceip1_out_ia_rdata[30], \cceip1_out_ia_rdata.r.part0 [30]);
tran (cceip1_out_ia_rdata[30], \cceip1_out_ia_rdata.f.bytes_vld [7]);
tran (cceip1_out_ia_rdata[29], \cceip1_out_ia_rdata.r.part0 [29]);
tran (cceip1_out_ia_rdata[29], \cceip1_out_ia_rdata.f.bytes_vld [6]);
tran (cceip1_out_ia_rdata[28], \cceip1_out_ia_rdata.r.part0 [28]);
tran (cceip1_out_ia_rdata[28], \cceip1_out_ia_rdata.f.bytes_vld [5]);
tran (cceip1_out_ia_rdata[27], \cceip1_out_ia_rdata.r.part0 [27]);
tran (cceip1_out_ia_rdata[27], \cceip1_out_ia_rdata.f.bytes_vld [4]);
tran (cceip1_out_ia_rdata[26], \cceip1_out_ia_rdata.r.part0 [26]);
tran (cceip1_out_ia_rdata[26], \cceip1_out_ia_rdata.f.bytes_vld [3]);
tran (cceip1_out_ia_rdata[25], \cceip1_out_ia_rdata.r.part0 [25]);
tran (cceip1_out_ia_rdata[25], \cceip1_out_ia_rdata.f.bytes_vld [2]);
tran (cceip1_out_ia_rdata[24], \cceip1_out_ia_rdata.r.part0 [24]);
tran (cceip1_out_ia_rdata[24], \cceip1_out_ia_rdata.f.bytes_vld [1]);
tran (cceip1_out_ia_rdata[23], \cceip1_out_ia_rdata.r.part0 [23]);
tran (cceip1_out_ia_rdata[23], \cceip1_out_ia_rdata.f.bytes_vld [0]);
tran (cceip1_out_ia_rdata[22], \cceip1_out_ia_rdata.r.part0 [22]);
tran (cceip1_out_ia_rdata[22], \cceip1_out_ia_rdata.f.unused1 [7]);
tran (cceip1_out_ia_rdata[21], \cceip1_out_ia_rdata.r.part0 [21]);
tran (cceip1_out_ia_rdata[21], \cceip1_out_ia_rdata.f.unused1 [6]);
tran (cceip1_out_ia_rdata[20], \cceip1_out_ia_rdata.r.part0 [20]);
tran (cceip1_out_ia_rdata[20], \cceip1_out_ia_rdata.f.unused1 [5]);
tran (cceip1_out_ia_rdata[19], \cceip1_out_ia_rdata.r.part0 [19]);
tran (cceip1_out_ia_rdata[19], \cceip1_out_ia_rdata.f.unused1 [4]);
tran (cceip1_out_ia_rdata[18], \cceip1_out_ia_rdata.r.part0 [18]);
tran (cceip1_out_ia_rdata[18], \cceip1_out_ia_rdata.f.unused1 [3]);
tran (cceip1_out_ia_rdata[17], \cceip1_out_ia_rdata.r.part0 [17]);
tran (cceip1_out_ia_rdata[17], \cceip1_out_ia_rdata.f.unused1 [2]);
tran (cceip1_out_ia_rdata[16], \cceip1_out_ia_rdata.r.part0 [16]);
tran (cceip1_out_ia_rdata[16], \cceip1_out_ia_rdata.f.unused1 [1]);
tran (cceip1_out_ia_rdata[15], \cceip1_out_ia_rdata.r.part0 [15]);
tran (cceip1_out_ia_rdata[15], \cceip1_out_ia_rdata.f.unused1 [0]);
tran (cceip1_out_ia_rdata[14], \cceip1_out_ia_rdata.r.part0 [14]);
tran (cceip1_out_ia_rdata[14], \cceip1_out_ia_rdata.f.tid );
tran (cceip1_out_ia_rdata[13], \cceip1_out_ia_rdata.r.part0 [13]);
tran (cceip1_out_ia_rdata[13], \cceip1_out_ia_rdata.f.tuser [7]);
tran (cceip1_out_ia_rdata[12], \cceip1_out_ia_rdata.r.part0 [12]);
tran (cceip1_out_ia_rdata[12], \cceip1_out_ia_rdata.f.tuser [6]);
tran (cceip1_out_ia_rdata[11], \cceip1_out_ia_rdata.r.part0 [11]);
tran (cceip1_out_ia_rdata[11], \cceip1_out_ia_rdata.f.tuser [5]);
tran (cceip1_out_ia_rdata[10], \cceip1_out_ia_rdata.r.part0 [10]);
tran (cceip1_out_ia_rdata[10], \cceip1_out_ia_rdata.f.tuser [4]);
tran (cceip1_out_ia_rdata[9], \cceip1_out_ia_rdata.r.part0 [9]);
tran (cceip1_out_ia_rdata[9], \cceip1_out_ia_rdata.f.tuser [3]);
tran (cceip1_out_ia_rdata[8], \cceip1_out_ia_rdata.r.part0 [8]);
tran (cceip1_out_ia_rdata[8], \cceip1_out_ia_rdata.f.tuser [2]);
tran (cceip1_out_ia_rdata[7], \cceip1_out_ia_rdata.r.part0 [7]);
tran (cceip1_out_ia_rdata[7], \cceip1_out_ia_rdata.f.tuser [1]);
tran (cceip1_out_ia_rdata[6], \cceip1_out_ia_rdata.r.part0 [6]);
tran (cceip1_out_ia_rdata[6], \cceip1_out_ia_rdata.f.tuser [0]);
tran (cceip1_out_ia_rdata[5], \cceip1_out_ia_rdata.r.part0 [5]);
tran (cceip1_out_ia_rdata[5], \cceip1_out_ia_rdata.f.unused0 [5]);
tran (cceip1_out_ia_rdata[4], \cceip1_out_ia_rdata.r.part0 [4]);
tran (cceip1_out_ia_rdata[4], \cceip1_out_ia_rdata.f.unused0 [4]);
tran (cceip1_out_ia_rdata[3], \cceip1_out_ia_rdata.r.part0 [3]);
tran (cceip1_out_ia_rdata[3], \cceip1_out_ia_rdata.f.unused0 [3]);
tran (cceip1_out_ia_rdata[2], \cceip1_out_ia_rdata.r.part0 [2]);
tran (cceip1_out_ia_rdata[2], \cceip1_out_ia_rdata.f.unused0 [2]);
tran (cceip1_out_ia_rdata[1], \cceip1_out_ia_rdata.r.part0 [1]);
tran (cceip1_out_ia_rdata[1], \cceip1_out_ia_rdata.f.unused0 [1]);
tran (cceip1_out_ia_rdata[0], \cceip1_out_ia_rdata.r.part0 [0]);
tran (cceip1_out_ia_rdata[0], \cceip1_out_ia_rdata.f.unused0 [0]);
tran (cceip1_out_im_status[11], \cceip1_out_im_status.r.part0 [11]);
tran (cceip1_out_im_status[11], \cceip1_out_im_status.f.bank_hi );
tran (cceip1_out_im_status[10], \cceip1_out_im_status.r.part0 [10]);
tran (cceip1_out_im_status[10], \cceip1_out_im_status.f.bank_lo );
tran (cceip1_out_im_status[9], \cceip1_out_im_status.r.part0 [9]);
tran (cceip1_out_im_status[9], \cceip1_out_im_status.f.overflow );
tran (cceip1_out_im_status[8], \cceip1_out_im_status.r.part0 [8]);
tran (cceip1_out_im_status[8], \cceip1_out_im_status.f.wr_pointer [8]);
tran (cceip1_out_im_status[7], \cceip1_out_im_status.r.part0 [7]);
tran (cceip1_out_im_status[7], \cceip1_out_im_status.f.wr_pointer [7]);
tran (cceip1_out_im_status[6], \cceip1_out_im_status.r.part0 [6]);
tran (cceip1_out_im_status[6], \cceip1_out_im_status.f.wr_pointer [6]);
tran (cceip1_out_im_status[5], \cceip1_out_im_status.r.part0 [5]);
tran (cceip1_out_im_status[5], \cceip1_out_im_status.f.wr_pointer [5]);
tran (cceip1_out_im_status[4], \cceip1_out_im_status.r.part0 [4]);
tran (cceip1_out_im_status[4], \cceip1_out_im_status.f.wr_pointer [4]);
tran (cceip1_out_im_status[3], \cceip1_out_im_status.r.part0 [3]);
tran (cceip1_out_im_status[3], \cceip1_out_im_status.f.wr_pointer [3]);
tran (cceip1_out_im_status[2], \cceip1_out_im_status.r.part0 [2]);
tran (cceip1_out_im_status[2], \cceip1_out_im_status.f.wr_pointer [2]);
tran (cceip1_out_im_status[1], \cceip1_out_im_status.r.part0 [1]);
tran (cceip1_out_im_status[1], \cceip1_out_im_status.f.wr_pointer [1]);
tran (cceip1_out_im_status[0], \cceip1_out_im_status.r.part0 [0]);
tran (cceip1_out_im_status[0], \cceip1_out_im_status.f.wr_pointer [0]);
tran (cceip2_out_ia_status[16], \cceip2_out_ia_status.r.part0 [16]);
tran (cceip2_out_ia_status[16], \cceip2_out_ia_status.f.code [2]);
tran (cceip2_out_ia_status[15], \cceip2_out_ia_status.r.part0 [15]);
tran (cceip2_out_ia_status[15], \cceip2_out_ia_status.f.code [1]);
tran (cceip2_out_ia_status[14], \cceip2_out_ia_status.r.part0 [14]);
tran (cceip2_out_ia_status[14], \cceip2_out_ia_status.f.code [0]);
tran (cceip2_out_ia_status[13], \cceip2_out_ia_status.r.part0 [13]);
tran (cceip2_out_ia_status[13], \cceip2_out_ia_status.f.datawords [4]);
tran (cceip2_out_ia_status[12], \cceip2_out_ia_status.r.part0 [12]);
tran (cceip2_out_ia_status[12], \cceip2_out_ia_status.f.datawords [3]);
tran (cceip2_out_ia_status[11], \cceip2_out_ia_status.r.part0 [11]);
tran (cceip2_out_ia_status[11], \cceip2_out_ia_status.f.datawords [2]);
tran (cceip2_out_ia_status[10], \cceip2_out_ia_status.r.part0 [10]);
tran (cceip2_out_ia_status[10], \cceip2_out_ia_status.f.datawords [1]);
tran (cceip2_out_ia_status[9], \cceip2_out_ia_status.r.part0 [9]);
tran (cceip2_out_ia_status[9], \cceip2_out_ia_status.f.datawords [0]);
tran (cceip2_out_ia_status[8], \cceip2_out_ia_status.r.part0 [8]);
tran (cceip2_out_ia_status[8], \cceip2_out_ia_status.f.addr [8]);
tran (cceip2_out_ia_status[7], \cceip2_out_ia_status.r.part0 [7]);
tran (cceip2_out_ia_status[7], \cceip2_out_ia_status.f.addr [7]);
tran (cceip2_out_ia_status[6], \cceip2_out_ia_status.r.part0 [6]);
tran (cceip2_out_ia_status[6], \cceip2_out_ia_status.f.addr [6]);
tran (cceip2_out_ia_status[5], \cceip2_out_ia_status.r.part0 [5]);
tran (cceip2_out_ia_status[5], \cceip2_out_ia_status.f.addr [5]);
tran (cceip2_out_ia_status[4], \cceip2_out_ia_status.r.part0 [4]);
tran (cceip2_out_ia_status[4], \cceip2_out_ia_status.f.addr [4]);
tran (cceip2_out_ia_status[3], \cceip2_out_ia_status.r.part0 [3]);
tran (cceip2_out_ia_status[3], \cceip2_out_ia_status.f.addr [3]);
tran (cceip2_out_ia_status[2], \cceip2_out_ia_status.r.part0 [2]);
tran (cceip2_out_ia_status[2], \cceip2_out_ia_status.f.addr [2]);
tran (cceip2_out_ia_status[1], \cceip2_out_ia_status.r.part0 [1]);
tran (cceip2_out_ia_status[1], \cceip2_out_ia_status.f.addr [1]);
tran (cceip2_out_ia_status[0], \cceip2_out_ia_status.r.part0 [0]);
tran (cceip2_out_ia_status[0], \cceip2_out_ia_status.f.addr [0]);
tran (cceip2_out_ia_capability[15], \cceip2_out_ia_capability.r.part0 [15]);
tran (cceip2_out_ia_capability[15], \cceip2_out_ia_capability.f.ack_error );
tran (cceip2_out_ia_capability[14], \cceip2_out_ia_capability.r.part0 [14]);
tran (cceip2_out_ia_capability[14], \cceip2_out_ia_capability.f.sim_tmo );
tran (cceip2_out_ia_capability[13], \cceip2_out_ia_capability.r.part0 [13]);
tran (cceip2_out_ia_capability[13], \cceip2_out_ia_capability.f.reserved_op [3]);
tran (cceip2_out_ia_capability[12], \cceip2_out_ia_capability.r.part0 [12]);
tran (cceip2_out_ia_capability[12], \cceip2_out_ia_capability.f.reserved_op [2]);
tran (cceip2_out_ia_capability[11], \cceip2_out_ia_capability.r.part0 [11]);
tran (cceip2_out_ia_capability[11], \cceip2_out_ia_capability.f.reserved_op [1]);
tran (cceip2_out_ia_capability[10], \cceip2_out_ia_capability.r.part0 [10]);
tran (cceip2_out_ia_capability[10], \cceip2_out_ia_capability.f.reserved_op [0]);
tran (cceip2_out_ia_capability[9], \cceip2_out_ia_capability.r.part0 [9]);
tran (cceip2_out_ia_capability[9], \cceip2_out_ia_capability.f.compare );
tran (cceip2_out_ia_capability[8], \cceip2_out_ia_capability.r.part0 [8]);
tran (cceip2_out_ia_capability[8], \cceip2_out_ia_capability.f.set_init_start );
tran (cceip2_out_ia_capability[7], \cceip2_out_ia_capability.r.part0 [7]);
tran (cceip2_out_ia_capability[7], \cceip2_out_ia_capability.f.initialize_inc );
tran (cceip2_out_ia_capability[6], \cceip2_out_ia_capability.r.part0 [6]);
tran (cceip2_out_ia_capability[6], \cceip2_out_ia_capability.f.initialize );
tran (cceip2_out_ia_capability[5], \cceip2_out_ia_capability.r.part0 [5]);
tran (cceip2_out_ia_capability[5], \cceip2_out_ia_capability.f.reset );
tran (cceip2_out_ia_capability[4], \cceip2_out_ia_capability.r.part0 [4]);
tran (cceip2_out_ia_capability[4], \cceip2_out_ia_capability.f.disabled );
tran (cceip2_out_ia_capability[3], \cceip2_out_ia_capability.r.part0 [3]);
tran (cceip2_out_ia_capability[3], \cceip2_out_ia_capability.f.enable );
tran (cceip2_out_ia_capability[2], \cceip2_out_ia_capability.r.part0 [2]);
tran (cceip2_out_ia_capability[2], \cceip2_out_ia_capability.f.write );
tran (cceip2_out_ia_capability[1], \cceip2_out_ia_capability.r.part0 [1]);
tran (cceip2_out_ia_capability[1], \cceip2_out_ia_capability.f.read );
tran (cceip2_out_ia_capability[0], \cceip2_out_ia_capability.r.part0 [0]);
tran (cceip2_out_ia_capability[0], \cceip2_out_ia_capability.f.nop );
tran (cceip2_out_ia_capability[19], \cceip2_out_ia_capability.r.part0 [19]);
tran (cceip2_out_ia_capability[19], \cceip2_out_ia_capability.f.mem_type [3]);
tran (cceip2_out_ia_capability[18], \cceip2_out_ia_capability.r.part0 [18]);
tran (cceip2_out_ia_capability[18], \cceip2_out_ia_capability.f.mem_type [2]);
tran (cceip2_out_ia_capability[17], \cceip2_out_ia_capability.r.part0 [17]);
tran (cceip2_out_ia_capability[17], \cceip2_out_ia_capability.f.mem_type [1]);
tran (cceip2_out_ia_capability[16], \cceip2_out_ia_capability.r.part0 [16]);
tran (cceip2_out_ia_capability[16], \cceip2_out_ia_capability.f.mem_type [0]);
tran (cceip2_out_ia_rdata[95], \cceip2_out_ia_rdata.r.part2 [31]);
tran (cceip2_out_ia_rdata[95], \cceip2_out_ia_rdata.f.tdata_hi [31]);
tran (cceip2_out_ia_rdata[94], \cceip2_out_ia_rdata.r.part2 [30]);
tran (cceip2_out_ia_rdata[94], \cceip2_out_ia_rdata.f.tdata_hi [30]);
tran (cceip2_out_ia_rdata[93], \cceip2_out_ia_rdata.r.part2 [29]);
tran (cceip2_out_ia_rdata[93], \cceip2_out_ia_rdata.f.tdata_hi [29]);
tran (cceip2_out_ia_rdata[92], \cceip2_out_ia_rdata.r.part2 [28]);
tran (cceip2_out_ia_rdata[92], \cceip2_out_ia_rdata.f.tdata_hi [28]);
tran (cceip2_out_ia_rdata[91], \cceip2_out_ia_rdata.r.part2 [27]);
tran (cceip2_out_ia_rdata[91], \cceip2_out_ia_rdata.f.tdata_hi [27]);
tran (cceip2_out_ia_rdata[90], \cceip2_out_ia_rdata.r.part2 [26]);
tran (cceip2_out_ia_rdata[90], \cceip2_out_ia_rdata.f.tdata_hi [26]);
tran (cceip2_out_ia_rdata[89], \cceip2_out_ia_rdata.r.part2 [25]);
tran (cceip2_out_ia_rdata[89], \cceip2_out_ia_rdata.f.tdata_hi [25]);
tran (cceip2_out_ia_rdata[88], \cceip2_out_ia_rdata.r.part2 [24]);
tran (cceip2_out_ia_rdata[88], \cceip2_out_ia_rdata.f.tdata_hi [24]);
tran (cceip2_out_ia_rdata[87], \cceip2_out_ia_rdata.r.part2 [23]);
tran (cceip2_out_ia_rdata[87], \cceip2_out_ia_rdata.f.tdata_hi [23]);
tran (cceip2_out_ia_rdata[86], \cceip2_out_ia_rdata.r.part2 [22]);
tran (cceip2_out_ia_rdata[86], \cceip2_out_ia_rdata.f.tdata_hi [22]);
tran (cceip2_out_ia_rdata[85], \cceip2_out_ia_rdata.r.part2 [21]);
tran (cceip2_out_ia_rdata[85], \cceip2_out_ia_rdata.f.tdata_hi [21]);
tran (cceip2_out_ia_rdata[84], \cceip2_out_ia_rdata.r.part2 [20]);
tran (cceip2_out_ia_rdata[84], \cceip2_out_ia_rdata.f.tdata_hi [20]);
tran (cceip2_out_ia_rdata[83], \cceip2_out_ia_rdata.r.part2 [19]);
tran (cceip2_out_ia_rdata[83], \cceip2_out_ia_rdata.f.tdata_hi [19]);
tran (cceip2_out_ia_rdata[82], \cceip2_out_ia_rdata.r.part2 [18]);
tran (cceip2_out_ia_rdata[82], \cceip2_out_ia_rdata.f.tdata_hi [18]);
tran (cceip2_out_ia_rdata[81], \cceip2_out_ia_rdata.r.part2 [17]);
tran (cceip2_out_ia_rdata[81], \cceip2_out_ia_rdata.f.tdata_hi [17]);
tran (cceip2_out_ia_rdata[80], \cceip2_out_ia_rdata.r.part2 [16]);
tran (cceip2_out_ia_rdata[80], \cceip2_out_ia_rdata.f.tdata_hi [16]);
tran (cceip2_out_ia_rdata[79], \cceip2_out_ia_rdata.r.part2 [15]);
tran (cceip2_out_ia_rdata[79], \cceip2_out_ia_rdata.f.tdata_hi [15]);
tran (cceip2_out_ia_rdata[78], \cceip2_out_ia_rdata.r.part2 [14]);
tran (cceip2_out_ia_rdata[78], \cceip2_out_ia_rdata.f.tdata_hi [14]);
tran (cceip2_out_ia_rdata[77], \cceip2_out_ia_rdata.r.part2 [13]);
tran (cceip2_out_ia_rdata[77], \cceip2_out_ia_rdata.f.tdata_hi [13]);
tran (cceip2_out_ia_rdata[76], \cceip2_out_ia_rdata.r.part2 [12]);
tran (cceip2_out_ia_rdata[76], \cceip2_out_ia_rdata.f.tdata_hi [12]);
tran (cceip2_out_ia_rdata[75], \cceip2_out_ia_rdata.r.part2 [11]);
tran (cceip2_out_ia_rdata[75], \cceip2_out_ia_rdata.f.tdata_hi [11]);
tran (cceip2_out_ia_rdata[74], \cceip2_out_ia_rdata.r.part2 [10]);
tran (cceip2_out_ia_rdata[74], \cceip2_out_ia_rdata.f.tdata_hi [10]);
tran (cceip2_out_ia_rdata[73], \cceip2_out_ia_rdata.r.part2 [9]);
tran (cceip2_out_ia_rdata[73], \cceip2_out_ia_rdata.f.tdata_hi [9]);
tran (cceip2_out_ia_rdata[72], \cceip2_out_ia_rdata.r.part2 [8]);
tran (cceip2_out_ia_rdata[72], \cceip2_out_ia_rdata.f.tdata_hi [8]);
tran (cceip2_out_ia_rdata[71], \cceip2_out_ia_rdata.r.part2 [7]);
tran (cceip2_out_ia_rdata[71], \cceip2_out_ia_rdata.f.tdata_hi [7]);
tran (cceip2_out_ia_rdata[70], \cceip2_out_ia_rdata.r.part2 [6]);
tran (cceip2_out_ia_rdata[70], \cceip2_out_ia_rdata.f.tdata_hi [6]);
tran (cceip2_out_ia_rdata[69], \cceip2_out_ia_rdata.r.part2 [5]);
tran (cceip2_out_ia_rdata[69], \cceip2_out_ia_rdata.f.tdata_hi [5]);
tran (cceip2_out_ia_rdata[68], \cceip2_out_ia_rdata.r.part2 [4]);
tran (cceip2_out_ia_rdata[68], \cceip2_out_ia_rdata.f.tdata_hi [4]);
tran (cceip2_out_ia_rdata[67], \cceip2_out_ia_rdata.r.part2 [3]);
tran (cceip2_out_ia_rdata[67], \cceip2_out_ia_rdata.f.tdata_hi [3]);
tran (cceip2_out_ia_rdata[66], \cceip2_out_ia_rdata.r.part2 [2]);
tran (cceip2_out_ia_rdata[66], \cceip2_out_ia_rdata.f.tdata_hi [2]);
tran (cceip2_out_ia_rdata[65], \cceip2_out_ia_rdata.r.part2 [1]);
tran (cceip2_out_ia_rdata[65], \cceip2_out_ia_rdata.f.tdata_hi [1]);
tran (cceip2_out_ia_rdata[64], \cceip2_out_ia_rdata.r.part2 [0]);
tran (cceip2_out_ia_rdata[64], \cceip2_out_ia_rdata.f.tdata_hi [0]);
tran (cceip2_out_ia_rdata[63], \cceip2_out_ia_rdata.r.part1 [31]);
tran (cceip2_out_ia_rdata[63], \cceip2_out_ia_rdata.f.tdata_lo [31]);
tran (cceip2_out_ia_rdata[62], \cceip2_out_ia_rdata.r.part1 [30]);
tran (cceip2_out_ia_rdata[62], \cceip2_out_ia_rdata.f.tdata_lo [30]);
tran (cceip2_out_ia_rdata[61], \cceip2_out_ia_rdata.r.part1 [29]);
tran (cceip2_out_ia_rdata[61], \cceip2_out_ia_rdata.f.tdata_lo [29]);
tran (cceip2_out_ia_rdata[60], \cceip2_out_ia_rdata.r.part1 [28]);
tran (cceip2_out_ia_rdata[60], \cceip2_out_ia_rdata.f.tdata_lo [28]);
tran (cceip2_out_ia_rdata[59], \cceip2_out_ia_rdata.r.part1 [27]);
tran (cceip2_out_ia_rdata[59], \cceip2_out_ia_rdata.f.tdata_lo [27]);
tran (cceip2_out_ia_rdata[58], \cceip2_out_ia_rdata.r.part1 [26]);
tran (cceip2_out_ia_rdata[58], \cceip2_out_ia_rdata.f.tdata_lo [26]);
tran (cceip2_out_ia_rdata[57], \cceip2_out_ia_rdata.r.part1 [25]);
tran (cceip2_out_ia_rdata[57], \cceip2_out_ia_rdata.f.tdata_lo [25]);
tran (cceip2_out_ia_rdata[56], \cceip2_out_ia_rdata.r.part1 [24]);
tran (cceip2_out_ia_rdata[56], \cceip2_out_ia_rdata.f.tdata_lo [24]);
tran (cceip2_out_ia_rdata[55], \cceip2_out_ia_rdata.r.part1 [23]);
tran (cceip2_out_ia_rdata[55], \cceip2_out_ia_rdata.f.tdata_lo [23]);
tran (cceip2_out_ia_rdata[54], \cceip2_out_ia_rdata.r.part1 [22]);
tran (cceip2_out_ia_rdata[54], \cceip2_out_ia_rdata.f.tdata_lo [22]);
tran (cceip2_out_ia_rdata[53], \cceip2_out_ia_rdata.r.part1 [21]);
tran (cceip2_out_ia_rdata[53], \cceip2_out_ia_rdata.f.tdata_lo [21]);
tran (cceip2_out_ia_rdata[52], \cceip2_out_ia_rdata.r.part1 [20]);
tran (cceip2_out_ia_rdata[52], \cceip2_out_ia_rdata.f.tdata_lo [20]);
tran (cceip2_out_ia_rdata[51], \cceip2_out_ia_rdata.r.part1 [19]);
tran (cceip2_out_ia_rdata[51], \cceip2_out_ia_rdata.f.tdata_lo [19]);
tran (cceip2_out_ia_rdata[50], \cceip2_out_ia_rdata.r.part1 [18]);
tran (cceip2_out_ia_rdata[50], \cceip2_out_ia_rdata.f.tdata_lo [18]);
tran (cceip2_out_ia_rdata[49], \cceip2_out_ia_rdata.r.part1 [17]);
tran (cceip2_out_ia_rdata[49], \cceip2_out_ia_rdata.f.tdata_lo [17]);
tran (cceip2_out_ia_rdata[48], \cceip2_out_ia_rdata.r.part1 [16]);
tran (cceip2_out_ia_rdata[48], \cceip2_out_ia_rdata.f.tdata_lo [16]);
tran (cceip2_out_ia_rdata[47], \cceip2_out_ia_rdata.r.part1 [15]);
tran (cceip2_out_ia_rdata[47], \cceip2_out_ia_rdata.f.tdata_lo [15]);
tran (cceip2_out_ia_rdata[46], \cceip2_out_ia_rdata.r.part1 [14]);
tran (cceip2_out_ia_rdata[46], \cceip2_out_ia_rdata.f.tdata_lo [14]);
tran (cceip2_out_ia_rdata[45], \cceip2_out_ia_rdata.r.part1 [13]);
tran (cceip2_out_ia_rdata[45], \cceip2_out_ia_rdata.f.tdata_lo [13]);
tran (cceip2_out_ia_rdata[44], \cceip2_out_ia_rdata.r.part1 [12]);
tran (cceip2_out_ia_rdata[44], \cceip2_out_ia_rdata.f.tdata_lo [12]);
tran (cceip2_out_ia_rdata[43], \cceip2_out_ia_rdata.r.part1 [11]);
tran (cceip2_out_ia_rdata[43], \cceip2_out_ia_rdata.f.tdata_lo [11]);
tran (cceip2_out_ia_rdata[42], \cceip2_out_ia_rdata.r.part1 [10]);
tran (cceip2_out_ia_rdata[42], \cceip2_out_ia_rdata.f.tdata_lo [10]);
tran (cceip2_out_ia_rdata[41], \cceip2_out_ia_rdata.r.part1 [9]);
tran (cceip2_out_ia_rdata[41], \cceip2_out_ia_rdata.f.tdata_lo [9]);
tran (cceip2_out_ia_rdata[40], \cceip2_out_ia_rdata.r.part1 [8]);
tran (cceip2_out_ia_rdata[40], \cceip2_out_ia_rdata.f.tdata_lo [8]);
tran (cceip2_out_ia_rdata[39], \cceip2_out_ia_rdata.r.part1 [7]);
tran (cceip2_out_ia_rdata[39], \cceip2_out_ia_rdata.f.tdata_lo [7]);
tran (cceip2_out_ia_rdata[38], \cceip2_out_ia_rdata.r.part1 [6]);
tran (cceip2_out_ia_rdata[38], \cceip2_out_ia_rdata.f.tdata_lo [6]);
tran (cceip2_out_ia_rdata[37], \cceip2_out_ia_rdata.r.part1 [5]);
tran (cceip2_out_ia_rdata[37], \cceip2_out_ia_rdata.f.tdata_lo [5]);
tran (cceip2_out_ia_rdata[36], \cceip2_out_ia_rdata.r.part1 [4]);
tran (cceip2_out_ia_rdata[36], \cceip2_out_ia_rdata.f.tdata_lo [4]);
tran (cceip2_out_ia_rdata[35], \cceip2_out_ia_rdata.r.part1 [3]);
tran (cceip2_out_ia_rdata[35], \cceip2_out_ia_rdata.f.tdata_lo [3]);
tran (cceip2_out_ia_rdata[34], \cceip2_out_ia_rdata.r.part1 [2]);
tran (cceip2_out_ia_rdata[34], \cceip2_out_ia_rdata.f.tdata_lo [2]);
tran (cceip2_out_ia_rdata[33], \cceip2_out_ia_rdata.r.part1 [1]);
tran (cceip2_out_ia_rdata[33], \cceip2_out_ia_rdata.f.tdata_lo [1]);
tran (cceip2_out_ia_rdata[32], \cceip2_out_ia_rdata.r.part1 [0]);
tran (cceip2_out_ia_rdata[32], \cceip2_out_ia_rdata.f.tdata_lo [0]);
tran (cceip2_out_ia_rdata[31], \cceip2_out_ia_rdata.r.part0 [31]);
tran (cceip2_out_ia_rdata[31], \cceip2_out_ia_rdata.f.eob );
tran (cceip2_out_ia_rdata[30], \cceip2_out_ia_rdata.r.part0 [30]);
tran (cceip2_out_ia_rdata[30], \cceip2_out_ia_rdata.f.bytes_vld [7]);
tran (cceip2_out_ia_rdata[29], \cceip2_out_ia_rdata.r.part0 [29]);
tran (cceip2_out_ia_rdata[29], \cceip2_out_ia_rdata.f.bytes_vld [6]);
tran (cceip2_out_ia_rdata[28], \cceip2_out_ia_rdata.r.part0 [28]);
tran (cceip2_out_ia_rdata[28], \cceip2_out_ia_rdata.f.bytes_vld [5]);
tran (cceip2_out_ia_rdata[27], \cceip2_out_ia_rdata.r.part0 [27]);
tran (cceip2_out_ia_rdata[27], \cceip2_out_ia_rdata.f.bytes_vld [4]);
tran (cceip2_out_ia_rdata[26], \cceip2_out_ia_rdata.r.part0 [26]);
tran (cceip2_out_ia_rdata[26], \cceip2_out_ia_rdata.f.bytes_vld [3]);
tran (cceip2_out_ia_rdata[25], \cceip2_out_ia_rdata.r.part0 [25]);
tran (cceip2_out_ia_rdata[25], \cceip2_out_ia_rdata.f.bytes_vld [2]);
tran (cceip2_out_ia_rdata[24], \cceip2_out_ia_rdata.r.part0 [24]);
tran (cceip2_out_ia_rdata[24], \cceip2_out_ia_rdata.f.bytes_vld [1]);
tran (cceip2_out_ia_rdata[23], \cceip2_out_ia_rdata.r.part0 [23]);
tran (cceip2_out_ia_rdata[23], \cceip2_out_ia_rdata.f.bytes_vld [0]);
tran (cceip2_out_ia_rdata[22], \cceip2_out_ia_rdata.r.part0 [22]);
tran (cceip2_out_ia_rdata[22], \cceip2_out_ia_rdata.f.unused1 [7]);
tran (cceip2_out_ia_rdata[21], \cceip2_out_ia_rdata.r.part0 [21]);
tran (cceip2_out_ia_rdata[21], \cceip2_out_ia_rdata.f.unused1 [6]);
tran (cceip2_out_ia_rdata[20], \cceip2_out_ia_rdata.r.part0 [20]);
tran (cceip2_out_ia_rdata[20], \cceip2_out_ia_rdata.f.unused1 [5]);
tran (cceip2_out_ia_rdata[19], \cceip2_out_ia_rdata.r.part0 [19]);
tran (cceip2_out_ia_rdata[19], \cceip2_out_ia_rdata.f.unused1 [4]);
tran (cceip2_out_ia_rdata[18], \cceip2_out_ia_rdata.r.part0 [18]);
tran (cceip2_out_ia_rdata[18], \cceip2_out_ia_rdata.f.unused1 [3]);
tran (cceip2_out_ia_rdata[17], \cceip2_out_ia_rdata.r.part0 [17]);
tran (cceip2_out_ia_rdata[17], \cceip2_out_ia_rdata.f.unused1 [2]);
tran (cceip2_out_ia_rdata[16], \cceip2_out_ia_rdata.r.part0 [16]);
tran (cceip2_out_ia_rdata[16], \cceip2_out_ia_rdata.f.unused1 [1]);
tran (cceip2_out_ia_rdata[15], \cceip2_out_ia_rdata.r.part0 [15]);
tran (cceip2_out_ia_rdata[15], \cceip2_out_ia_rdata.f.unused1 [0]);
tran (cceip2_out_ia_rdata[14], \cceip2_out_ia_rdata.r.part0 [14]);
tran (cceip2_out_ia_rdata[14], \cceip2_out_ia_rdata.f.tid );
tran (cceip2_out_ia_rdata[13], \cceip2_out_ia_rdata.r.part0 [13]);
tran (cceip2_out_ia_rdata[13], \cceip2_out_ia_rdata.f.tuser [7]);
tran (cceip2_out_ia_rdata[12], \cceip2_out_ia_rdata.r.part0 [12]);
tran (cceip2_out_ia_rdata[12], \cceip2_out_ia_rdata.f.tuser [6]);
tran (cceip2_out_ia_rdata[11], \cceip2_out_ia_rdata.r.part0 [11]);
tran (cceip2_out_ia_rdata[11], \cceip2_out_ia_rdata.f.tuser [5]);
tran (cceip2_out_ia_rdata[10], \cceip2_out_ia_rdata.r.part0 [10]);
tran (cceip2_out_ia_rdata[10], \cceip2_out_ia_rdata.f.tuser [4]);
tran (cceip2_out_ia_rdata[9], \cceip2_out_ia_rdata.r.part0 [9]);
tran (cceip2_out_ia_rdata[9], \cceip2_out_ia_rdata.f.tuser [3]);
tran (cceip2_out_ia_rdata[8], \cceip2_out_ia_rdata.r.part0 [8]);
tran (cceip2_out_ia_rdata[8], \cceip2_out_ia_rdata.f.tuser [2]);
tran (cceip2_out_ia_rdata[7], \cceip2_out_ia_rdata.r.part0 [7]);
tran (cceip2_out_ia_rdata[7], \cceip2_out_ia_rdata.f.tuser [1]);
tran (cceip2_out_ia_rdata[6], \cceip2_out_ia_rdata.r.part0 [6]);
tran (cceip2_out_ia_rdata[6], \cceip2_out_ia_rdata.f.tuser [0]);
tran (cceip2_out_ia_rdata[5], \cceip2_out_ia_rdata.r.part0 [5]);
tran (cceip2_out_ia_rdata[5], \cceip2_out_ia_rdata.f.unused0 [5]);
tran (cceip2_out_ia_rdata[4], \cceip2_out_ia_rdata.r.part0 [4]);
tran (cceip2_out_ia_rdata[4], \cceip2_out_ia_rdata.f.unused0 [4]);
tran (cceip2_out_ia_rdata[3], \cceip2_out_ia_rdata.r.part0 [3]);
tran (cceip2_out_ia_rdata[3], \cceip2_out_ia_rdata.f.unused0 [3]);
tran (cceip2_out_ia_rdata[2], \cceip2_out_ia_rdata.r.part0 [2]);
tran (cceip2_out_ia_rdata[2], \cceip2_out_ia_rdata.f.unused0 [2]);
tran (cceip2_out_ia_rdata[1], \cceip2_out_ia_rdata.r.part0 [1]);
tran (cceip2_out_ia_rdata[1], \cceip2_out_ia_rdata.f.unused0 [1]);
tran (cceip2_out_ia_rdata[0], \cceip2_out_ia_rdata.r.part0 [0]);
tran (cceip2_out_ia_rdata[0], \cceip2_out_ia_rdata.f.unused0 [0]);
tran (cceip2_out_im_status[11], \cceip2_out_im_status.r.part0 [11]);
tran (cceip2_out_im_status[11], \cceip2_out_im_status.f.bank_hi );
tran (cceip2_out_im_status[10], \cceip2_out_im_status.r.part0 [10]);
tran (cceip2_out_im_status[10], \cceip2_out_im_status.f.bank_lo );
tran (cceip2_out_im_status[9], \cceip2_out_im_status.r.part0 [9]);
tran (cceip2_out_im_status[9], \cceip2_out_im_status.f.overflow );
tran (cceip2_out_im_status[8], \cceip2_out_im_status.r.part0 [8]);
tran (cceip2_out_im_status[8], \cceip2_out_im_status.f.wr_pointer [8]);
tran (cceip2_out_im_status[7], \cceip2_out_im_status.r.part0 [7]);
tran (cceip2_out_im_status[7], \cceip2_out_im_status.f.wr_pointer [7]);
tran (cceip2_out_im_status[6], \cceip2_out_im_status.r.part0 [6]);
tran (cceip2_out_im_status[6], \cceip2_out_im_status.f.wr_pointer [6]);
tran (cceip2_out_im_status[5], \cceip2_out_im_status.r.part0 [5]);
tran (cceip2_out_im_status[5], \cceip2_out_im_status.f.wr_pointer [5]);
tran (cceip2_out_im_status[4], \cceip2_out_im_status.r.part0 [4]);
tran (cceip2_out_im_status[4], \cceip2_out_im_status.f.wr_pointer [4]);
tran (cceip2_out_im_status[3], \cceip2_out_im_status.r.part0 [3]);
tran (cceip2_out_im_status[3], \cceip2_out_im_status.f.wr_pointer [3]);
tran (cceip2_out_im_status[2], \cceip2_out_im_status.r.part0 [2]);
tran (cceip2_out_im_status[2], \cceip2_out_im_status.f.wr_pointer [2]);
tran (cceip2_out_im_status[1], \cceip2_out_im_status.r.part0 [1]);
tran (cceip2_out_im_status[1], \cceip2_out_im_status.f.wr_pointer [1]);
tran (cceip2_out_im_status[0], \cceip2_out_im_status.r.part0 [0]);
tran (cceip2_out_im_status[0], \cceip2_out_im_status.f.wr_pointer [0]);
tran (cceip3_out_ia_status[16], \cceip3_out_ia_status.r.part0 [16]);
tran (cceip3_out_ia_status[16], \cceip3_out_ia_status.f.code [2]);
tran (cceip3_out_ia_status[15], \cceip3_out_ia_status.r.part0 [15]);
tran (cceip3_out_ia_status[15], \cceip3_out_ia_status.f.code [1]);
tran (cceip3_out_ia_status[14], \cceip3_out_ia_status.r.part0 [14]);
tran (cceip3_out_ia_status[14], \cceip3_out_ia_status.f.code [0]);
tran (cceip3_out_ia_status[13], \cceip3_out_ia_status.r.part0 [13]);
tran (cceip3_out_ia_status[13], \cceip3_out_ia_status.f.datawords [4]);
tran (cceip3_out_ia_status[12], \cceip3_out_ia_status.r.part0 [12]);
tran (cceip3_out_ia_status[12], \cceip3_out_ia_status.f.datawords [3]);
tran (cceip3_out_ia_status[11], \cceip3_out_ia_status.r.part0 [11]);
tran (cceip3_out_ia_status[11], \cceip3_out_ia_status.f.datawords [2]);
tran (cceip3_out_ia_status[10], \cceip3_out_ia_status.r.part0 [10]);
tran (cceip3_out_ia_status[10], \cceip3_out_ia_status.f.datawords [1]);
tran (cceip3_out_ia_status[9], \cceip3_out_ia_status.r.part0 [9]);
tran (cceip3_out_ia_status[9], \cceip3_out_ia_status.f.datawords [0]);
tran (cceip3_out_ia_status[8], \cceip3_out_ia_status.r.part0 [8]);
tran (cceip3_out_ia_status[8], \cceip3_out_ia_status.f.addr [8]);
tran (cceip3_out_ia_status[7], \cceip3_out_ia_status.r.part0 [7]);
tran (cceip3_out_ia_status[7], \cceip3_out_ia_status.f.addr [7]);
tran (cceip3_out_ia_status[6], \cceip3_out_ia_status.r.part0 [6]);
tran (cceip3_out_ia_status[6], \cceip3_out_ia_status.f.addr [6]);
tran (cceip3_out_ia_status[5], \cceip3_out_ia_status.r.part0 [5]);
tran (cceip3_out_ia_status[5], \cceip3_out_ia_status.f.addr [5]);
tran (cceip3_out_ia_status[4], \cceip3_out_ia_status.r.part0 [4]);
tran (cceip3_out_ia_status[4], \cceip3_out_ia_status.f.addr [4]);
tran (cceip3_out_ia_status[3], \cceip3_out_ia_status.r.part0 [3]);
tran (cceip3_out_ia_status[3], \cceip3_out_ia_status.f.addr [3]);
tran (cceip3_out_ia_status[2], \cceip3_out_ia_status.r.part0 [2]);
tran (cceip3_out_ia_status[2], \cceip3_out_ia_status.f.addr [2]);
tran (cceip3_out_ia_status[1], \cceip3_out_ia_status.r.part0 [1]);
tran (cceip3_out_ia_status[1], \cceip3_out_ia_status.f.addr [1]);
tran (cceip3_out_ia_status[0], \cceip3_out_ia_status.r.part0 [0]);
tran (cceip3_out_ia_status[0], \cceip3_out_ia_status.f.addr [0]);
tran (cceip3_out_ia_capability[15], \cceip3_out_ia_capability.r.part0 [15]);
tran (cceip3_out_ia_capability[15], \cceip3_out_ia_capability.f.ack_error );
tran (cceip3_out_ia_capability[14], \cceip3_out_ia_capability.r.part0 [14]);
tran (cceip3_out_ia_capability[14], \cceip3_out_ia_capability.f.sim_tmo );
tran (cceip3_out_ia_capability[13], \cceip3_out_ia_capability.r.part0 [13]);
tran (cceip3_out_ia_capability[13], \cceip3_out_ia_capability.f.reserved_op [3]);
tran (cceip3_out_ia_capability[12], \cceip3_out_ia_capability.r.part0 [12]);
tran (cceip3_out_ia_capability[12], \cceip3_out_ia_capability.f.reserved_op [2]);
tran (cceip3_out_ia_capability[11], \cceip3_out_ia_capability.r.part0 [11]);
tran (cceip3_out_ia_capability[11], \cceip3_out_ia_capability.f.reserved_op [1]);
tran (cceip3_out_ia_capability[10], \cceip3_out_ia_capability.r.part0 [10]);
tran (cceip3_out_ia_capability[10], \cceip3_out_ia_capability.f.reserved_op [0]);
tran (cceip3_out_ia_capability[9], \cceip3_out_ia_capability.r.part0 [9]);
tran (cceip3_out_ia_capability[9], \cceip3_out_ia_capability.f.compare );
tran (cceip3_out_ia_capability[8], \cceip3_out_ia_capability.r.part0 [8]);
tran (cceip3_out_ia_capability[8], \cceip3_out_ia_capability.f.set_init_start );
tran (cceip3_out_ia_capability[7], \cceip3_out_ia_capability.r.part0 [7]);
tran (cceip3_out_ia_capability[7], \cceip3_out_ia_capability.f.initialize_inc );
tran (cceip3_out_ia_capability[6], \cceip3_out_ia_capability.r.part0 [6]);
tran (cceip3_out_ia_capability[6], \cceip3_out_ia_capability.f.initialize );
tran (cceip3_out_ia_capability[5], \cceip3_out_ia_capability.r.part0 [5]);
tran (cceip3_out_ia_capability[5], \cceip3_out_ia_capability.f.reset );
tran (cceip3_out_ia_capability[4], \cceip3_out_ia_capability.r.part0 [4]);
tran (cceip3_out_ia_capability[4], \cceip3_out_ia_capability.f.disabled );
tran (cceip3_out_ia_capability[3], \cceip3_out_ia_capability.r.part0 [3]);
tran (cceip3_out_ia_capability[3], \cceip3_out_ia_capability.f.enable );
tran (cceip3_out_ia_capability[2], \cceip3_out_ia_capability.r.part0 [2]);
tran (cceip3_out_ia_capability[2], \cceip3_out_ia_capability.f.write );
tran (cceip3_out_ia_capability[1], \cceip3_out_ia_capability.r.part0 [1]);
tran (cceip3_out_ia_capability[1], \cceip3_out_ia_capability.f.read );
tran (cceip3_out_ia_capability[0], \cceip3_out_ia_capability.r.part0 [0]);
tran (cceip3_out_ia_capability[0], \cceip3_out_ia_capability.f.nop );
tran (cceip3_out_ia_capability[19], \cceip3_out_ia_capability.r.part0 [19]);
tran (cceip3_out_ia_capability[19], \cceip3_out_ia_capability.f.mem_type [3]);
tran (cceip3_out_ia_capability[18], \cceip3_out_ia_capability.r.part0 [18]);
tran (cceip3_out_ia_capability[18], \cceip3_out_ia_capability.f.mem_type [2]);
tran (cceip3_out_ia_capability[17], \cceip3_out_ia_capability.r.part0 [17]);
tran (cceip3_out_ia_capability[17], \cceip3_out_ia_capability.f.mem_type [1]);
tran (cceip3_out_ia_capability[16], \cceip3_out_ia_capability.r.part0 [16]);
tran (cceip3_out_ia_capability[16], \cceip3_out_ia_capability.f.mem_type [0]);
tran (cceip3_out_ia_rdata[95], \cceip3_out_ia_rdata.r.part2 [31]);
tran (cceip3_out_ia_rdata[95], \cceip3_out_ia_rdata.f.tdata_hi [31]);
tran (cceip3_out_ia_rdata[94], \cceip3_out_ia_rdata.r.part2 [30]);
tran (cceip3_out_ia_rdata[94], \cceip3_out_ia_rdata.f.tdata_hi [30]);
tran (cceip3_out_ia_rdata[93], \cceip3_out_ia_rdata.r.part2 [29]);
tran (cceip3_out_ia_rdata[93], \cceip3_out_ia_rdata.f.tdata_hi [29]);
tran (cceip3_out_ia_rdata[92], \cceip3_out_ia_rdata.r.part2 [28]);
tran (cceip3_out_ia_rdata[92], \cceip3_out_ia_rdata.f.tdata_hi [28]);
tran (cceip3_out_ia_rdata[91], \cceip3_out_ia_rdata.r.part2 [27]);
tran (cceip3_out_ia_rdata[91], \cceip3_out_ia_rdata.f.tdata_hi [27]);
tran (cceip3_out_ia_rdata[90], \cceip3_out_ia_rdata.r.part2 [26]);
tran (cceip3_out_ia_rdata[90], \cceip3_out_ia_rdata.f.tdata_hi [26]);
tran (cceip3_out_ia_rdata[89], \cceip3_out_ia_rdata.r.part2 [25]);
tran (cceip3_out_ia_rdata[89], \cceip3_out_ia_rdata.f.tdata_hi [25]);
tran (cceip3_out_ia_rdata[88], \cceip3_out_ia_rdata.r.part2 [24]);
tran (cceip3_out_ia_rdata[88], \cceip3_out_ia_rdata.f.tdata_hi [24]);
tran (cceip3_out_ia_rdata[87], \cceip3_out_ia_rdata.r.part2 [23]);
tran (cceip3_out_ia_rdata[87], \cceip3_out_ia_rdata.f.tdata_hi [23]);
tran (cceip3_out_ia_rdata[86], \cceip3_out_ia_rdata.r.part2 [22]);
tran (cceip3_out_ia_rdata[86], \cceip3_out_ia_rdata.f.tdata_hi [22]);
tran (cceip3_out_ia_rdata[85], \cceip3_out_ia_rdata.r.part2 [21]);
tran (cceip3_out_ia_rdata[85], \cceip3_out_ia_rdata.f.tdata_hi [21]);
tran (cceip3_out_ia_rdata[84], \cceip3_out_ia_rdata.r.part2 [20]);
tran (cceip3_out_ia_rdata[84], \cceip3_out_ia_rdata.f.tdata_hi [20]);
tran (cceip3_out_ia_rdata[83], \cceip3_out_ia_rdata.r.part2 [19]);
tran (cceip3_out_ia_rdata[83], \cceip3_out_ia_rdata.f.tdata_hi [19]);
tran (cceip3_out_ia_rdata[82], \cceip3_out_ia_rdata.r.part2 [18]);
tran (cceip3_out_ia_rdata[82], \cceip3_out_ia_rdata.f.tdata_hi [18]);
tran (cceip3_out_ia_rdata[81], \cceip3_out_ia_rdata.r.part2 [17]);
tran (cceip3_out_ia_rdata[81], \cceip3_out_ia_rdata.f.tdata_hi [17]);
tran (cceip3_out_ia_rdata[80], \cceip3_out_ia_rdata.r.part2 [16]);
tran (cceip3_out_ia_rdata[80], \cceip3_out_ia_rdata.f.tdata_hi [16]);
tran (cceip3_out_ia_rdata[79], \cceip3_out_ia_rdata.r.part2 [15]);
tran (cceip3_out_ia_rdata[79], \cceip3_out_ia_rdata.f.tdata_hi [15]);
tran (cceip3_out_ia_rdata[78], \cceip3_out_ia_rdata.r.part2 [14]);
tran (cceip3_out_ia_rdata[78], \cceip3_out_ia_rdata.f.tdata_hi [14]);
tran (cceip3_out_ia_rdata[77], \cceip3_out_ia_rdata.r.part2 [13]);
tran (cceip3_out_ia_rdata[77], \cceip3_out_ia_rdata.f.tdata_hi [13]);
tran (cceip3_out_ia_rdata[76], \cceip3_out_ia_rdata.r.part2 [12]);
tran (cceip3_out_ia_rdata[76], \cceip3_out_ia_rdata.f.tdata_hi [12]);
tran (cceip3_out_ia_rdata[75], \cceip3_out_ia_rdata.r.part2 [11]);
tran (cceip3_out_ia_rdata[75], \cceip3_out_ia_rdata.f.tdata_hi [11]);
tran (cceip3_out_ia_rdata[74], \cceip3_out_ia_rdata.r.part2 [10]);
tran (cceip3_out_ia_rdata[74], \cceip3_out_ia_rdata.f.tdata_hi [10]);
tran (cceip3_out_ia_rdata[73], \cceip3_out_ia_rdata.r.part2 [9]);
tran (cceip3_out_ia_rdata[73], \cceip3_out_ia_rdata.f.tdata_hi [9]);
tran (cceip3_out_ia_rdata[72], \cceip3_out_ia_rdata.r.part2 [8]);
tran (cceip3_out_ia_rdata[72], \cceip3_out_ia_rdata.f.tdata_hi [8]);
tran (cceip3_out_ia_rdata[71], \cceip3_out_ia_rdata.r.part2 [7]);
tran (cceip3_out_ia_rdata[71], \cceip3_out_ia_rdata.f.tdata_hi [7]);
tran (cceip3_out_ia_rdata[70], \cceip3_out_ia_rdata.r.part2 [6]);
tran (cceip3_out_ia_rdata[70], \cceip3_out_ia_rdata.f.tdata_hi [6]);
tran (cceip3_out_ia_rdata[69], \cceip3_out_ia_rdata.r.part2 [5]);
tran (cceip3_out_ia_rdata[69], \cceip3_out_ia_rdata.f.tdata_hi [5]);
tran (cceip3_out_ia_rdata[68], \cceip3_out_ia_rdata.r.part2 [4]);
tran (cceip3_out_ia_rdata[68], \cceip3_out_ia_rdata.f.tdata_hi [4]);
tran (cceip3_out_ia_rdata[67], \cceip3_out_ia_rdata.r.part2 [3]);
tran (cceip3_out_ia_rdata[67], \cceip3_out_ia_rdata.f.tdata_hi [3]);
tran (cceip3_out_ia_rdata[66], \cceip3_out_ia_rdata.r.part2 [2]);
tran (cceip3_out_ia_rdata[66], \cceip3_out_ia_rdata.f.tdata_hi [2]);
tran (cceip3_out_ia_rdata[65], \cceip3_out_ia_rdata.r.part2 [1]);
tran (cceip3_out_ia_rdata[65], \cceip3_out_ia_rdata.f.tdata_hi [1]);
tran (cceip3_out_ia_rdata[64], \cceip3_out_ia_rdata.r.part2 [0]);
tran (cceip3_out_ia_rdata[64], \cceip3_out_ia_rdata.f.tdata_hi [0]);
tran (cceip3_out_ia_rdata[63], \cceip3_out_ia_rdata.r.part1 [31]);
tran (cceip3_out_ia_rdata[63], \cceip3_out_ia_rdata.f.tdata_lo [31]);
tran (cceip3_out_ia_rdata[62], \cceip3_out_ia_rdata.r.part1 [30]);
tran (cceip3_out_ia_rdata[62], \cceip3_out_ia_rdata.f.tdata_lo [30]);
tran (cceip3_out_ia_rdata[61], \cceip3_out_ia_rdata.r.part1 [29]);
tran (cceip3_out_ia_rdata[61], \cceip3_out_ia_rdata.f.tdata_lo [29]);
tran (cceip3_out_ia_rdata[60], \cceip3_out_ia_rdata.r.part1 [28]);
tran (cceip3_out_ia_rdata[60], \cceip3_out_ia_rdata.f.tdata_lo [28]);
tran (cceip3_out_ia_rdata[59], \cceip3_out_ia_rdata.r.part1 [27]);
tran (cceip3_out_ia_rdata[59], \cceip3_out_ia_rdata.f.tdata_lo [27]);
tran (cceip3_out_ia_rdata[58], \cceip3_out_ia_rdata.r.part1 [26]);
tran (cceip3_out_ia_rdata[58], \cceip3_out_ia_rdata.f.tdata_lo [26]);
tran (cceip3_out_ia_rdata[57], \cceip3_out_ia_rdata.r.part1 [25]);
tran (cceip3_out_ia_rdata[57], \cceip3_out_ia_rdata.f.tdata_lo [25]);
tran (cceip3_out_ia_rdata[56], \cceip3_out_ia_rdata.r.part1 [24]);
tran (cceip3_out_ia_rdata[56], \cceip3_out_ia_rdata.f.tdata_lo [24]);
tran (cceip3_out_ia_rdata[55], \cceip3_out_ia_rdata.r.part1 [23]);
tran (cceip3_out_ia_rdata[55], \cceip3_out_ia_rdata.f.tdata_lo [23]);
tran (cceip3_out_ia_rdata[54], \cceip3_out_ia_rdata.r.part1 [22]);
tran (cceip3_out_ia_rdata[54], \cceip3_out_ia_rdata.f.tdata_lo [22]);
tran (cceip3_out_ia_rdata[53], \cceip3_out_ia_rdata.r.part1 [21]);
tran (cceip3_out_ia_rdata[53], \cceip3_out_ia_rdata.f.tdata_lo [21]);
tran (cceip3_out_ia_rdata[52], \cceip3_out_ia_rdata.r.part1 [20]);
tran (cceip3_out_ia_rdata[52], \cceip3_out_ia_rdata.f.tdata_lo [20]);
tran (cceip3_out_ia_rdata[51], \cceip3_out_ia_rdata.r.part1 [19]);
tran (cceip3_out_ia_rdata[51], \cceip3_out_ia_rdata.f.tdata_lo [19]);
tran (cceip3_out_ia_rdata[50], \cceip3_out_ia_rdata.r.part1 [18]);
tran (cceip3_out_ia_rdata[50], \cceip3_out_ia_rdata.f.tdata_lo [18]);
tran (cceip3_out_ia_rdata[49], \cceip3_out_ia_rdata.r.part1 [17]);
tran (cceip3_out_ia_rdata[49], \cceip3_out_ia_rdata.f.tdata_lo [17]);
tran (cceip3_out_ia_rdata[48], \cceip3_out_ia_rdata.r.part1 [16]);
tran (cceip3_out_ia_rdata[48], \cceip3_out_ia_rdata.f.tdata_lo [16]);
tran (cceip3_out_ia_rdata[47], \cceip3_out_ia_rdata.r.part1 [15]);
tran (cceip3_out_ia_rdata[47], \cceip3_out_ia_rdata.f.tdata_lo [15]);
tran (cceip3_out_ia_rdata[46], \cceip3_out_ia_rdata.r.part1 [14]);
tran (cceip3_out_ia_rdata[46], \cceip3_out_ia_rdata.f.tdata_lo [14]);
tran (cceip3_out_ia_rdata[45], \cceip3_out_ia_rdata.r.part1 [13]);
tran (cceip3_out_ia_rdata[45], \cceip3_out_ia_rdata.f.tdata_lo [13]);
tran (cceip3_out_ia_rdata[44], \cceip3_out_ia_rdata.r.part1 [12]);
tran (cceip3_out_ia_rdata[44], \cceip3_out_ia_rdata.f.tdata_lo [12]);
tran (cceip3_out_ia_rdata[43], \cceip3_out_ia_rdata.r.part1 [11]);
tran (cceip3_out_ia_rdata[43], \cceip3_out_ia_rdata.f.tdata_lo [11]);
tran (cceip3_out_ia_rdata[42], \cceip3_out_ia_rdata.r.part1 [10]);
tran (cceip3_out_ia_rdata[42], \cceip3_out_ia_rdata.f.tdata_lo [10]);
tran (cceip3_out_ia_rdata[41], \cceip3_out_ia_rdata.r.part1 [9]);
tran (cceip3_out_ia_rdata[41], \cceip3_out_ia_rdata.f.tdata_lo [9]);
tran (cceip3_out_ia_rdata[40], \cceip3_out_ia_rdata.r.part1 [8]);
tran (cceip3_out_ia_rdata[40], \cceip3_out_ia_rdata.f.tdata_lo [8]);
tran (cceip3_out_ia_rdata[39], \cceip3_out_ia_rdata.r.part1 [7]);
tran (cceip3_out_ia_rdata[39], \cceip3_out_ia_rdata.f.tdata_lo [7]);
tran (cceip3_out_ia_rdata[38], \cceip3_out_ia_rdata.r.part1 [6]);
tran (cceip3_out_ia_rdata[38], \cceip3_out_ia_rdata.f.tdata_lo [6]);
tran (cceip3_out_ia_rdata[37], \cceip3_out_ia_rdata.r.part1 [5]);
tran (cceip3_out_ia_rdata[37], \cceip3_out_ia_rdata.f.tdata_lo [5]);
tran (cceip3_out_ia_rdata[36], \cceip3_out_ia_rdata.r.part1 [4]);
tran (cceip3_out_ia_rdata[36], \cceip3_out_ia_rdata.f.tdata_lo [4]);
tran (cceip3_out_ia_rdata[35], \cceip3_out_ia_rdata.r.part1 [3]);
tran (cceip3_out_ia_rdata[35], \cceip3_out_ia_rdata.f.tdata_lo [3]);
tran (cceip3_out_ia_rdata[34], \cceip3_out_ia_rdata.r.part1 [2]);
tran (cceip3_out_ia_rdata[34], \cceip3_out_ia_rdata.f.tdata_lo [2]);
tran (cceip3_out_ia_rdata[33], \cceip3_out_ia_rdata.r.part1 [1]);
tran (cceip3_out_ia_rdata[33], \cceip3_out_ia_rdata.f.tdata_lo [1]);
tran (cceip3_out_ia_rdata[32], \cceip3_out_ia_rdata.r.part1 [0]);
tran (cceip3_out_ia_rdata[32], \cceip3_out_ia_rdata.f.tdata_lo [0]);
tran (cceip3_out_ia_rdata[31], \cceip3_out_ia_rdata.r.part0 [31]);
tran (cceip3_out_ia_rdata[31], \cceip3_out_ia_rdata.f.eob );
tran (cceip3_out_ia_rdata[30], \cceip3_out_ia_rdata.r.part0 [30]);
tran (cceip3_out_ia_rdata[30], \cceip3_out_ia_rdata.f.bytes_vld [7]);
tran (cceip3_out_ia_rdata[29], \cceip3_out_ia_rdata.r.part0 [29]);
tran (cceip3_out_ia_rdata[29], \cceip3_out_ia_rdata.f.bytes_vld [6]);
tran (cceip3_out_ia_rdata[28], \cceip3_out_ia_rdata.r.part0 [28]);
tran (cceip3_out_ia_rdata[28], \cceip3_out_ia_rdata.f.bytes_vld [5]);
tran (cceip3_out_ia_rdata[27], \cceip3_out_ia_rdata.r.part0 [27]);
tran (cceip3_out_ia_rdata[27], \cceip3_out_ia_rdata.f.bytes_vld [4]);
tran (cceip3_out_ia_rdata[26], \cceip3_out_ia_rdata.r.part0 [26]);
tran (cceip3_out_ia_rdata[26], \cceip3_out_ia_rdata.f.bytes_vld [3]);
tran (cceip3_out_ia_rdata[25], \cceip3_out_ia_rdata.r.part0 [25]);
tran (cceip3_out_ia_rdata[25], \cceip3_out_ia_rdata.f.bytes_vld [2]);
tran (cceip3_out_ia_rdata[24], \cceip3_out_ia_rdata.r.part0 [24]);
tran (cceip3_out_ia_rdata[24], \cceip3_out_ia_rdata.f.bytes_vld [1]);
tran (cceip3_out_ia_rdata[23], \cceip3_out_ia_rdata.r.part0 [23]);
tran (cceip3_out_ia_rdata[23], \cceip3_out_ia_rdata.f.bytes_vld [0]);
tran (cceip3_out_ia_rdata[22], \cceip3_out_ia_rdata.r.part0 [22]);
tran (cceip3_out_ia_rdata[22], \cceip3_out_ia_rdata.f.unused1 [7]);
tran (cceip3_out_ia_rdata[21], \cceip3_out_ia_rdata.r.part0 [21]);
tran (cceip3_out_ia_rdata[21], \cceip3_out_ia_rdata.f.unused1 [6]);
tran (cceip3_out_ia_rdata[20], \cceip3_out_ia_rdata.r.part0 [20]);
tran (cceip3_out_ia_rdata[20], \cceip3_out_ia_rdata.f.unused1 [5]);
tran (cceip3_out_ia_rdata[19], \cceip3_out_ia_rdata.r.part0 [19]);
tran (cceip3_out_ia_rdata[19], \cceip3_out_ia_rdata.f.unused1 [4]);
tran (cceip3_out_ia_rdata[18], \cceip3_out_ia_rdata.r.part0 [18]);
tran (cceip3_out_ia_rdata[18], \cceip3_out_ia_rdata.f.unused1 [3]);
tran (cceip3_out_ia_rdata[17], \cceip3_out_ia_rdata.r.part0 [17]);
tran (cceip3_out_ia_rdata[17], \cceip3_out_ia_rdata.f.unused1 [2]);
tran (cceip3_out_ia_rdata[16], \cceip3_out_ia_rdata.r.part0 [16]);
tran (cceip3_out_ia_rdata[16], \cceip3_out_ia_rdata.f.unused1 [1]);
tran (cceip3_out_ia_rdata[15], \cceip3_out_ia_rdata.r.part0 [15]);
tran (cceip3_out_ia_rdata[15], \cceip3_out_ia_rdata.f.unused1 [0]);
tran (cceip3_out_ia_rdata[14], \cceip3_out_ia_rdata.r.part0 [14]);
tran (cceip3_out_ia_rdata[14], \cceip3_out_ia_rdata.f.tid );
tran (cceip3_out_ia_rdata[13], \cceip3_out_ia_rdata.r.part0 [13]);
tran (cceip3_out_ia_rdata[13], \cceip3_out_ia_rdata.f.tuser [7]);
tran (cceip3_out_ia_rdata[12], \cceip3_out_ia_rdata.r.part0 [12]);
tran (cceip3_out_ia_rdata[12], \cceip3_out_ia_rdata.f.tuser [6]);
tran (cceip3_out_ia_rdata[11], \cceip3_out_ia_rdata.r.part0 [11]);
tran (cceip3_out_ia_rdata[11], \cceip3_out_ia_rdata.f.tuser [5]);
tran (cceip3_out_ia_rdata[10], \cceip3_out_ia_rdata.r.part0 [10]);
tran (cceip3_out_ia_rdata[10], \cceip3_out_ia_rdata.f.tuser [4]);
tran (cceip3_out_ia_rdata[9], \cceip3_out_ia_rdata.r.part0 [9]);
tran (cceip3_out_ia_rdata[9], \cceip3_out_ia_rdata.f.tuser [3]);
tran (cceip3_out_ia_rdata[8], \cceip3_out_ia_rdata.r.part0 [8]);
tran (cceip3_out_ia_rdata[8], \cceip3_out_ia_rdata.f.tuser [2]);
tran (cceip3_out_ia_rdata[7], \cceip3_out_ia_rdata.r.part0 [7]);
tran (cceip3_out_ia_rdata[7], \cceip3_out_ia_rdata.f.tuser [1]);
tran (cceip3_out_ia_rdata[6], \cceip3_out_ia_rdata.r.part0 [6]);
tran (cceip3_out_ia_rdata[6], \cceip3_out_ia_rdata.f.tuser [0]);
tran (cceip3_out_ia_rdata[5], \cceip3_out_ia_rdata.r.part0 [5]);
tran (cceip3_out_ia_rdata[5], \cceip3_out_ia_rdata.f.unused0 [5]);
tran (cceip3_out_ia_rdata[4], \cceip3_out_ia_rdata.r.part0 [4]);
tran (cceip3_out_ia_rdata[4], \cceip3_out_ia_rdata.f.unused0 [4]);
tran (cceip3_out_ia_rdata[3], \cceip3_out_ia_rdata.r.part0 [3]);
tran (cceip3_out_ia_rdata[3], \cceip3_out_ia_rdata.f.unused0 [3]);
tran (cceip3_out_ia_rdata[2], \cceip3_out_ia_rdata.r.part0 [2]);
tran (cceip3_out_ia_rdata[2], \cceip3_out_ia_rdata.f.unused0 [2]);
tran (cceip3_out_ia_rdata[1], \cceip3_out_ia_rdata.r.part0 [1]);
tran (cceip3_out_ia_rdata[1], \cceip3_out_ia_rdata.f.unused0 [1]);
tran (cceip3_out_ia_rdata[0], \cceip3_out_ia_rdata.r.part0 [0]);
tran (cceip3_out_ia_rdata[0], \cceip3_out_ia_rdata.f.unused0 [0]);
tran (cceip3_out_im_status[11], \cceip3_out_im_status.r.part0 [11]);
tran (cceip3_out_im_status[11], \cceip3_out_im_status.f.bank_hi );
tran (cceip3_out_im_status[10], \cceip3_out_im_status.r.part0 [10]);
tran (cceip3_out_im_status[10], \cceip3_out_im_status.f.bank_lo );
tran (cceip3_out_im_status[9], \cceip3_out_im_status.r.part0 [9]);
tran (cceip3_out_im_status[9], \cceip3_out_im_status.f.overflow );
tran (cceip3_out_im_status[8], \cceip3_out_im_status.r.part0 [8]);
tran (cceip3_out_im_status[8], \cceip3_out_im_status.f.wr_pointer [8]);
tran (cceip3_out_im_status[7], \cceip3_out_im_status.r.part0 [7]);
tran (cceip3_out_im_status[7], \cceip3_out_im_status.f.wr_pointer [7]);
tran (cceip3_out_im_status[6], \cceip3_out_im_status.r.part0 [6]);
tran (cceip3_out_im_status[6], \cceip3_out_im_status.f.wr_pointer [6]);
tran (cceip3_out_im_status[5], \cceip3_out_im_status.r.part0 [5]);
tran (cceip3_out_im_status[5], \cceip3_out_im_status.f.wr_pointer [5]);
tran (cceip3_out_im_status[4], \cceip3_out_im_status.r.part0 [4]);
tran (cceip3_out_im_status[4], \cceip3_out_im_status.f.wr_pointer [4]);
tran (cceip3_out_im_status[3], \cceip3_out_im_status.r.part0 [3]);
tran (cceip3_out_im_status[3], \cceip3_out_im_status.f.wr_pointer [3]);
tran (cceip3_out_im_status[2], \cceip3_out_im_status.r.part0 [2]);
tran (cceip3_out_im_status[2], \cceip3_out_im_status.f.wr_pointer [2]);
tran (cceip3_out_im_status[1], \cceip3_out_im_status.r.part0 [1]);
tran (cceip3_out_im_status[1], \cceip3_out_im_status.f.wr_pointer [1]);
tran (cceip3_out_im_status[0], \cceip3_out_im_status.r.part0 [0]);
tran (cceip3_out_im_status[0], \cceip3_out_im_status.f.wr_pointer [0]);
tran (cddip0_out_ia_status[16], \cddip0_out_ia_status.r.part0 [16]);
tran (cddip0_out_ia_status[16], \cddip0_out_ia_status.f.code [2]);
tran (cddip0_out_ia_status[15], \cddip0_out_ia_status.r.part0 [15]);
tran (cddip0_out_ia_status[15], \cddip0_out_ia_status.f.code [1]);
tran (cddip0_out_ia_status[14], \cddip0_out_ia_status.r.part0 [14]);
tran (cddip0_out_ia_status[14], \cddip0_out_ia_status.f.code [0]);
tran (cddip0_out_ia_status[13], \cddip0_out_ia_status.r.part0 [13]);
tran (cddip0_out_ia_status[13], \cddip0_out_ia_status.f.datawords [4]);
tran (cddip0_out_ia_status[12], \cddip0_out_ia_status.r.part0 [12]);
tran (cddip0_out_ia_status[12], \cddip0_out_ia_status.f.datawords [3]);
tran (cddip0_out_ia_status[11], \cddip0_out_ia_status.r.part0 [11]);
tran (cddip0_out_ia_status[11], \cddip0_out_ia_status.f.datawords [2]);
tran (cddip0_out_ia_status[10], \cddip0_out_ia_status.r.part0 [10]);
tran (cddip0_out_ia_status[10], \cddip0_out_ia_status.f.datawords [1]);
tran (cddip0_out_ia_status[9], \cddip0_out_ia_status.r.part0 [9]);
tran (cddip0_out_ia_status[9], \cddip0_out_ia_status.f.datawords [0]);
tran (cddip0_out_ia_status[8], \cddip0_out_ia_status.r.part0 [8]);
tran (cddip0_out_ia_status[8], \cddip0_out_ia_status.f.addr [8]);
tran (cddip0_out_ia_status[7], \cddip0_out_ia_status.r.part0 [7]);
tran (cddip0_out_ia_status[7], \cddip0_out_ia_status.f.addr [7]);
tran (cddip0_out_ia_status[6], \cddip0_out_ia_status.r.part0 [6]);
tran (cddip0_out_ia_status[6], \cddip0_out_ia_status.f.addr [6]);
tran (cddip0_out_ia_status[5], \cddip0_out_ia_status.r.part0 [5]);
tran (cddip0_out_ia_status[5], \cddip0_out_ia_status.f.addr [5]);
tran (cddip0_out_ia_status[4], \cddip0_out_ia_status.r.part0 [4]);
tran (cddip0_out_ia_status[4], \cddip0_out_ia_status.f.addr [4]);
tran (cddip0_out_ia_status[3], \cddip0_out_ia_status.r.part0 [3]);
tran (cddip0_out_ia_status[3], \cddip0_out_ia_status.f.addr [3]);
tran (cddip0_out_ia_status[2], \cddip0_out_ia_status.r.part0 [2]);
tran (cddip0_out_ia_status[2], \cddip0_out_ia_status.f.addr [2]);
tran (cddip0_out_ia_status[1], \cddip0_out_ia_status.r.part0 [1]);
tran (cddip0_out_ia_status[1], \cddip0_out_ia_status.f.addr [1]);
tran (cddip0_out_ia_status[0], \cddip0_out_ia_status.r.part0 [0]);
tran (cddip0_out_ia_status[0], \cddip0_out_ia_status.f.addr [0]);
tran (cddip0_out_ia_capability[15], \cddip0_out_ia_capability.r.part0 [15]);
tran (cddip0_out_ia_capability[15], \cddip0_out_ia_capability.f.ack_error );
tran (cddip0_out_ia_capability[14], \cddip0_out_ia_capability.r.part0 [14]);
tran (cddip0_out_ia_capability[14], \cddip0_out_ia_capability.f.sim_tmo );
tran (cddip0_out_ia_capability[13], \cddip0_out_ia_capability.r.part0 [13]);
tran (cddip0_out_ia_capability[13], \cddip0_out_ia_capability.f.reserved_op [3]);
tran (cddip0_out_ia_capability[12], \cddip0_out_ia_capability.r.part0 [12]);
tran (cddip0_out_ia_capability[12], \cddip0_out_ia_capability.f.reserved_op [2]);
tran (cddip0_out_ia_capability[11], \cddip0_out_ia_capability.r.part0 [11]);
tran (cddip0_out_ia_capability[11], \cddip0_out_ia_capability.f.reserved_op [1]);
tran (cddip0_out_ia_capability[10], \cddip0_out_ia_capability.r.part0 [10]);
tran (cddip0_out_ia_capability[10], \cddip0_out_ia_capability.f.reserved_op [0]);
tran (cddip0_out_ia_capability[9], \cddip0_out_ia_capability.r.part0 [9]);
tran (cddip0_out_ia_capability[9], \cddip0_out_ia_capability.f.compare );
tran (cddip0_out_ia_capability[8], \cddip0_out_ia_capability.r.part0 [8]);
tran (cddip0_out_ia_capability[8], \cddip0_out_ia_capability.f.set_init_start );
tran (cddip0_out_ia_capability[7], \cddip0_out_ia_capability.r.part0 [7]);
tran (cddip0_out_ia_capability[7], \cddip0_out_ia_capability.f.initialize_inc );
tran (cddip0_out_ia_capability[6], \cddip0_out_ia_capability.r.part0 [6]);
tran (cddip0_out_ia_capability[6], \cddip0_out_ia_capability.f.initialize );
tran (cddip0_out_ia_capability[5], \cddip0_out_ia_capability.r.part0 [5]);
tran (cddip0_out_ia_capability[5], \cddip0_out_ia_capability.f.reset );
tran (cddip0_out_ia_capability[4], \cddip0_out_ia_capability.r.part0 [4]);
tran (cddip0_out_ia_capability[4], \cddip0_out_ia_capability.f.disabled );
tran (cddip0_out_ia_capability[3], \cddip0_out_ia_capability.r.part0 [3]);
tran (cddip0_out_ia_capability[3], \cddip0_out_ia_capability.f.enable );
tran (cddip0_out_ia_capability[2], \cddip0_out_ia_capability.r.part0 [2]);
tran (cddip0_out_ia_capability[2], \cddip0_out_ia_capability.f.write );
tran (cddip0_out_ia_capability[1], \cddip0_out_ia_capability.r.part0 [1]);
tran (cddip0_out_ia_capability[1], \cddip0_out_ia_capability.f.read );
tran (cddip0_out_ia_capability[0], \cddip0_out_ia_capability.r.part0 [0]);
tran (cddip0_out_ia_capability[0], \cddip0_out_ia_capability.f.nop );
tran (cddip0_out_ia_capability[19], \cddip0_out_ia_capability.r.part0 [19]);
tran (cddip0_out_ia_capability[19], \cddip0_out_ia_capability.f.mem_type [3]);
tran (cddip0_out_ia_capability[18], \cddip0_out_ia_capability.r.part0 [18]);
tran (cddip0_out_ia_capability[18], \cddip0_out_ia_capability.f.mem_type [2]);
tran (cddip0_out_ia_capability[17], \cddip0_out_ia_capability.r.part0 [17]);
tran (cddip0_out_ia_capability[17], \cddip0_out_ia_capability.f.mem_type [1]);
tran (cddip0_out_ia_capability[16], \cddip0_out_ia_capability.r.part0 [16]);
tran (cddip0_out_ia_capability[16], \cddip0_out_ia_capability.f.mem_type [0]);
tran (cddip0_out_ia_rdata[95], \cddip0_out_ia_rdata.r.part2 [31]);
tran (cddip0_out_ia_rdata[95], \cddip0_out_ia_rdata.f.tdata_hi [31]);
tran (cddip0_out_ia_rdata[94], \cddip0_out_ia_rdata.r.part2 [30]);
tran (cddip0_out_ia_rdata[94], \cddip0_out_ia_rdata.f.tdata_hi [30]);
tran (cddip0_out_ia_rdata[93], \cddip0_out_ia_rdata.r.part2 [29]);
tran (cddip0_out_ia_rdata[93], \cddip0_out_ia_rdata.f.tdata_hi [29]);
tran (cddip0_out_ia_rdata[92], \cddip0_out_ia_rdata.r.part2 [28]);
tran (cddip0_out_ia_rdata[92], \cddip0_out_ia_rdata.f.tdata_hi [28]);
tran (cddip0_out_ia_rdata[91], \cddip0_out_ia_rdata.r.part2 [27]);
tran (cddip0_out_ia_rdata[91], \cddip0_out_ia_rdata.f.tdata_hi [27]);
tran (cddip0_out_ia_rdata[90], \cddip0_out_ia_rdata.r.part2 [26]);
tran (cddip0_out_ia_rdata[90], \cddip0_out_ia_rdata.f.tdata_hi [26]);
tran (cddip0_out_ia_rdata[89], \cddip0_out_ia_rdata.r.part2 [25]);
tran (cddip0_out_ia_rdata[89], \cddip0_out_ia_rdata.f.tdata_hi [25]);
tran (cddip0_out_ia_rdata[88], \cddip0_out_ia_rdata.r.part2 [24]);
tran (cddip0_out_ia_rdata[88], \cddip0_out_ia_rdata.f.tdata_hi [24]);
tran (cddip0_out_ia_rdata[87], \cddip0_out_ia_rdata.r.part2 [23]);
tran (cddip0_out_ia_rdata[87], \cddip0_out_ia_rdata.f.tdata_hi [23]);
tran (cddip0_out_ia_rdata[86], \cddip0_out_ia_rdata.r.part2 [22]);
tran (cddip0_out_ia_rdata[86], \cddip0_out_ia_rdata.f.tdata_hi [22]);
tran (cddip0_out_ia_rdata[85], \cddip0_out_ia_rdata.r.part2 [21]);
tran (cddip0_out_ia_rdata[85], \cddip0_out_ia_rdata.f.tdata_hi [21]);
tran (cddip0_out_ia_rdata[84], \cddip0_out_ia_rdata.r.part2 [20]);
tran (cddip0_out_ia_rdata[84], \cddip0_out_ia_rdata.f.tdata_hi [20]);
tran (cddip0_out_ia_rdata[83], \cddip0_out_ia_rdata.r.part2 [19]);
tran (cddip0_out_ia_rdata[83], \cddip0_out_ia_rdata.f.tdata_hi [19]);
tran (cddip0_out_ia_rdata[82], \cddip0_out_ia_rdata.r.part2 [18]);
tran (cddip0_out_ia_rdata[82], \cddip0_out_ia_rdata.f.tdata_hi [18]);
tran (cddip0_out_ia_rdata[81], \cddip0_out_ia_rdata.r.part2 [17]);
tran (cddip0_out_ia_rdata[81], \cddip0_out_ia_rdata.f.tdata_hi [17]);
tran (cddip0_out_ia_rdata[80], \cddip0_out_ia_rdata.r.part2 [16]);
tran (cddip0_out_ia_rdata[80], \cddip0_out_ia_rdata.f.tdata_hi [16]);
tran (cddip0_out_ia_rdata[79], \cddip0_out_ia_rdata.r.part2 [15]);
tran (cddip0_out_ia_rdata[79], \cddip0_out_ia_rdata.f.tdata_hi [15]);
tran (cddip0_out_ia_rdata[78], \cddip0_out_ia_rdata.r.part2 [14]);
tran (cddip0_out_ia_rdata[78], \cddip0_out_ia_rdata.f.tdata_hi [14]);
tran (cddip0_out_ia_rdata[77], \cddip0_out_ia_rdata.r.part2 [13]);
tran (cddip0_out_ia_rdata[77], \cddip0_out_ia_rdata.f.tdata_hi [13]);
tran (cddip0_out_ia_rdata[76], \cddip0_out_ia_rdata.r.part2 [12]);
tran (cddip0_out_ia_rdata[76], \cddip0_out_ia_rdata.f.tdata_hi [12]);
tran (cddip0_out_ia_rdata[75], \cddip0_out_ia_rdata.r.part2 [11]);
tran (cddip0_out_ia_rdata[75], \cddip0_out_ia_rdata.f.tdata_hi [11]);
tran (cddip0_out_ia_rdata[74], \cddip0_out_ia_rdata.r.part2 [10]);
tran (cddip0_out_ia_rdata[74], \cddip0_out_ia_rdata.f.tdata_hi [10]);
tran (cddip0_out_ia_rdata[73], \cddip0_out_ia_rdata.r.part2 [9]);
tran (cddip0_out_ia_rdata[73], \cddip0_out_ia_rdata.f.tdata_hi [9]);
tran (cddip0_out_ia_rdata[72], \cddip0_out_ia_rdata.r.part2 [8]);
tran (cddip0_out_ia_rdata[72], \cddip0_out_ia_rdata.f.tdata_hi [8]);
tran (cddip0_out_ia_rdata[71], \cddip0_out_ia_rdata.r.part2 [7]);
tran (cddip0_out_ia_rdata[71], \cddip0_out_ia_rdata.f.tdata_hi [7]);
tran (cddip0_out_ia_rdata[70], \cddip0_out_ia_rdata.r.part2 [6]);
tran (cddip0_out_ia_rdata[70], \cddip0_out_ia_rdata.f.tdata_hi [6]);
tran (cddip0_out_ia_rdata[69], \cddip0_out_ia_rdata.r.part2 [5]);
tran (cddip0_out_ia_rdata[69], \cddip0_out_ia_rdata.f.tdata_hi [5]);
tran (cddip0_out_ia_rdata[68], \cddip0_out_ia_rdata.r.part2 [4]);
tran (cddip0_out_ia_rdata[68], \cddip0_out_ia_rdata.f.tdata_hi [4]);
tran (cddip0_out_ia_rdata[67], \cddip0_out_ia_rdata.r.part2 [3]);
tran (cddip0_out_ia_rdata[67], \cddip0_out_ia_rdata.f.tdata_hi [3]);
tran (cddip0_out_ia_rdata[66], \cddip0_out_ia_rdata.r.part2 [2]);
tran (cddip0_out_ia_rdata[66], \cddip0_out_ia_rdata.f.tdata_hi [2]);
tran (cddip0_out_ia_rdata[65], \cddip0_out_ia_rdata.r.part2 [1]);
tran (cddip0_out_ia_rdata[65], \cddip0_out_ia_rdata.f.tdata_hi [1]);
tran (cddip0_out_ia_rdata[64], \cddip0_out_ia_rdata.r.part2 [0]);
tran (cddip0_out_ia_rdata[64], \cddip0_out_ia_rdata.f.tdata_hi [0]);
tran (cddip0_out_ia_rdata[63], \cddip0_out_ia_rdata.r.part1 [31]);
tran (cddip0_out_ia_rdata[63], \cddip0_out_ia_rdata.f.tdata_lo [31]);
tran (cddip0_out_ia_rdata[62], \cddip0_out_ia_rdata.r.part1 [30]);
tran (cddip0_out_ia_rdata[62], \cddip0_out_ia_rdata.f.tdata_lo [30]);
tran (cddip0_out_ia_rdata[61], \cddip0_out_ia_rdata.r.part1 [29]);
tran (cddip0_out_ia_rdata[61], \cddip0_out_ia_rdata.f.tdata_lo [29]);
tran (cddip0_out_ia_rdata[60], \cddip0_out_ia_rdata.r.part1 [28]);
tran (cddip0_out_ia_rdata[60], \cddip0_out_ia_rdata.f.tdata_lo [28]);
tran (cddip0_out_ia_rdata[59], \cddip0_out_ia_rdata.r.part1 [27]);
tran (cddip0_out_ia_rdata[59], \cddip0_out_ia_rdata.f.tdata_lo [27]);
tran (cddip0_out_ia_rdata[58], \cddip0_out_ia_rdata.r.part1 [26]);
tran (cddip0_out_ia_rdata[58], \cddip0_out_ia_rdata.f.tdata_lo [26]);
tran (cddip0_out_ia_rdata[57], \cddip0_out_ia_rdata.r.part1 [25]);
tran (cddip0_out_ia_rdata[57], \cddip0_out_ia_rdata.f.tdata_lo [25]);
tran (cddip0_out_ia_rdata[56], \cddip0_out_ia_rdata.r.part1 [24]);
tran (cddip0_out_ia_rdata[56], \cddip0_out_ia_rdata.f.tdata_lo [24]);
tran (cddip0_out_ia_rdata[55], \cddip0_out_ia_rdata.r.part1 [23]);
tran (cddip0_out_ia_rdata[55], \cddip0_out_ia_rdata.f.tdata_lo [23]);
tran (cddip0_out_ia_rdata[54], \cddip0_out_ia_rdata.r.part1 [22]);
tran (cddip0_out_ia_rdata[54], \cddip0_out_ia_rdata.f.tdata_lo [22]);
tran (cddip0_out_ia_rdata[53], \cddip0_out_ia_rdata.r.part1 [21]);
tran (cddip0_out_ia_rdata[53], \cddip0_out_ia_rdata.f.tdata_lo [21]);
tran (cddip0_out_ia_rdata[52], \cddip0_out_ia_rdata.r.part1 [20]);
tran (cddip0_out_ia_rdata[52], \cddip0_out_ia_rdata.f.tdata_lo [20]);
tran (cddip0_out_ia_rdata[51], \cddip0_out_ia_rdata.r.part1 [19]);
tran (cddip0_out_ia_rdata[51], \cddip0_out_ia_rdata.f.tdata_lo [19]);
tran (cddip0_out_ia_rdata[50], \cddip0_out_ia_rdata.r.part1 [18]);
tran (cddip0_out_ia_rdata[50], \cddip0_out_ia_rdata.f.tdata_lo [18]);
tran (cddip0_out_ia_rdata[49], \cddip0_out_ia_rdata.r.part1 [17]);
tran (cddip0_out_ia_rdata[49], \cddip0_out_ia_rdata.f.tdata_lo [17]);
tran (cddip0_out_ia_rdata[48], \cddip0_out_ia_rdata.r.part1 [16]);
tran (cddip0_out_ia_rdata[48], \cddip0_out_ia_rdata.f.tdata_lo [16]);
tran (cddip0_out_ia_rdata[47], \cddip0_out_ia_rdata.r.part1 [15]);
tran (cddip0_out_ia_rdata[47], \cddip0_out_ia_rdata.f.tdata_lo [15]);
tran (cddip0_out_ia_rdata[46], \cddip0_out_ia_rdata.r.part1 [14]);
tran (cddip0_out_ia_rdata[46], \cddip0_out_ia_rdata.f.tdata_lo [14]);
tran (cddip0_out_ia_rdata[45], \cddip0_out_ia_rdata.r.part1 [13]);
tran (cddip0_out_ia_rdata[45], \cddip0_out_ia_rdata.f.tdata_lo [13]);
tran (cddip0_out_ia_rdata[44], \cddip0_out_ia_rdata.r.part1 [12]);
tran (cddip0_out_ia_rdata[44], \cddip0_out_ia_rdata.f.tdata_lo [12]);
tran (cddip0_out_ia_rdata[43], \cddip0_out_ia_rdata.r.part1 [11]);
tran (cddip0_out_ia_rdata[43], \cddip0_out_ia_rdata.f.tdata_lo [11]);
tran (cddip0_out_ia_rdata[42], \cddip0_out_ia_rdata.r.part1 [10]);
tran (cddip0_out_ia_rdata[42], \cddip0_out_ia_rdata.f.tdata_lo [10]);
tran (cddip0_out_ia_rdata[41], \cddip0_out_ia_rdata.r.part1 [9]);
tran (cddip0_out_ia_rdata[41], \cddip0_out_ia_rdata.f.tdata_lo [9]);
tran (cddip0_out_ia_rdata[40], \cddip0_out_ia_rdata.r.part1 [8]);
tran (cddip0_out_ia_rdata[40], \cddip0_out_ia_rdata.f.tdata_lo [8]);
tran (cddip0_out_ia_rdata[39], \cddip0_out_ia_rdata.r.part1 [7]);
tran (cddip0_out_ia_rdata[39], \cddip0_out_ia_rdata.f.tdata_lo [7]);
tran (cddip0_out_ia_rdata[38], \cddip0_out_ia_rdata.r.part1 [6]);
tran (cddip0_out_ia_rdata[38], \cddip0_out_ia_rdata.f.tdata_lo [6]);
tran (cddip0_out_ia_rdata[37], \cddip0_out_ia_rdata.r.part1 [5]);
tran (cddip0_out_ia_rdata[37], \cddip0_out_ia_rdata.f.tdata_lo [5]);
tran (cddip0_out_ia_rdata[36], \cddip0_out_ia_rdata.r.part1 [4]);
tran (cddip0_out_ia_rdata[36], \cddip0_out_ia_rdata.f.tdata_lo [4]);
tran (cddip0_out_ia_rdata[35], \cddip0_out_ia_rdata.r.part1 [3]);
tran (cddip0_out_ia_rdata[35], \cddip0_out_ia_rdata.f.tdata_lo [3]);
tran (cddip0_out_ia_rdata[34], \cddip0_out_ia_rdata.r.part1 [2]);
tran (cddip0_out_ia_rdata[34], \cddip0_out_ia_rdata.f.tdata_lo [2]);
tran (cddip0_out_ia_rdata[33], \cddip0_out_ia_rdata.r.part1 [1]);
tran (cddip0_out_ia_rdata[33], \cddip0_out_ia_rdata.f.tdata_lo [1]);
tran (cddip0_out_ia_rdata[32], \cddip0_out_ia_rdata.r.part1 [0]);
tran (cddip0_out_ia_rdata[32], \cddip0_out_ia_rdata.f.tdata_lo [0]);
tran (cddip0_out_ia_rdata[31], \cddip0_out_ia_rdata.r.part0 [31]);
tran (cddip0_out_ia_rdata[31], \cddip0_out_ia_rdata.f.eob );
tran (cddip0_out_ia_rdata[30], \cddip0_out_ia_rdata.r.part0 [30]);
tran (cddip0_out_ia_rdata[30], \cddip0_out_ia_rdata.f.bytes_vld [7]);
tran (cddip0_out_ia_rdata[29], \cddip0_out_ia_rdata.r.part0 [29]);
tran (cddip0_out_ia_rdata[29], \cddip0_out_ia_rdata.f.bytes_vld [6]);
tran (cddip0_out_ia_rdata[28], \cddip0_out_ia_rdata.r.part0 [28]);
tran (cddip0_out_ia_rdata[28], \cddip0_out_ia_rdata.f.bytes_vld [5]);
tran (cddip0_out_ia_rdata[27], \cddip0_out_ia_rdata.r.part0 [27]);
tran (cddip0_out_ia_rdata[27], \cddip0_out_ia_rdata.f.bytes_vld [4]);
tran (cddip0_out_ia_rdata[26], \cddip0_out_ia_rdata.r.part0 [26]);
tran (cddip0_out_ia_rdata[26], \cddip0_out_ia_rdata.f.bytes_vld [3]);
tran (cddip0_out_ia_rdata[25], \cddip0_out_ia_rdata.r.part0 [25]);
tran (cddip0_out_ia_rdata[25], \cddip0_out_ia_rdata.f.bytes_vld [2]);
tran (cddip0_out_ia_rdata[24], \cddip0_out_ia_rdata.r.part0 [24]);
tran (cddip0_out_ia_rdata[24], \cddip0_out_ia_rdata.f.bytes_vld [1]);
tran (cddip0_out_ia_rdata[23], \cddip0_out_ia_rdata.r.part0 [23]);
tran (cddip0_out_ia_rdata[23], \cddip0_out_ia_rdata.f.bytes_vld [0]);
tran (cddip0_out_ia_rdata[22], \cddip0_out_ia_rdata.r.part0 [22]);
tran (cddip0_out_ia_rdata[22], \cddip0_out_ia_rdata.f.unused1 [7]);
tran (cddip0_out_ia_rdata[21], \cddip0_out_ia_rdata.r.part0 [21]);
tran (cddip0_out_ia_rdata[21], \cddip0_out_ia_rdata.f.unused1 [6]);
tran (cddip0_out_ia_rdata[20], \cddip0_out_ia_rdata.r.part0 [20]);
tran (cddip0_out_ia_rdata[20], \cddip0_out_ia_rdata.f.unused1 [5]);
tran (cddip0_out_ia_rdata[19], \cddip0_out_ia_rdata.r.part0 [19]);
tran (cddip0_out_ia_rdata[19], \cddip0_out_ia_rdata.f.unused1 [4]);
tran (cddip0_out_ia_rdata[18], \cddip0_out_ia_rdata.r.part0 [18]);
tran (cddip0_out_ia_rdata[18], \cddip0_out_ia_rdata.f.unused1 [3]);
tran (cddip0_out_ia_rdata[17], \cddip0_out_ia_rdata.r.part0 [17]);
tran (cddip0_out_ia_rdata[17], \cddip0_out_ia_rdata.f.unused1 [2]);
tran (cddip0_out_ia_rdata[16], \cddip0_out_ia_rdata.r.part0 [16]);
tran (cddip0_out_ia_rdata[16], \cddip0_out_ia_rdata.f.unused1 [1]);
tran (cddip0_out_ia_rdata[15], \cddip0_out_ia_rdata.r.part0 [15]);
tran (cddip0_out_ia_rdata[15], \cddip0_out_ia_rdata.f.unused1 [0]);
tran (cddip0_out_ia_rdata[14], \cddip0_out_ia_rdata.r.part0 [14]);
tran (cddip0_out_ia_rdata[14], \cddip0_out_ia_rdata.f.tid );
tran (cddip0_out_ia_rdata[13], \cddip0_out_ia_rdata.r.part0 [13]);
tran (cddip0_out_ia_rdata[13], \cddip0_out_ia_rdata.f.tuser [7]);
tran (cddip0_out_ia_rdata[12], \cddip0_out_ia_rdata.r.part0 [12]);
tran (cddip0_out_ia_rdata[12], \cddip0_out_ia_rdata.f.tuser [6]);
tran (cddip0_out_ia_rdata[11], \cddip0_out_ia_rdata.r.part0 [11]);
tran (cddip0_out_ia_rdata[11], \cddip0_out_ia_rdata.f.tuser [5]);
tran (cddip0_out_ia_rdata[10], \cddip0_out_ia_rdata.r.part0 [10]);
tran (cddip0_out_ia_rdata[10], \cddip0_out_ia_rdata.f.tuser [4]);
tran (cddip0_out_ia_rdata[9], \cddip0_out_ia_rdata.r.part0 [9]);
tran (cddip0_out_ia_rdata[9], \cddip0_out_ia_rdata.f.tuser [3]);
tran (cddip0_out_ia_rdata[8], \cddip0_out_ia_rdata.r.part0 [8]);
tran (cddip0_out_ia_rdata[8], \cddip0_out_ia_rdata.f.tuser [2]);
tran (cddip0_out_ia_rdata[7], \cddip0_out_ia_rdata.r.part0 [7]);
tran (cddip0_out_ia_rdata[7], \cddip0_out_ia_rdata.f.tuser [1]);
tran (cddip0_out_ia_rdata[6], \cddip0_out_ia_rdata.r.part0 [6]);
tran (cddip0_out_ia_rdata[6], \cddip0_out_ia_rdata.f.tuser [0]);
tran (cddip0_out_ia_rdata[5], \cddip0_out_ia_rdata.r.part0 [5]);
tran (cddip0_out_ia_rdata[5], \cddip0_out_ia_rdata.f.unused0 [5]);
tran (cddip0_out_ia_rdata[4], \cddip0_out_ia_rdata.r.part0 [4]);
tran (cddip0_out_ia_rdata[4], \cddip0_out_ia_rdata.f.unused0 [4]);
tran (cddip0_out_ia_rdata[3], \cddip0_out_ia_rdata.r.part0 [3]);
tran (cddip0_out_ia_rdata[3], \cddip0_out_ia_rdata.f.unused0 [3]);
tran (cddip0_out_ia_rdata[2], \cddip0_out_ia_rdata.r.part0 [2]);
tran (cddip0_out_ia_rdata[2], \cddip0_out_ia_rdata.f.unused0 [2]);
tran (cddip0_out_ia_rdata[1], \cddip0_out_ia_rdata.r.part0 [1]);
tran (cddip0_out_ia_rdata[1], \cddip0_out_ia_rdata.f.unused0 [1]);
tran (cddip0_out_ia_rdata[0], \cddip0_out_ia_rdata.r.part0 [0]);
tran (cddip0_out_ia_rdata[0], \cddip0_out_ia_rdata.f.unused0 [0]);
tran (cddip0_out_im_status[11], \cddip0_out_im_status.r.part0 [11]);
tran (cddip0_out_im_status[11], \cddip0_out_im_status.f.bank_hi );
tran (cddip0_out_im_status[10], \cddip0_out_im_status.r.part0 [10]);
tran (cddip0_out_im_status[10], \cddip0_out_im_status.f.bank_lo );
tran (cddip0_out_im_status[9], \cddip0_out_im_status.r.part0 [9]);
tran (cddip0_out_im_status[9], \cddip0_out_im_status.f.overflow );
tran (cddip0_out_im_status[8], \cddip0_out_im_status.r.part0 [8]);
tran (cddip0_out_im_status[8], \cddip0_out_im_status.f.wr_pointer [8]);
tran (cddip0_out_im_status[7], \cddip0_out_im_status.r.part0 [7]);
tran (cddip0_out_im_status[7], \cddip0_out_im_status.f.wr_pointer [7]);
tran (cddip0_out_im_status[6], \cddip0_out_im_status.r.part0 [6]);
tran (cddip0_out_im_status[6], \cddip0_out_im_status.f.wr_pointer [6]);
tran (cddip0_out_im_status[5], \cddip0_out_im_status.r.part0 [5]);
tran (cddip0_out_im_status[5], \cddip0_out_im_status.f.wr_pointer [5]);
tran (cddip0_out_im_status[4], \cddip0_out_im_status.r.part0 [4]);
tran (cddip0_out_im_status[4], \cddip0_out_im_status.f.wr_pointer [4]);
tran (cddip0_out_im_status[3], \cddip0_out_im_status.r.part0 [3]);
tran (cddip0_out_im_status[3], \cddip0_out_im_status.f.wr_pointer [3]);
tran (cddip0_out_im_status[2], \cddip0_out_im_status.r.part0 [2]);
tran (cddip0_out_im_status[2], \cddip0_out_im_status.f.wr_pointer [2]);
tran (cddip0_out_im_status[1], \cddip0_out_im_status.r.part0 [1]);
tran (cddip0_out_im_status[1], \cddip0_out_im_status.f.wr_pointer [1]);
tran (cddip0_out_im_status[0], \cddip0_out_im_status.r.part0 [0]);
tran (cddip0_out_im_status[0], \cddip0_out_im_status.f.wr_pointer [0]);
tran (cddip1_out_ia_status[16], \cddip1_out_ia_status.r.part0 [16]);
tran (cddip1_out_ia_status[16], \cddip1_out_ia_status.f.code [2]);
tran (cddip1_out_ia_status[15], \cddip1_out_ia_status.r.part0 [15]);
tran (cddip1_out_ia_status[15], \cddip1_out_ia_status.f.code [1]);
tran (cddip1_out_ia_status[14], \cddip1_out_ia_status.r.part0 [14]);
tran (cddip1_out_ia_status[14], \cddip1_out_ia_status.f.code [0]);
tran (cddip1_out_ia_status[13], \cddip1_out_ia_status.r.part0 [13]);
tran (cddip1_out_ia_status[13], \cddip1_out_ia_status.f.datawords [4]);
tran (cddip1_out_ia_status[12], \cddip1_out_ia_status.r.part0 [12]);
tran (cddip1_out_ia_status[12], \cddip1_out_ia_status.f.datawords [3]);
tran (cddip1_out_ia_status[11], \cddip1_out_ia_status.r.part0 [11]);
tran (cddip1_out_ia_status[11], \cddip1_out_ia_status.f.datawords [2]);
tran (cddip1_out_ia_status[10], \cddip1_out_ia_status.r.part0 [10]);
tran (cddip1_out_ia_status[10], \cddip1_out_ia_status.f.datawords [1]);
tran (cddip1_out_ia_status[9], \cddip1_out_ia_status.r.part0 [9]);
tran (cddip1_out_ia_status[9], \cddip1_out_ia_status.f.datawords [0]);
tran (cddip1_out_ia_status[8], \cddip1_out_ia_status.r.part0 [8]);
tran (cddip1_out_ia_status[8], \cddip1_out_ia_status.f.addr [8]);
tran (cddip1_out_ia_status[7], \cddip1_out_ia_status.r.part0 [7]);
tran (cddip1_out_ia_status[7], \cddip1_out_ia_status.f.addr [7]);
tran (cddip1_out_ia_status[6], \cddip1_out_ia_status.r.part0 [6]);
tran (cddip1_out_ia_status[6], \cddip1_out_ia_status.f.addr [6]);
tran (cddip1_out_ia_status[5], \cddip1_out_ia_status.r.part0 [5]);
tran (cddip1_out_ia_status[5], \cddip1_out_ia_status.f.addr [5]);
tran (cddip1_out_ia_status[4], \cddip1_out_ia_status.r.part0 [4]);
tran (cddip1_out_ia_status[4], \cddip1_out_ia_status.f.addr [4]);
tran (cddip1_out_ia_status[3], \cddip1_out_ia_status.r.part0 [3]);
tran (cddip1_out_ia_status[3], \cddip1_out_ia_status.f.addr [3]);
tran (cddip1_out_ia_status[2], \cddip1_out_ia_status.r.part0 [2]);
tran (cddip1_out_ia_status[2], \cddip1_out_ia_status.f.addr [2]);
tran (cddip1_out_ia_status[1], \cddip1_out_ia_status.r.part0 [1]);
tran (cddip1_out_ia_status[1], \cddip1_out_ia_status.f.addr [1]);
tran (cddip1_out_ia_status[0], \cddip1_out_ia_status.r.part0 [0]);
tran (cddip1_out_ia_status[0], \cddip1_out_ia_status.f.addr [0]);
tran (cddip1_out_ia_capability[15], \cddip1_out_ia_capability.r.part0 [15]);
tran (cddip1_out_ia_capability[15], \cddip1_out_ia_capability.f.ack_error );
tran (cddip1_out_ia_capability[14], \cddip1_out_ia_capability.r.part0 [14]);
tran (cddip1_out_ia_capability[14], \cddip1_out_ia_capability.f.sim_tmo );
tran (cddip1_out_ia_capability[13], \cddip1_out_ia_capability.r.part0 [13]);
tran (cddip1_out_ia_capability[13], \cddip1_out_ia_capability.f.reserved_op [3]);
tran (cddip1_out_ia_capability[12], \cddip1_out_ia_capability.r.part0 [12]);
tran (cddip1_out_ia_capability[12], \cddip1_out_ia_capability.f.reserved_op [2]);
tran (cddip1_out_ia_capability[11], \cddip1_out_ia_capability.r.part0 [11]);
tran (cddip1_out_ia_capability[11], \cddip1_out_ia_capability.f.reserved_op [1]);
tran (cddip1_out_ia_capability[10], \cddip1_out_ia_capability.r.part0 [10]);
tran (cddip1_out_ia_capability[10], \cddip1_out_ia_capability.f.reserved_op [0]);
tran (cddip1_out_ia_capability[9], \cddip1_out_ia_capability.r.part0 [9]);
tran (cddip1_out_ia_capability[9], \cddip1_out_ia_capability.f.compare );
tran (cddip1_out_ia_capability[8], \cddip1_out_ia_capability.r.part0 [8]);
tran (cddip1_out_ia_capability[8], \cddip1_out_ia_capability.f.set_init_start );
tran (cddip1_out_ia_capability[7], \cddip1_out_ia_capability.r.part0 [7]);
tran (cddip1_out_ia_capability[7], \cddip1_out_ia_capability.f.initialize_inc );
tran (cddip1_out_ia_capability[6], \cddip1_out_ia_capability.r.part0 [6]);
tran (cddip1_out_ia_capability[6], \cddip1_out_ia_capability.f.initialize );
tran (cddip1_out_ia_capability[5], \cddip1_out_ia_capability.r.part0 [5]);
tran (cddip1_out_ia_capability[5], \cddip1_out_ia_capability.f.reset );
tran (cddip1_out_ia_capability[4], \cddip1_out_ia_capability.r.part0 [4]);
tran (cddip1_out_ia_capability[4], \cddip1_out_ia_capability.f.disabled );
tran (cddip1_out_ia_capability[3], \cddip1_out_ia_capability.r.part0 [3]);
tran (cddip1_out_ia_capability[3], \cddip1_out_ia_capability.f.enable );
tran (cddip1_out_ia_capability[2], \cddip1_out_ia_capability.r.part0 [2]);
tran (cddip1_out_ia_capability[2], \cddip1_out_ia_capability.f.write );
tran (cddip1_out_ia_capability[1], \cddip1_out_ia_capability.r.part0 [1]);
tran (cddip1_out_ia_capability[1], \cddip1_out_ia_capability.f.read );
tran (cddip1_out_ia_capability[0], \cddip1_out_ia_capability.r.part0 [0]);
tran (cddip1_out_ia_capability[0], \cddip1_out_ia_capability.f.nop );
tran (cddip1_out_ia_capability[19], \cddip1_out_ia_capability.r.part0 [19]);
tran (cddip1_out_ia_capability[19], \cddip1_out_ia_capability.f.mem_type [3]);
tran (cddip1_out_ia_capability[18], \cddip1_out_ia_capability.r.part0 [18]);
tran (cddip1_out_ia_capability[18], \cddip1_out_ia_capability.f.mem_type [2]);
tran (cddip1_out_ia_capability[17], \cddip1_out_ia_capability.r.part0 [17]);
tran (cddip1_out_ia_capability[17], \cddip1_out_ia_capability.f.mem_type [1]);
tran (cddip1_out_ia_capability[16], \cddip1_out_ia_capability.r.part0 [16]);
tran (cddip1_out_ia_capability[16], \cddip1_out_ia_capability.f.mem_type [0]);
tran (cddip1_out_ia_rdata[95], \cddip1_out_ia_rdata.r.part2 [31]);
tran (cddip1_out_ia_rdata[95], \cddip1_out_ia_rdata.f.tdata_hi [31]);
tran (cddip1_out_ia_rdata[94], \cddip1_out_ia_rdata.r.part2 [30]);
tran (cddip1_out_ia_rdata[94], \cddip1_out_ia_rdata.f.tdata_hi [30]);
tran (cddip1_out_ia_rdata[93], \cddip1_out_ia_rdata.r.part2 [29]);
tran (cddip1_out_ia_rdata[93], \cddip1_out_ia_rdata.f.tdata_hi [29]);
tran (cddip1_out_ia_rdata[92], \cddip1_out_ia_rdata.r.part2 [28]);
tran (cddip1_out_ia_rdata[92], \cddip1_out_ia_rdata.f.tdata_hi [28]);
tran (cddip1_out_ia_rdata[91], \cddip1_out_ia_rdata.r.part2 [27]);
tran (cddip1_out_ia_rdata[91], \cddip1_out_ia_rdata.f.tdata_hi [27]);
tran (cddip1_out_ia_rdata[90], \cddip1_out_ia_rdata.r.part2 [26]);
tran (cddip1_out_ia_rdata[90], \cddip1_out_ia_rdata.f.tdata_hi [26]);
tran (cddip1_out_ia_rdata[89], \cddip1_out_ia_rdata.r.part2 [25]);
tran (cddip1_out_ia_rdata[89], \cddip1_out_ia_rdata.f.tdata_hi [25]);
tran (cddip1_out_ia_rdata[88], \cddip1_out_ia_rdata.r.part2 [24]);
tran (cddip1_out_ia_rdata[88], \cddip1_out_ia_rdata.f.tdata_hi [24]);
tran (cddip1_out_ia_rdata[87], \cddip1_out_ia_rdata.r.part2 [23]);
tran (cddip1_out_ia_rdata[87], \cddip1_out_ia_rdata.f.tdata_hi [23]);
tran (cddip1_out_ia_rdata[86], \cddip1_out_ia_rdata.r.part2 [22]);
tran (cddip1_out_ia_rdata[86], \cddip1_out_ia_rdata.f.tdata_hi [22]);
tran (cddip1_out_ia_rdata[85], \cddip1_out_ia_rdata.r.part2 [21]);
tran (cddip1_out_ia_rdata[85], \cddip1_out_ia_rdata.f.tdata_hi [21]);
tran (cddip1_out_ia_rdata[84], \cddip1_out_ia_rdata.r.part2 [20]);
tran (cddip1_out_ia_rdata[84], \cddip1_out_ia_rdata.f.tdata_hi [20]);
tran (cddip1_out_ia_rdata[83], \cddip1_out_ia_rdata.r.part2 [19]);
tran (cddip1_out_ia_rdata[83], \cddip1_out_ia_rdata.f.tdata_hi [19]);
tran (cddip1_out_ia_rdata[82], \cddip1_out_ia_rdata.r.part2 [18]);
tran (cddip1_out_ia_rdata[82], \cddip1_out_ia_rdata.f.tdata_hi [18]);
tran (cddip1_out_ia_rdata[81], \cddip1_out_ia_rdata.r.part2 [17]);
tran (cddip1_out_ia_rdata[81], \cddip1_out_ia_rdata.f.tdata_hi [17]);
tran (cddip1_out_ia_rdata[80], \cddip1_out_ia_rdata.r.part2 [16]);
tran (cddip1_out_ia_rdata[80], \cddip1_out_ia_rdata.f.tdata_hi [16]);
tran (cddip1_out_ia_rdata[79], \cddip1_out_ia_rdata.r.part2 [15]);
tran (cddip1_out_ia_rdata[79], \cddip1_out_ia_rdata.f.tdata_hi [15]);
tran (cddip1_out_ia_rdata[78], \cddip1_out_ia_rdata.r.part2 [14]);
tran (cddip1_out_ia_rdata[78], \cddip1_out_ia_rdata.f.tdata_hi [14]);
tran (cddip1_out_ia_rdata[77], \cddip1_out_ia_rdata.r.part2 [13]);
tran (cddip1_out_ia_rdata[77], \cddip1_out_ia_rdata.f.tdata_hi [13]);
tran (cddip1_out_ia_rdata[76], \cddip1_out_ia_rdata.r.part2 [12]);
tran (cddip1_out_ia_rdata[76], \cddip1_out_ia_rdata.f.tdata_hi [12]);
tran (cddip1_out_ia_rdata[75], \cddip1_out_ia_rdata.r.part2 [11]);
tran (cddip1_out_ia_rdata[75], \cddip1_out_ia_rdata.f.tdata_hi [11]);
tran (cddip1_out_ia_rdata[74], \cddip1_out_ia_rdata.r.part2 [10]);
tran (cddip1_out_ia_rdata[74], \cddip1_out_ia_rdata.f.tdata_hi [10]);
tran (cddip1_out_ia_rdata[73], \cddip1_out_ia_rdata.r.part2 [9]);
tran (cddip1_out_ia_rdata[73], \cddip1_out_ia_rdata.f.tdata_hi [9]);
tran (cddip1_out_ia_rdata[72], \cddip1_out_ia_rdata.r.part2 [8]);
tran (cddip1_out_ia_rdata[72], \cddip1_out_ia_rdata.f.tdata_hi [8]);
tran (cddip1_out_ia_rdata[71], \cddip1_out_ia_rdata.r.part2 [7]);
tran (cddip1_out_ia_rdata[71], \cddip1_out_ia_rdata.f.tdata_hi [7]);
tran (cddip1_out_ia_rdata[70], \cddip1_out_ia_rdata.r.part2 [6]);
tran (cddip1_out_ia_rdata[70], \cddip1_out_ia_rdata.f.tdata_hi [6]);
tran (cddip1_out_ia_rdata[69], \cddip1_out_ia_rdata.r.part2 [5]);
tran (cddip1_out_ia_rdata[69], \cddip1_out_ia_rdata.f.tdata_hi [5]);
tran (cddip1_out_ia_rdata[68], \cddip1_out_ia_rdata.r.part2 [4]);
tran (cddip1_out_ia_rdata[68], \cddip1_out_ia_rdata.f.tdata_hi [4]);
tran (cddip1_out_ia_rdata[67], \cddip1_out_ia_rdata.r.part2 [3]);
tran (cddip1_out_ia_rdata[67], \cddip1_out_ia_rdata.f.tdata_hi [3]);
tran (cddip1_out_ia_rdata[66], \cddip1_out_ia_rdata.r.part2 [2]);
tran (cddip1_out_ia_rdata[66], \cddip1_out_ia_rdata.f.tdata_hi [2]);
tran (cddip1_out_ia_rdata[65], \cddip1_out_ia_rdata.r.part2 [1]);
tran (cddip1_out_ia_rdata[65], \cddip1_out_ia_rdata.f.tdata_hi [1]);
tran (cddip1_out_ia_rdata[64], \cddip1_out_ia_rdata.r.part2 [0]);
tran (cddip1_out_ia_rdata[64], \cddip1_out_ia_rdata.f.tdata_hi [0]);
tran (cddip1_out_ia_rdata[63], \cddip1_out_ia_rdata.r.part1 [31]);
tran (cddip1_out_ia_rdata[63], \cddip1_out_ia_rdata.f.tdata_lo [31]);
tran (cddip1_out_ia_rdata[62], \cddip1_out_ia_rdata.r.part1 [30]);
tran (cddip1_out_ia_rdata[62], \cddip1_out_ia_rdata.f.tdata_lo [30]);
tran (cddip1_out_ia_rdata[61], \cddip1_out_ia_rdata.r.part1 [29]);
tran (cddip1_out_ia_rdata[61], \cddip1_out_ia_rdata.f.tdata_lo [29]);
tran (cddip1_out_ia_rdata[60], \cddip1_out_ia_rdata.r.part1 [28]);
tran (cddip1_out_ia_rdata[60], \cddip1_out_ia_rdata.f.tdata_lo [28]);
tran (cddip1_out_ia_rdata[59], \cddip1_out_ia_rdata.r.part1 [27]);
tran (cddip1_out_ia_rdata[59], \cddip1_out_ia_rdata.f.tdata_lo [27]);
tran (cddip1_out_ia_rdata[58], \cddip1_out_ia_rdata.r.part1 [26]);
tran (cddip1_out_ia_rdata[58], \cddip1_out_ia_rdata.f.tdata_lo [26]);
tran (cddip1_out_ia_rdata[57], \cddip1_out_ia_rdata.r.part1 [25]);
tran (cddip1_out_ia_rdata[57], \cddip1_out_ia_rdata.f.tdata_lo [25]);
tran (cddip1_out_ia_rdata[56], \cddip1_out_ia_rdata.r.part1 [24]);
tran (cddip1_out_ia_rdata[56], \cddip1_out_ia_rdata.f.tdata_lo [24]);
tran (cddip1_out_ia_rdata[55], \cddip1_out_ia_rdata.r.part1 [23]);
tran (cddip1_out_ia_rdata[55], \cddip1_out_ia_rdata.f.tdata_lo [23]);
tran (cddip1_out_ia_rdata[54], \cddip1_out_ia_rdata.r.part1 [22]);
tran (cddip1_out_ia_rdata[54], \cddip1_out_ia_rdata.f.tdata_lo [22]);
tran (cddip1_out_ia_rdata[53], \cddip1_out_ia_rdata.r.part1 [21]);
tran (cddip1_out_ia_rdata[53], \cddip1_out_ia_rdata.f.tdata_lo [21]);
tran (cddip1_out_ia_rdata[52], \cddip1_out_ia_rdata.r.part1 [20]);
tran (cddip1_out_ia_rdata[52], \cddip1_out_ia_rdata.f.tdata_lo [20]);
tran (cddip1_out_ia_rdata[51], \cddip1_out_ia_rdata.r.part1 [19]);
tran (cddip1_out_ia_rdata[51], \cddip1_out_ia_rdata.f.tdata_lo [19]);
tran (cddip1_out_ia_rdata[50], \cddip1_out_ia_rdata.r.part1 [18]);
tran (cddip1_out_ia_rdata[50], \cddip1_out_ia_rdata.f.tdata_lo [18]);
tran (cddip1_out_ia_rdata[49], \cddip1_out_ia_rdata.r.part1 [17]);
tran (cddip1_out_ia_rdata[49], \cddip1_out_ia_rdata.f.tdata_lo [17]);
tran (cddip1_out_ia_rdata[48], \cddip1_out_ia_rdata.r.part1 [16]);
tran (cddip1_out_ia_rdata[48], \cddip1_out_ia_rdata.f.tdata_lo [16]);
tran (cddip1_out_ia_rdata[47], \cddip1_out_ia_rdata.r.part1 [15]);
tran (cddip1_out_ia_rdata[47], \cddip1_out_ia_rdata.f.tdata_lo [15]);
tran (cddip1_out_ia_rdata[46], \cddip1_out_ia_rdata.r.part1 [14]);
tran (cddip1_out_ia_rdata[46], \cddip1_out_ia_rdata.f.tdata_lo [14]);
tran (cddip1_out_ia_rdata[45], \cddip1_out_ia_rdata.r.part1 [13]);
tran (cddip1_out_ia_rdata[45], \cddip1_out_ia_rdata.f.tdata_lo [13]);
tran (cddip1_out_ia_rdata[44], \cddip1_out_ia_rdata.r.part1 [12]);
tran (cddip1_out_ia_rdata[44], \cddip1_out_ia_rdata.f.tdata_lo [12]);
tran (cddip1_out_ia_rdata[43], \cddip1_out_ia_rdata.r.part1 [11]);
tran (cddip1_out_ia_rdata[43], \cddip1_out_ia_rdata.f.tdata_lo [11]);
tran (cddip1_out_ia_rdata[42], \cddip1_out_ia_rdata.r.part1 [10]);
tran (cddip1_out_ia_rdata[42], \cddip1_out_ia_rdata.f.tdata_lo [10]);
tran (cddip1_out_ia_rdata[41], \cddip1_out_ia_rdata.r.part1 [9]);
tran (cddip1_out_ia_rdata[41], \cddip1_out_ia_rdata.f.tdata_lo [9]);
tran (cddip1_out_ia_rdata[40], \cddip1_out_ia_rdata.r.part1 [8]);
tran (cddip1_out_ia_rdata[40], \cddip1_out_ia_rdata.f.tdata_lo [8]);
tran (cddip1_out_ia_rdata[39], \cddip1_out_ia_rdata.r.part1 [7]);
tran (cddip1_out_ia_rdata[39], \cddip1_out_ia_rdata.f.tdata_lo [7]);
tran (cddip1_out_ia_rdata[38], \cddip1_out_ia_rdata.r.part1 [6]);
tran (cddip1_out_ia_rdata[38], \cddip1_out_ia_rdata.f.tdata_lo [6]);
tran (cddip1_out_ia_rdata[37], \cddip1_out_ia_rdata.r.part1 [5]);
tran (cddip1_out_ia_rdata[37], \cddip1_out_ia_rdata.f.tdata_lo [5]);
tran (cddip1_out_ia_rdata[36], \cddip1_out_ia_rdata.r.part1 [4]);
tran (cddip1_out_ia_rdata[36], \cddip1_out_ia_rdata.f.tdata_lo [4]);
tran (cddip1_out_ia_rdata[35], \cddip1_out_ia_rdata.r.part1 [3]);
tran (cddip1_out_ia_rdata[35], \cddip1_out_ia_rdata.f.tdata_lo [3]);
tran (cddip1_out_ia_rdata[34], \cddip1_out_ia_rdata.r.part1 [2]);
tran (cddip1_out_ia_rdata[34], \cddip1_out_ia_rdata.f.tdata_lo [2]);
tran (cddip1_out_ia_rdata[33], \cddip1_out_ia_rdata.r.part1 [1]);
tran (cddip1_out_ia_rdata[33], \cddip1_out_ia_rdata.f.tdata_lo [1]);
tran (cddip1_out_ia_rdata[32], \cddip1_out_ia_rdata.r.part1 [0]);
tran (cddip1_out_ia_rdata[32], \cddip1_out_ia_rdata.f.tdata_lo [0]);
tran (cddip1_out_ia_rdata[31], \cddip1_out_ia_rdata.r.part0 [31]);
tran (cddip1_out_ia_rdata[31], \cddip1_out_ia_rdata.f.eob );
tran (cddip1_out_ia_rdata[30], \cddip1_out_ia_rdata.r.part0 [30]);
tran (cddip1_out_ia_rdata[30], \cddip1_out_ia_rdata.f.bytes_vld [7]);
tran (cddip1_out_ia_rdata[29], \cddip1_out_ia_rdata.r.part0 [29]);
tran (cddip1_out_ia_rdata[29], \cddip1_out_ia_rdata.f.bytes_vld [6]);
tran (cddip1_out_ia_rdata[28], \cddip1_out_ia_rdata.r.part0 [28]);
tran (cddip1_out_ia_rdata[28], \cddip1_out_ia_rdata.f.bytes_vld [5]);
tran (cddip1_out_ia_rdata[27], \cddip1_out_ia_rdata.r.part0 [27]);
tran (cddip1_out_ia_rdata[27], \cddip1_out_ia_rdata.f.bytes_vld [4]);
tran (cddip1_out_ia_rdata[26], \cddip1_out_ia_rdata.r.part0 [26]);
tran (cddip1_out_ia_rdata[26], \cddip1_out_ia_rdata.f.bytes_vld [3]);
tran (cddip1_out_ia_rdata[25], \cddip1_out_ia_rdata.r.part0 [25]);
tran (cddip1_out_ia_rdata[25], \cddip1_out_ia_rdata.f.bytes_vld [2]);
tran (cddip1_out_ia_rdata[24], \cddip1_out_ia_rdata.r.part0 [24]);
tran (cddip1_out_ia_rdata[24], \cddip1_out_ia_rdata.f.bytes_vld [1]);
tran (cddip1_out_ia_rdata[23], \cddip1_out_ia_rdata.r.part0 [23]);
tran (cddip1_out_ia_rdata[23], \cddip1_out_ia_rdata.f.bytes_vld [0]);
tran (cddip1_out_ia_rdata[22], \cddip1_out_ia_rdata.r.part0 [22]);
tran (cddip1_out_ia_rdata[22], \cddip1_out_ia_rdata.f.unused1 [7]);
tran (cddip1_out_ia_rdata[21], \cddip1_out_ia_rdata.r.part0 [21]);
tran (cddip1_out_ia_rdata[21], \cddip1_out_ia_rdata.f.unused1 [6]);
tran (cddip1_out_ia_rdata[20], \cddip1_out_ia_rdata.r.part0 [20]);
tran (cddip1_out_ia_rdata[20], \cddip1_out_ia_rdata.f.unused1 [5]);
tran (cddip1_out_ia_rdata[19], \cddip1_out_ia_rdata.r.part0 [19]);
tran (cddip1_out_ia_rdata[19], \cddip1_out_ia_rdata.f.unused1 [4]);
tran (cddip1_out_ia_rdata[18], \cddip1_out_ia_rdata.r.part0 [18]);
tran (cddip1_out_ia_rdata[18], \cddip1_out_ia_rdata.f.unused1 [3]);
tran (cddip1_out_ia_rdata[17], \cddip1_out_ia_rdata.r.part0 [17]);
tran (cddip1_out_ia_rdata[17], \cddip1_out_ia_rdata.f.unused1 [2]);
tran (cddip1_out_ia_rdata[16], \cddip1_out_ia_rdata.r.part0 [16]);
tran (cddip1_out_ia_rdata[16], \cddip1_out_ia_rdata.f.unused1 [1]);
tran (cddip1_out_ia_rdata[15], \cddip1_out_ia_rdata.r.part0 [15]);
tran (cddip1_out_ia_rdata[15], \cddip1_out_ia_rdata.f.unused1 [0]);
tran (cddip1_out_ia_rdata[14], \cddip1_out_ia_rdata.r.part0 [14]);
tran (cddip1_out_ia_rdata[14], \cddip1_out_ia_rdata.f.tid );
tran (cddip1_out_ia_rdata[13], \cddip1_out_ia_rdata.r.part0 [13]);
tran (cddip1_out_ia_rdata[13], \cddip1_out_ia_rdata.f.tuser [7]);
tran (cddip1_out_ia_rdata[12], \cddip1_out_ia_rdata.r.part0 [12]);
tran (cddip1_out_ia_rdata[12], \cddip1_out_ia_rdata.f.tuser [6]);
tran (cddip1_out_ia_rdata[11], \cddip1_out_ia_rdata.r.part0 [11]);
tran (cddip1_out_ia_rdata[11], \cddip1_out_ia_rdata.f.tuser [5]);
tran (cddip1_out_ia_rdata[10], \cddip1_out_ia_rdata.r.part0 [10]);
tran (cddip1_out_ia_rdata[10], \cddip1_out_ia_rdata.f.tuser [4]);
tran (cddip1_out_ia_rdata[9], \cddip1_out_ia_rdata.r.part0 [9]);
tran (cddip1_out_ia_rdata[9], \cddip1_out_ia_rdata.f.tuser [3]);
tran (cddip1_out_ia_rdata[8], \cddip1_out_ia_rdata.r.part0 [8]);
tran (cddip1_out_ia_rdata[8], \cddip1_out_ia_rdata.f.tuser [2]);
tran (cddip1_out_ia_rdata[7], \cddip1_out_ia_rdata.r.part0 [7]);
tran (cddip1_out_ia_rdata[7], \cddip1_out_ia_rdata.f.tuser [1]);
tran (cddip1_out_ia_rdata[6], \cddip1_out_ia_rdata.r.part0 [6]);
tran (cddip1_out_ia_rdata[6], \cddip1_out_ia_rdata.f.tuser [0]);
tran (cddip1_out_ia_rdata[5], \cddip1_out_ia_rdata.r.part0 [5]);
tran (cddip1_out_ia_rdata[5], \cddip1_out_ia_rdata.f.unused0 [5]);
tran (cddip1_out_ia_rdata[4], \cddip1_out_ia_rdata.r.part0 [4]);
tran (cddip1_out_ia_rdata[4], \cddip1_out_ia_rdata.f.unused0 [4]);
tran (cddip1_out_ia_rdata[3], \cddip1_out_ia_rdata.r.part0 [3]);
tran (cddip1_out_ia_rdata[3], \cddip1_out_ia_rdata.f.unused0 [3]);
tran (cddip1_out_ia_rdata[2], \cddip1_out_ia_rdata.r.part0 [2]);
tran (cddip1_out_ia_rdata[2], \cddip1_out_ia_rdata.f.unused0 [2]);
tran (cddip1_out_ia_rdata[1], \cddip1_out_ia_rdata.r.part0 [1]);
tran (cddip1_out_ia_rdata[1], \cddip1_out_ia_rdata.f.unused0 [1]);
tran (cddip1_out_ia_rdata[0], \cddip1_out_ia_rdata.r.part0 [0]);
tran (cddip1_out_ia_rdata[0], \cddip1_out_ia_rdata.f.unused0 [0]);
tran (cddip1_out_im_status[11], \cddip1_out_im_status.r.part0 [11]);
tran (cddip1_out_im_status[11], \cddip1_out_im_status.f.bank_hi );
tran (cddip1_out_im_status[10], \cddip1_out_im_status.r.part0 [10]);
tran (cddip1_out_im_status[10], \cddip1_out_im_status.f.bank_lo );
tran (cddip1_out_im_status[9], \cddip1_out_im_status.r.part0 [9]);
tran (cddip1_out_im_status[9], \cddip1_out_im_status.f.overflow );
tran (cddip1_out_im_status[8], \cddip1_out_im_status.r.part0 [8]);
tran (cddip1_out_im_status[8], \cddip1_out_im_status.f.wr_pointer [8]);
tran (cddip1_out_im_status[7], \cddip1_out_im_status.r.part0 [7]);
tran (cddip1_out_im_status[7], \cddip1_out_im_status.f.wr_pointer [7]);
tran (cddip1_out_im_status[6], \cddip1_out_im_status.r.part0 [6]);
tran (cddip1_out_im_status[6], \cddip1_out_im_status.f.wr_pointer [6]);
tran (cddip1_out_im_status[5], \cddip1_out_im_status.r.part0 [5]);
tran (cddip1_out_im_status[5], \cddip1_out_im_status.f.wr_pointer [5]);
tran (cddip1_out_im_status[4], \cddip1_out_im_status.r.part0 [4]);
tran (cddip1_out_im_status[4], \cddip1_out_im_status.f.wr_pointer [4]);
tran (cddip1_out_im_status[3], \cddip1_out_im_status.r.part0 [3]);
tran (cddip1_out_im_status[3], \cddip1_out_im_status.f.wr_pointer [3]);
tran (cddip1_out_im_status[2], \cddip1_out_im_status.r.part0 [2]);
tran (cddip1_out_im_status[2], \cddip1_out_im_status.f.wr_pointer [2]);
tran (cddip1_out_im_status[1], \cddip1_out_im_status.r.part0 [1]);
tran (cddip1_out_im_status[1], \cddip1_out_im_status.f.wr_pointer [1]);
tran (cddip1_out_im_status[0], \cddip1_out_im_status.r.part0 [0]);
tran (cddip1_out_im_status[0], \cddip1_out_im_status.f.wr_pointer [0]);
tran (cddip2_out_ia_status[16], \cddip2_out_ia_status.r.part0 [16]);
tran (cddip2_out_ia_status[16], \cddip2_out_ia_status.f.code [2]);
tran (cddip2_out_ia_status[15], \cddip2_out_ia_status.r.part0 [15]);
tran (cddip2_out_ia_status[15], \cddip2_out_ia_status.f.code [1]);
tran (cddip2_out_ia_status[14], \cddip2_out_ia_status.r.part0 [14]);
tran (cddip2_out_ia_status[14], \cddip2_out_ia_status.f.code [0]);
tran (cddip2_out_ia_status[13], \cddip2_out_ia_status.r.part0 [13]);
tran (cddip2_out_ia_status[13], \cddip2_out_ia_status.f.datawords [4]);
tran (cddip2_out_ia_status[12], \cddip2_out_ia_status.r.part0 [12]);
tran (cddip2_out_ia_status[12], \cddip2_out_ia_status.f.datawords [3]);
tran (cddip2_out_ia_status[11], \cddip2_out_ia_status.r.part0 [11]);
tran (cddip2_out_ia_status[11], \cddip2_out_ia_status.f.datawords [2]);
tran (cddip2_out_ia_status[10], \cddip2_out_ia_status.r.part0 [10]);
tran (cddip2_out_ia_status[10], \cddip2_out_ia_status.f.datawords [1]);
tran (cddip2_out_ia_status[9], \cddip2_out_ia_status.r.part0 [9]);
tran (cddip2_out_ia_status[9], \cddip2_out_ia_status.f.datawords [0]);
tran (cddip2_out_ia_status[8], \cddip2_out_ia_status.r.part0 [8]);
tran (cddip2_out_ia_status[8], \cddip2_out_ia_status.f.addr [8]);
tran (cddip2_out_ia_status[7], \cddip2_out_ia_status.r.part0 [7]);
tran (cddip2_out_ia_status[7], \cddip2_out_ia_status.f.addr [7]);
tran (cddip2_out_ia_status[6], \cddip2_out_ia_status.r.part0 [6]);
tran (cddip2_out_ia_status[6], \cddip2_out_ia_status.f.addr [6]);
tran (cddip2_out_ia_status[5], \cddip2_out_ia_status.r.part0 [5]);
tran (cddip2_out_ia_status[5], \cddip2_out_ia_status.f.addr [5]);
tran (cddip2_out_ia_status[4], \cddip2_out_ia_status.r.part0 [4]);
tran (cddip2_out_ia_status[4], \cddip2_out_ia_status.f.addr [4]);
tran (cddip2_out_ia_status[3], \cddip2_out_ia_status.r.part0 [3]);
tran (cddip2_out_ia_status[3], \cddip2_out_ia_status.f.addr [3]);
tran (cddip2_out_ia_status[2], \cddip2_out_ia_status.r.part0 [2]);
tran (cddip2_out_ia_status[2], \cddip2_out_ia_status.f.addr [2]);
tran (cddip2_out_ia_status[1], \cddip2_out_ia_status.r.part0 [1]);
tran (cddip2_out_ia_status[1], \cddip2_out_ia_status.f.addr [1]);
tran (cddip2_out_ia_status[0], \cddip2_out_ia_status.r.part0 [0]);
tran (cddip2_out_ia_status[0], \cddip2_out_ia_status.f.addr [0]);
tran (cddip2_out_ia_capability[15], \cddip2_out_ia_capability.r.part0 [15]);
tran (cddip2_out_ia_capability[15], \cddip2_out_ia_capability.f.ack_error );
tran (cddip2_out_ia_capability[14], \cddip2_out_ia_capability.r.part0 [14]);
tran (cddip2_out_ia_capability[14], \cddip2_out_ia_capability.f.sim_tmo );
tran (cddip2_out_ia_capability[13], \cddip2_out_ia_capability.r.part0 [13]);
tran (cddip2_out_ia_capability[13], \cddip2_out_ia_capability.f.reserved_op [3]);
tran (cddip2_out_ia_capability[12], \cddip2_out_ia_capability.r.part0 [12]);
tran (cddip2_out_ia_capability[12], \cddip2_out_ia_capability.f.reserved_op [2]);
tran (cddip2_out_ia_capability[11], \cddip2_out_ia_capability.r.part0 [11]);
tran (cddip2_out_ia_capability[11], \cddip2_out_ia_capability.f.reserved_op [1]);
tran (cddip2_out_ia_capability[10], \cddip2_out_ia_capability.r.part0 [10]);
tran (cddip2_out_ia_capability[10], \cddip2_out_ia_capability.f.reserved_op [0]);
tran (cddip2_out_ia_capability[9], \cddip2_out_ia_capability.r.part0 [9]);
tran (cddip2_out_ia_capability[9], \cddip2_out_ia_capability.f.compare );
tran (cddip2_out_ia_capability[8], \cddip2_out_ia_capability.r.part0 [8]);
tran (cddip2_out_ia_capability[8], \cddip2_out_ia_capability.f.set_init_start );
tran (cddip2_out_ia_capability[7], \cddip2_out_ia_capability.r.part0 [7]);
tran (cddip2_out_ia_capability[7], \cddip2_out_ia_capability.f.initialize_inc );
tran (cddip2_out_ia_capability[6], \cddip2_out_ia_capability.r.part0 [6]);
tran (cddip2_out_ia_capability[6], \cddip2_out_ia_capability.f.initialize );
tran (cddip2_out_ia_capability[5], \cddip2_out_ia_capability.r.part0 [5]);
tran (cddip2_out_ia_capability[5], \cddip2_out_ia_capability.f.reset );
tran (cddip2_out_ia_capability[4], \cddip2_out_ia_capability.r.part0 [4]);
tran (cddip2_out_ia_capability[4], \cddip2_out_ia_capability.f.disabled );
tran (cddip2_out_ia_capability[3], \cddip2_out_ia_capability.r.part0 [3]);
tran (cddip2_out_ia_capability[3], \cddip2_out_ia_capability.f.enable );
tran (cddip2_out_ia_capability[2], \cddip2_out_ia_capability.r.part0 [2]);
tran (cddip2_out_ia_capability[2], \cddip2_out_ia_capability.f.write );
tran (cddip2_out_ia_capability[1], \cddip2_out_ia_capability.r.part0 [1]);
tran (cddip2_out_ia_capability[1], \cddip2_out_ia_capability.f.read );
tran (cddip2_out_ia_capability[0], \cddip2_out_ia_capability.r.part0 [0]);
tran (cddip2_out_ia_capability[0], \cddip2_out_ia_capability.f.nop );
tran (cddip2_out_ia_capability[19], \cddip2_out_ia_capability.r.part0 [19]);
tran (cddip2_out_ia_capability[19], \cddip2_out_ia_capability.f.mem_type [3]);
tran (cddip2_out_ia_capability[18], \cddip2_out_ia_capability.r.part0 [18]);
tran (cddip2_out_ia_capability[18], \cddip2_out_ia_capability.f.mem_type [2]);
tran (cddip2_out_ia_capability[17], \cddip2_out_ia_capability.r.part0 [17]);
tran (cddip2_out_ia_capability[17], \cddip2_out_ia_capability.f.mem_type [1]);
tran (cddip2_out_ia_capability[16], \cddip2_out_ia_capability.r.part0 [16]);
tran (cddip2_out_ia_capability[16], \cddip2_out_ia_capability.f.mem_type [0]);
tran (cddip2_out_ia_rdata[95], \cddip2_out_ia_rdata.r.part2 [31]);
tran (cddip2_out_ia_rdata[95], \cddip2_out_ia_rdata.f.tdata_hi [31]);
tran (cddip2_out_ia_rdata[94], \cddip2_out_ia_rdata.r.part2 [30]);
tran (cddip2_out_ia_rdata[94], \cddip2_out_ia_rdata.f.tdata_hi [30]);
tran (cddip2_out_ia_rdata[93], \cddip2_out_ia_rdata.r.part2 [29]);
tran (cddip2_out_ia_rdata[93], \cddip2_out_ia_rdata.f.tdata_hi [29]);
tran (cddip2_out_ia_rdata[92], \cddip2_out_ia_rdata.r.part2 [28]);
tran (cddip2_out_ia_rdata[92], \cddip2_out_ia_rdata.f.tdata_hi [28]);
tran (cddip2_out_ia_rdata[91], \cddip2_out_ia_rdata.r.part2 [27]);
tran (cddip2_out_ia_rdata[91], \cddip2_out_ia_rdata.f.tdata_hi [27]);
tran (cddip2_out_ia_rdata[90], \cddip2_out_ia_rdata.r.part2 [26]);
tran (cddip2_out_ia_rdata[90], \cddip2_out_ia_rdata.f.tdata_hi [26]);
tran (cddip2_out_ia_rdata[89], \cddip2_out_ia_rdata.r.part2 [25]);
tran (cddip2_out_ia_rdata[89], \cddip2_out_ia_rdata.f.tdata_hi [25]);
tran (cddip2_out_ia_rdata[88], \cddip2_out_ia_rdata.r.part2 [24]);
tran (cddip2_out_ia_rdata[88], \cddip2_out_ia_rdata.f.tdata_hi [24]);
tran (cddip2_out_ia_rdata[87], \cddip2_out_ia_rdata.r.part2 [23]);
tran (cddip2_out_ia_rdata[87], \cddip2_out_ia_rdata.f.tdata_hi [23]);
tran (cddip2_out_ia_rdata[86], \cddip2_out_ia_rdata.r.part2 [22]);
tran (cddip2_out_ia_rdata[86], \cddip2_out_ia_rdata.f.tdata_hi [22]);
tran (cddip2_out_ia_rdata[85], \cddip2_out_ia_rdata.r.part2 [21]);
tran (cddip2_out_ia_rdata[85], \cddip2_out_ia_rdata.f.tdata_hi [21]);
tran (cddip2_out_ia_rdata[84], \cddip2_out_ia_rdata.r.part2 [20]);
tran (cddip2_out_ia_rdata[84], \cddip2_out_ia_rdata.f.tdata_hi [20]);
tran (cddip2_out_ia_rdata[83], \cddip2_out_ia_rdata.r.part2 [19]);
tran (cddip2_out_ia_rdata[83], \cddip2_out_ia_rdata.f.tdata_hi [19]);
tran (cddip2_out_ia_rdata[82], \cddip2_out_ia_rdata.r.part2 [18]);
tran (cddip2_out_ia_rdata[82], \cddip2_out_ia_rdata.f.tdata_hi [18]);
tran (cddip2_out_ia_rdata[81], \cddip2_out_ia_rdata.r.part2 [17]);
tran (cddip2_out_ia_rdata[81], \cddip2_out_ia_rdata.f.tdata_hi [17]);
tran (cddip2_out_ia_rdata[80], \cddip2_out_ia_rdata.r.part2 [16]);
tran (cddip2_out_ia_rdata[80], \cddip2_out_ia_rdata.f.tdata_hi [16]);
tran (cddip2_out_ia_rdata[79], \cddip2_out_ia_rdata.r.part2 [15]);
tran (cddip2_out_ia_rdata[79], \cddip2_out_ia_rdata.f.tdata_hi [15]);
tran (cddip2_out_ia_rdata[78], \cddip2_out_ia_rdata.r.part2 [14]);
tran (cddip2_out_ia_rdata[78], \cddip2_out_ia_rdata.f.tdata_hi [14]);
tran (cddip2_out_ia_rdata[77], \cddip2_out_ia_rdata.r.part2 [13]);
tran (cddip2_out_ia_rdata[77], \cddip2_out_ia_rdata.f.tdata_hi [13]);
tran (cddip2_out_ia_rdata[76], \cddip2_out_ia_rdata.r.part2 [12]);
tran (cddip2_out_ia_rdata[76], \cddip2_out_ia_rdata.f.tdata_hi [12]);
tran (cddip2_out_ia_rdata[75], \cddip2_out_ia_rdata.r.part2 [11]);
tran (cddip2_out_ia_rdata[75], \cddip2_out_ia_rdata.f.tdata_hi [11]);
tran (cddip2_out_ia_rdata[74], \cddip2_out_ia_rdata.r.part2 [10]);
tran (cddip2_out_ia_rdata[74], \cddip2_out_ia_rdata.f.tdata_hi [10]);
tran (cddip2_out_ia_rdata[73], \cddip2_out_ia_rdata.r.part2 [9]);
tran (cddip2_out_ia_rdata[73], \cddip2_out_ia_rdata.f.tdata_hi [9]);
tran (cddip2_out_ia_rdata[72], \cddip2_out_ia_rdata.r.part2 [8]);
tran (cddip2_out_ia_rdata[72], \cddip2_out_ia_rdata.f.tdata_hi [8]);
tran (cddip2_out_ia_rdata[71], \cddip2_out_ia_rdata.r.part2 [7]);
tran (cddip2_out_ia_rdata[71], \cddip2_out_ia_rdata.f.tdata_hi [7]);
tran (cddip2_out_ia_rdata[70], \cddip2_out_ia_rdata.r.part2 [6]);
tran (cddip2_out_ia_rdata[70], \cddip2_out_ia_rdata.f.tdata_hi [6]);
tran (cddip2_out_ia_rdata[69], \cddip2_out_ia_rdata.r.part2 [5]);
tran (cddip2_out_ia_rdata[69], \cddip2_out_ia_rdata.f.tdata_hi [5]);
tran (cddip2_out_ia_rdata[68], \cddip2_out_ia_rdata.r.part2 [4]);
tran (cddip2_out_ia_rdata[68], \cddip2_out_ia_rdata.f.tdata_hi [4]);
tran (cddip2_out_ia_rdata[67], \cddip2_out_ia_rdata.r.part2 [3]);
tran (cddip2_out_ia_rdata[67], \cddip2_out_ia_rdata.f.tdata_hi [3]);
tran (cddip2_out_ia_rdata[66], \cddip2_out_ia_rdata.r.part2 [2]);
tran (cddip2_out_ia_rdata[66], \cddip2_out_ia_rdata.f.tdata_hi [2]);
tran (cddip2_out_ia_rdata[65], \cddip2_out_ia_rdata.r.part2 [1]);
tran (cddip2_out_ia_rdata[65], \cddip2_out_ia_rdata.f.tdata_hi [1]);
tran (cddip2_out_ia_rdata[64], \cddip2_out_ia_rdata.r.part2 [0]);
tran (cddip2_out_ia_rdata[64], \cddip2_out_ia_rdata.f.tdata_hi [0]);
tran (cddip2_out_ia_rdata[63], \cddip2_out_ia_rdata.r.part1 [31]);
tran (cddip2_out_ia_rdata[63], \cddip2_out_ia_rdata.f.tdata_lo [31]);
tran (cddip2_out_ia_rdata[62], \cddip2_out_ia_rdata.r.part1 [30]);
tran (cddip2_out_ia_rdata[62], \cddip2_out_ia_rdata.f.tdata_lo [30]);
tran (cddip2_out_ia_rdata[61], \cddip2_out_ia_rdata.r.part1 [29]);
tran (cddip2_out_ia_rdata[61], \cddip2_out_ia_rdata.f.tdata_lo [29]);
tran (cddip2_out_ia_rdata[60], \cddip2_out_ia_rdata.r.part1 [28]);
tran (cddip2_out_ia_rdata[60], \cddip2_out_ia_rdata.f.tdata_lo [28]);
tran (cddip2_out_ia_rdata[59], \cddip2_out_ia_rdata.r.part1 [27]);
tran (cddip2_out_ia_rdata[59], \cddip2_out_ia_rdata.f.tdata_lo [27]);
tran (cddip2_out_ia_rdata[58], \cddip2_out_ia_rdata.r.part1 [26]);
tran (cddip2_out_ia_rdata[58], \cddip2_out_ia_rdata.f.tdata_lo [26]);
tran (cddip2_out_ia_rdata[57], \cddip2_out_ia_rdata.r.part1 [25]);
tran (cddip2_out_ia_rdata[57], \cddip2_out_ia_rdata.f.tdata_lo [25]);
tran (cddip2_out_ia_rdata[56], \cddip2_out_ia_rdata.r.part1 [24]);
tran (cddip2_out_ia_rdata[56], \cddip2_out_ia_rdata.f.tdata_lo [24]);
tran (cddip2_out_ia_rdata[55], \cddip2_out_ia_rdata.r.part1 [23]);
tran (cddip2_out_ia_rdata[55], \cddip2_out_ia_rdata.f.tdata_lo [23]);
tran (cddip2_out_ia_rdata[54], \cddip2_out_ia_rdata.r.part1 [22]);
tran (cddip2_out_ia_rdata[54], \cddip2_out_ia_rdata.f.tdata_lo [22]);
tran (cddip2_out_ia_rdata[53], \cddip2_out_ia_rdata.r.part1 [21]);
tran (cddip2_out_ia_rdata[53], \cddip2_out_ia_rdata.f.tdata_lo [21]);
tran (cddip2_out_ia_rdata[52], \cddip2_out_ia_rdata.r.part1 [20]);
tran (cddip2_out_ia_rdata[52], \cddip2_out_ia_rdata.f.tdata_lo [20]);
tran (cddip2_out_ia_rdata[51], \cddip2_out_ia_rdata.r.part1 [19]);
tran (cddip2_out_ia_rdata[51], \cddip2_out_ia_rdata.f.tdata_lo [19]);
tran (cddip2_out_ia_rdata[50], \cddip2_out_ia_rdata.r.part1 [18]);
tran (cddip2_out_ia_rdata[50], \cddip2_out_ia_rdata.f.tdata_lo [18]);
tran (cddip2_out_ia_rdata[49], \cddip2_out_ia_rdata.r.part1 [17]);
tran (cddip2_out_ia_rdata[49], \cddip2_out_ia_rdata.f.tdata_lo [17]);
tran (cddip2_out_ia_rdata[48], \cddip2_out_ia_rdata.r.part1 [16]);
tran (cddip2_out_ia_rdata[48], \cddip2_out_ia_rdata.f.tdata_lo [16]);
tran (cddip2_out_ia_rdata[47], \cddip2_out_ia_rdata.r.part1 [15]);
tran (cddip2_out_ia_rdata[47], \cddip2_out_ia_rdata.f.tdata_lo [15]);
tran (cddip2_out_ia_rdata[46], \cddip2_out_ia_rdata.r.part1 [14]);
tran (cddip2_out_ia_rdata[46], \cddip2_out_ia_rdata.f.tdata_lo [14]);
tran (cddip2_out_ia_rdata[45], \cddip2_out_ia_rdata.r.part1 [13]);
tran (cddip2_out_ia_rdata[45], \cddip2_out_ia_rdata.f.tdata_lo [13]);
tran (cddip2_out_ia_rdata[44], \cddip2_out_ia_rdata.r.part1 [12]);
tran (cddip2_out_ia_rdata[44], \cddip2_out_ia_rdata.f.tdata_lo [12]);
tran (cddip2_out_ia_rdata[43], \cddip2_out_ia_rdata.r.part1 [11]);
tran (cddip2_out_ia_rdata[43], \cddip2_out_ia_rdata.f.tdata_lo [11]);
tran (cddip2_out_ia_rdata[42], \cddip2_out_ia_rdata.r.part1 [10]);
tran (cddip2_out_ia_rdata[42], \cddip2_out_ia_rdata.f.tdata_lo [10]);
tran (cddip2_out_ia_rdata[41], \cddip2_out_ia_rdata.r.part1 [9]);
tran (cddip2_out_ia_rdata[41], \cddip2_out_ia_rdata.f.tdata_lo [9]);
tran (cddip2_out_ia_rdata[40], \cddip2_out_ia_rdata.r.part1 [8]);
tran (cddip2_out_ia_rdata[40], \cddip2_out_ia_rdata.f.tdata_lo [8]);
tran (cddip2_out_ia_rdata[39], \cddip2_out_ia_rdata.r.part1 [7]);
tran (cddip2_out_ia_rdata[39], \cddip2_out_ia_rdata.f.tdata_lo [7]);
tran (cddip2_out_ia_rdata[38], \cddip2_out_ia_rdata.r.part1 [6]);
tran (cddip2_out_ia_rdata[38], \cddip2_out_ia_rdata.f.tdata_lo [6]);
tran (cddip2_out_ia_rdata[37], \cddip2_out_ia_rdata.r.part1 [5]);
tran (cddip2_out_ia_rdata[37], \cddip2_out_ia_rdata.f.tdata_lo [5]);
tran (cddip2_out_ia_rdata[36], \cddip2_out_ia_rdata.r.part1 [4]);
tran (cddip2_out_ia_rdata[36], \cddip2_out_ia_rdata.f.tdata_lo [4]);
tran (cddip2_out_ia_rdata[35], \cddip2_out_ia_rdata.r.part1 [3]);
tran (cddip2_out_ia_rdata[35], \cddip2_out_ia_rdata.f.tdata_lo [3]);
tran (cddip2_out_ia_rdata[34], \cddip2_out_ia_rdata.r.part1 [2]);
tran (cddip2_out_ia_rdata[34], \cddip2_out_ia_rdata.f.tdata_lo [2]);
tran (cddip2_out_ia_rdata[33], \cddip2_out_ia_rdata.r.part1 [1]);
tran (cddip2_out_ia_rdata[33], \cddip2_out_ia_rdata.f.tdata_lo [1]);
tran (cddip2_out_ia_rdata[32], \cddip2_out_ia_rdata.r.part1 [0]);
tran (cddip2_out_ia_rdata[32], \cddip2_out_ia_rdata.f.tdata_lo [0]);
tran (cddip2_out_ia_rdata[31], \cddip2_out_ia_rdata.r.part0 [31]);
tran (cddip2_out_ia_rdata[31], \cddip2_out_ia_rdata.f.eob );
tran (cddip2_out_ia_rdata[30], \cddip2_out_ia_rdata.r.part0 [30]);
tran (cddip2_out_ia_rdata[30], \cddip2_out_ia_rdata.f.bytes_vld [7]);
tran (cddip2_out_ia_rdata[29], \cddip2_out_ia_rdata.r.part0 [29]);
tran (cddip2_out_ia_rdata[29], \cddip2_out_ia_rdata.f.bytes_vld [6]);
tran (cddip2_out_ia_rdata[28], \cddip2_out_ia_rdata.r.part0 [28]);
tran (cddip2_out_ia_rdata[28], \cddip2_out_ia_rdata.f.bytes_vld [5]);
tran (cddip2_out_ia_rdata[27], \cddip2_out_ia_rdata.r.part0 [27]);
tran (cddip2_out_ia_rdata[27], \cddip2_out_ia_rdata.f.bytes_vld [4]);
tran (cddip2_out_ia_rdata[26], \cddip2_out_ia_rdata.r.part0 [26]);
tran (cddip2_out_ia_rdata[26], \cddip2_out_ia_rdata.f.bytes_vld [3]);
tran (cddip2_out_ia_rdata[25], \cddip2_out_ia_rdata.r.part0 [25]);
tran (cddip2_out_ia_rdata[25], \cddip2_out_ia_rdata.f.bytes_vld [2]);
tran (cddip2_out_ia_rdata[24], \cddip2_out_ia_rdata.r.part0 [24]);
tran (cddip2_out_ia_rdata[24], \cddip2_out_ia_rdata.f.bytes_vld [1]);
tran (cddip2_out_ia_rdata[23], \cddip2_out_ia_rdata.r.part0 [23]);
tran (cddip2_out_ia_rdata[23], \cddip2_out_ia_rdata.f.bytes_vld [0]);
tran (cddip2_out_ia_rdata[22], \cddip2_out_ia_rdata.r.part0 [22]);
tran (cddip2_out_ia_rdata[22], \cddip2_out_ia_rdata.f.unused1 [7]);
tran (cddip2_out_ia_rdata[21], \cddip2_out_ia_rdata.r.part0 [21]);
tran (cddip2_out_ia_rdata[21], \cddip2_out_ia_rdata.f.unused1 [6]);
tran (cddip2_out_ia_rdata[20], \cddip2_out_ia_rdata.r.part0 [20]);
tran (cddip2_out_ia_rdata[20], \cddip2_out_ia_rdata.f.unused1 [5]);
tran (cddip2_out_ia_rdata[19], \cddip2_out_ia_rdata.r.part0 [19]);
tran (cddip2_out_ia_rdata[19], \cddip2_out_ia_rdata.f.unused1 [4]);
tran (cddip2_out_ia_rdata[18], \cddip2_out_ia_rdata.r.part0 [18]);
tran (cddip2_out_ia_rdata[18], \cddip2_out_ia_rdata.f.unused1 [3]);
tran (cddip2_out_ia_rdata[17], \cddip2_out_ia_rdata.r.part0 [17]);
tran (cddip2_out_ia_rdata[17], \cddip2_out_ia_rdata.f.unused1 [2]);
tran (cddip2_out_ia_rdata[16], \cddip2_out_ia_rdata.r.part0 [16]);
tran (cddip2_out_ia_rdata[16], \cddip2_out_ia_rdata.f.unused1 [1]);
tran (cddip2_out_ia_rdata[15], \cddip2_out_ia_rdata.r.part0 [15]);
tran (cddip2_out_ia_rdata[15], \cddip2_out_ia_rdata.f.unused1 [0]);
tran (cddip2_out_ia_rdata[14], \cddip2_out_ia_rdata.r.part0 [14]);
tran (cddip2_out_ia_rdata[14], \cddip2_out_ia_rdata.f.tid );
tran (cddip2_out_ia_rdata[13], \cddip2_out_ia_rdata.r.part0 [13]);
tran (cddip2_out_ia_rdata[13], \cddip2_out_ia_rdata.f.tuser [7]);
tran (cddip2_out_ia_rdata[12], \cddip2_out_ia_rdata.r.part0 [12]);
tran (cddip2_out_ia_rdata[12], \cddip2_out_ia_rdata.f.tuser [6]);
tran (cddip2_out_ia_rdata[11], \cddip2_out_ia_rdata.r.part0 [11]);
tran (cddip2_out_ia_rdata[11], \cddip2_out_ia_rdata.f.tuser [5]);
tran (cddip2_out_ia_rdata[10], \cddip2_out_ia_rdata.r.part0 [10]);
tran (cddip2_out_ia_rdata[10], \cddip2_out_ia_rdata.f.tuser [4]);
tran (cddip2_out_ia_rdata[9], \cddip2_out_ia_rdata.r.part0 [9]);
tran (cddip2_out_ia_rdata[9], \cddip2_out_ia_rdata.f.tuser [3]);
tran (cddip2_out_ia_rdata[8], \cddip2_out_ia_rdata.r.part0 [8]);
tran (cddip2_out_ia_rdata[8], \cddip2_out_ia_rdata.f.tuser [2]);
tran (cddip2_out_ia_rdata[7], \cddip2_out_ia_rdata.r.part0 [7]);
tran (cddip2_out_ia_rdata[7], \cddip2_out_ia_rdata.f.tuser [1]);
tran (cddip2_out_ia_rdata[6], \cddip2_out_ia_rdata.r.part0 [6]);
tran (cddip2_out_ia_rdata[6], \cddip2_out_ia_rdata.f.tuser [0]);
tran (cddip2_out_ia_rdata[5], \cddip2_out_ia_rdata.r.part0 [5]);
tran (cddip2_out_ia_rdata[5], \cddip2_out_ia_rdata.f.unused0 [5]);
tran (cddip2_out_ia_rdata[4], \cddip2_out_ia_rdata.r.part0 [4]);
tran (cddip2_out_ia_rdata[4], \cddip2_out_ia_rdata.f.unused0 [4]);
tran (cddip2_out_ia_rdata[3], \cddip2_out_ia_rdata.r.part0 [3]);
tran (cddip2_out_ia_rdata[3], \cddip2_out_ia_rdata.f.unused0 [3]);
tran (cddip2_out_ia_rdata[2], \cddip2_out_ia_rdata.r.part0 [2]);
tran (cddip2_out_ia_rdata[2], \cddip2_out_ia_rdata.f.unused0 [2]);
tran (cddip2_out_ia_rdata[1], \cddip2_out_ia_rdata.r.part0 [1]);
tran (cddip2_out_ia_rdata[1], \cddip2_out_ia_rdata.f.unused0 [1]);
tran (cddip2_out_ia_rdata[0], \cddip2_out_ia_rdata.r.part0 [0]);
tran (cddip2_out_ia_rdata[0], \cddip2_out_ia_rdata.f.unused0 [0]);
tran (cddip2_out_im_status[11], \cddip2_out_im_status.r.part0 [11]);
tran (cddip2_out_im_status[11], \cddip2_out_im_status.f.bank_hi );
tran (cddip2_out_im_status[10], \cddip2_out_im_status.r.part0 [10]);
tran (cddip2_out_im_status[10], \cddip2_out_im_status.f.bank_lo );
tran (cddip2_out_im_status[9], \cddip2_out_im_status.r.part0 [9]);
tran (cddip2_out_im_status[9], \cddip2_out_im_status.f.overflow );
tran (cddip2_out_im_status[8], \cddip2_out_im_status.r.part0 [8]);
tran (cddip2_out_im_status[8], \cddip2_out_im_status.f.wr_pointer [8]);
tran (cddip2_out_im_status[7], \cddip2_out_im_status.r.part0 [7]);
tran (cddip2_out_im_status[7], \cddip2_out_im_status.f.wr_pointer [7]);
tran (cddip2_out_im_status[6], \cddip2_out_im_status.r.part0 [6]);
tran (cddip2_out_im_status[6], \cddip2_out_im_status.f.wr_pointer [6]);
tran (cddip2_out_im_status[5], \cddip2_out_im_status.r.part0 [5]);
tran (cddip2_out_im_status[5], \cddip2_out_im_status.f.wr_pointer [5]);
tran (cddip2_out_im_status[4], \cddip2_out_im_status.r.part0 [4]);
tran (cddip2_out_im_status[4], \cddip2_out_im_status.f.wr_pointer [4]);
tran (cddip2_out_im_status[3], \cddip2_out_im_status.r.part0 [3]);
tran (cddip2_out_im_status[3], \cddip2_out_im_status.f.wr_pointer [3]);
tran (cddip2_out_im_status[2], \cddip2_out_im_status.r.part0 [2]);
tran (cddip2_out_im_status[2], \cddip2_out_im_status.f.wr_pointer [2]);
tran (cddip2_out_im_status[1], \cddip2_out_im_status.r.part0 [1]);
tran (cddip2_out_im_status[1], \cddip2_out_im_status.f.wr_pointer [1]);
tran (cddip2_out_im_status[0], \cddip2_out_im_status.r.part0 [0]);
tran (cddip2_out_im_status[0], \cddip2_out_im_status.f.wr_pointer [0]);
tran (cddip3_out_ia_status[16], \cddip3_out_ia_status.r.part0 [16]);
tran (cddip3_out_ia_status[16], \cddip3_out_ia_status.f.code [2]);
tran (cddip3_out_ia_status[15], \cddip3_out_ia_status.r.part0 [15]);
tran (cddip3_out_ia_status[15], \cddip3_out_ia_status.f.code [1]);
tran (cddip3_out_ia_status[14], \cddip3_out_ia_status.r.part0 [14]);
tran (cddip3_out_ia_status[14], \cddip3_out_ia_status.f.code [0]);
tran (cddip3_out_ia_status[13], \cddip3_out_ia_status.r.part0 [13]);
tran (cddip3_out_ia_status[13], \cddip3_out_ia_status.f.datawords [4]);
tran (cddip3_out_ia_status[12], \cddip3_out_ia_status.r.part0 [12]);
tran (cddip3_out_ia_status[12], \cddip3_out_ia_status.f.datawords [3]);
tran (cddip3_out_ia_status[11], \cddip3_out_ia_status.r.part0 [11]);
tran (cddip3_out_ia_status[11], \cddip3_out_ia_status.f.datawords [2]);
tran (cddip3_out_ia_status[10], \cddip3_out_ia_status.r.part0 [10]);
tran (cddip3_out_ia_status[10], \cddip3_out_ia_status.f.datawords [1]);
tran (cddip3_out_ia_status[9], \cddip3_out_ia_status.r.part0 [9]);
tran (cddip3_out_ia_status[9], \cddip3_out_ia_status.f.datawords [0]);
tran (cddip3_out_ia_status[8], \cddip3_out_ia_status.r.part0 [8]);
tran (cddip3_out_ia_status[8], \cddip3_out_ia_status.f.addr [8]);
tran (cddip3_out_ia_status[7], \cddip3_out_ia_status.r.part0 [7]);
tran (cddip3_out_ia_status[7], \cddip3_out_ia_status.f.addr [7]);
tran (cddip3_out_ia_status[6], \cddip3_out_ia_status.r.part0 [6]);
tran (cddip3_out_ia_status[6], \cddip3_out_ia_status.f.addr [6]);
tran (cddip3_out_ia_status[5], \cddip3_out_ia_status.r.part0 [5]);
tran (cddip3_out_ia_status[5], \cddip3_out_ia_status.f.addr [5]);
tran (cddip3_out_ia_status[4], \cddip3_out_ia_status.r.part0 [4]);
tran (cddip3_out_ia_status[4], \cddip3_out_ia_status.f.addr [4]);
tran (cddip3_out_ia_status[3], \cddip3_out_ia_status.r.part0 [3]);
tran (cddip3_out_ia_status[3], \cddip3_out_ia_status.f.addr [3]);
tran (cddip3_out_ia_status[2], \cddip3_out_ia_status.r.part0 [2]);
tran (cddip3_out_ia_status[2], \cddip3_out_ia_status.f.addr [2]);
tran (cddip3_out_ia_status[1], \cddip3_out_ia_status.r.part0 [1]);
tran (cddip3_out_ia_status[1], \cddip3_out_ia_status.f.addr [1]);
tran (cddip3_out_ia_status[0], \cddip3_out_ia_status.r.part0 [0]);
tran (cddip3_out_ia_status[0], \cddip3_out_ia_status.f.addr [0]);
tran (cddip3_out_ia_capability[15], \cddip3_out_ia_capability.r.part0 [15]);
tran (cddip3_out_ia_capability[15], \cddip3_out_ia_capability.f.ack_error );
tran (cddip3_out_ia_capability[14], \cddip3_out_ia_capability.r.part0 [14]);
tran (cddip3_out_ia_capability[14], \cddip3_out_ia_capability.f.sim_tmo );
tran (cddip3_out_ia_capability[13], \cddip3_out_ia_capability.r.part0 [13]);
tran (cddip3_out_ia_capability[13], \cddip3_out_ia_capability.f.reserved_op [3]);
tran (cddip3_out_ia_capability[12], \cddip3_out_ia_capability.r.part0 [12]);
tran (cddip3_out_ia_capability[12], \cddip3_out_ia_capability.f.reserved_op [2]);
tran (cddip3_out_ia_capability[11], \cddip3_out_ia_capability.r.part0 [11]);
tran (cddip3_out_ia_capability[11], \cddip3_out_ia_capability.f.reserved_op [1]);
tran (cddip3_out_ia_capability[10], \cddip3_out_ia_capability.r.part0 [10]);
tran (cddip3_out_ia_capability[10], \cddip3_out_ia_capability.f.reserved_op [0]);
tran (cddip3_out_ia_capability[9], \cddip3_out_ia_capability.r.part0 [9]);
tran (cddip3_out_ia_capability[9], \cddip3_out_ia_capability.f.compare );
tran (cddip3_out_ia_capability[8], \cddip3_out_ia_capability.r.part0 [8]);
tran (cddip3_out_ia_capability[8], \cddip3_out_ia_capability.f.set_init_start );
tran (cddip3_out_ia_capability[7], \cddip3_out_ia_capability.r.part0 [7]);
tran (cddip3_out_ia_capability[7], \cddip3_out_ia_capability.f.initialize_inc );
tran (cddip3_out_ia_capability[6], \cddip3_out_ia_capability.r.part0 [6]);
tran (cddip3_out_ia_capability[6], \cddip3_out_ia_capability.f.initialize );
tran (cddip3_out_ia_capability[5], \cddip3_out_ia_capability.r.part0 [5]);
tran (cddip3_out_ia_capability[5], \cddip3_out_ia_capability.f.reset );
tran (cddip3_out_ia_capability[4], \cddip3_out_ia_capability.r.part0 [4]);
tran (cddip3_out_ia_capability[4], \cddip3_out_ia_capability.f.disabled );
tran (cddip3_out_ia_capability[3], \cddip3_out_ia_capability.r.part0 [3]);
tran (cddip3_out_ia_capability[3], \cddip3_out_ia_capability.f.enable );
tran (cddip3_out_ia_capability[2], \cddip3_out_ia_capability.r.part0 [2]);
tran (cddip3_out_ia_capability[2], \cddip3_out_ia_capability.f.write );
tran (cddip3_out_ia_capability[1], \cddip3_out_ia_capability.r.part0 [1]);
tran (cddip3_out_ia_capability[1], \cddip3_out_ia_capability.f.read );
tran (cddip3_out_ia_capability[0], \cddip3_out_ia_capability.r.part0 [0]);
tran (cddip3_out_ia_capability[0], \cddip3_out_ia_capability.f.nop );
tran (cddip3_out_ia_capability[19], \cddip3_out_ia_capability.r.part0 [19]);
tran (cddip3_out_ia_capability[19], \cddip3_out_ia_capability.f.mem_type [3]);
tran (cddip3_out_ia_capability[18], \cddip3_out_ia_capability.r.part0 [18]);
tran (cddip3_out_ia_capability[18], \cddip3_out_ia_capability.f.mem_type [2]);
tran (cddip3_out_ia_capability[17], \cddip3_out_ia_capability.r.part0 [17]);
tran (cddip3_out_ia_capability[17], \cddip3_out_ia_capability.f.mem_type [1]);
tran (cddip3_out_ia_capability[16], \cddip3_out_ia_capability.r.part0 [16]);
tran (cddip3_out_ia_capability[16], \cddip3_out_ia_capability.f.mem_type [0]);
tran (cddip3_out_ia_rdata[95], \cddip3_out_ia_rdata.r.part2 [31]);
tran (cddip3_out_ia_rdata[95], \cddip3_out_ia_rdata.f.tdata_hi [31]);
tran (cddip3_out_ia_rdata[94], \cddip3_out_ia_rdata.r.part2 [30]);
tran (cddip3_out_ia_rdata[94], \cddip3_out_ia_rdata.f.tdata_hi [30]);
tran (cddip3_out_ia_rdata[93], \cddip3_out_ia_rdata.r.part2 [29]);
tran (cddip3_out_ia_rdata[93], \cddip3_out_ia_rdata.f.tdata_hi [29]);
tran (cddip3_out_ia_rdata[92], \cddip3_out_ia_rdata.r.part2 [28]);
tran (cddip3_out_ia_rdata[92], \cddip3_out_ia_rdata.f.tdata_hi [28]);
tran (cddip3_out_ia_rdata[91], \cddip3_out_ia_rdata.r.part2 [27]);
tran (cddip3_out_ia_rdata[91], \cddip3_out_ia_rdata.f.tdata_hi [27]);
tran (cddip3_out_ia_rdata[90], \cddip3_out_ia_rdata.r.part2 [26]);
tran (cddip3_out_ia_rdata[90], \cddip3_out_ia_rdata.f.tdata_hi [26]);
tran (cddip3_out_ia_rdata[89], \cddip3_out_ia_rdata.r.part2 [25]);
tran (cddip3_out_ia_rdata[89], \cddip3_out_ia_rdata.f.tdata_hi [25]);
tran (cddip3_out_ia_rdata[88], \cddip3_out_ia_rdata.r.part2 [24]);
tran (cddip3_out_ia_rdata[88], \cddip3_out_ia_rdata.f.tdata_hi [24]);
tran (cddip3_out_ia_rdata[87], \cddip3_out_ia_rdata.r.part2 [23]);
tran (cddip3_out_ia_rdata[87], \cddip3_out_ia_rdata.f.tdata_hi [23]);
tran (cddip3_out_ia_rdata[86], \cddip3_out_ia_rdata.r.part2 [22]);
tran (cddip3_out_ia_rdata[86], \cddip3_out_ia_rdata.f.tdata_hi [22]);
tran (cddip3_out_ia_rdata[85], \cddip3_out_ia_rdata.r.part2 [21]);
tran (cddip3_out_ia_rdata[85], \cddip3_out_ia_rdata.f.tdata_hi [21]);
tran (cddip3_out_ia_rdata[84], \cddip3_out_ia_rdata.r.part2 [20]);
tran (cddip3_out_ia_rdata[84], \cddip3_out_ia_rdata.f.tdata_hi [20]);
tran (cddip3_out_ia_rdata[83], \cddip3_out_ia_rdata.r.part2 [19]);
tran (cddip3_out_ia_rdata[83], \cddip3_out_ia_rdata.f.tdata_hi [19]);
tran (cddip3_out_ia_rdata[82], \cddip3_out_ia_rdata.r.part2 [18]);
tran (cddip3_out_ia_rdata[82], \cddip3_out_ia_rdata.f.tdata_hi [18]);
tran (cddip3_out_ia_rdata[81], \cddip3_out_ia_rdata.r.part2 [17]);
tran (cddip3_out_ia_rdata[81], \cddip3_out_ia_rdata.f.tdata_hi [17]);
tran (cddip3_out_ia_rdata[80], \cddip3_out_ia_rdata.r.part2 [16]);
tran (cddip3_out_ia_rdata[80], \cddip3_out_ia_rdata.f.tdata_hi [16]);
tran (cddip3_out_ia_rdata[79], \cddip3_out_ia_rdata.r.part2 [15]);
tran (cddip3_out_ia_rdata[79], \cddip3_out_ia_rdata.f.tdata_hi [15]);
tran (cddip3_out_ia_rdata[78], \cddip3_out_ia_rdata.r.part2 [14]);
tran (cddip3_out_ia_rdata[78], \cddip3_out_ia_rdata.f.tdata_hi [14]);
tran (cddip3_out_ia_rdata[77], \cddip3_out_ia_rdata.r.part2 [13]);
tran (cddip3_out_ia_rdata[77], \cddip3_out_ia_rdata.f.tdata_hi [13]);
tran (cddip3_out_ia_rdata[76], \cddip3_out_ia_rdata.r.part2 [12]);
tran (cddip3_out_ia_rdata[76], \cddip3_out_ia_rdata.f.tdata_hi [12]);
tran (cddip3_out_ia_rdata[75], \cddip3_out_ia_rdata.r.part2 [11]);
tran (cddip3_out_ia_rdata[75], \cddip3_out_ia_rdata.f.tdata_hi [11]);
tran (cddip3_out_ia_rdata[74], \cddip3_out_ia_rdata.r.part2 [10]);
tran (cddip3_out_ia_rdata[74], \cddip3_out_ia_rdata.f.tdata_hi [10]);
tran (cddip3_out_ia_rdata[73], \cddip3_out_ia_rdata.r.part2 [9]);
tran (cddip3_out_ia_rdata[73], \cddip3_out_ia_rdata.f.tdata_hi [9]);
tran (cddip3_out_ia_rdata[72], \cddip3_out_ia_rdata.r.part2 [8]);
tran (cddip3_out_ia_rdata[72], \cddip3_out_ia_rdata.f.tdata_hi [8]);
tran (cddip3_out_ia_rdata[71], \cddip3_out_ia_rdata.r.part2 [7]);
tran (cddip3_out_ia_rdata[71], \cddip3_out_ia_rdata.f.tdata_hi [7]);
tran (cddip3_out_ia_rdata[70], \cddip3_out_ia_rdata.r.part2 [6]);
tran (cddip3_out_ia_rdata[70], \cddip3_out_ia_rdata.f.tdata_hi [6]);
tran (cddip3_out_ia_rdata[69], \cddip3_out_ia_rdata.r.part2 [5]);
tran (cddip3_out_ia_rdata[69], \cddip3_out_ia_rdata.f.tdata_hi [5]);
tran (cddip3_out_ia_rdata[68], \cddip3_out_ia_rdata.r.part2 [4]);
tran (cddip3_out_ia_rdata[68], \cddip3_out_ia_rdata.f.tdata_hi [4]);
tran (cddip3_out_ia_rdata[67], \cddip3_out_ia_rdata.r.part2 [3]);
tran (cddip3_out_ia_rdata[67], \cddip3_out_ia_rdata.f.tdata_hi [3]);
tran (cddip3_out_ia_rdata[66], \cddip3_out_ia_rdata.r.part2 [2]);
tran (cddip3_out_ia_rdata[66], \cddip3_out_ia_rdata.f.tdata_hi [2]);
tran (cddip3_out_ia_rdata[65], \cddip3_out_ia_rdata.r.part2 [1]);
tran (cddip3_out_ia_rdata[65], \cddip3_out_ia_rdata.f.tdata_hi [1]);
tran (cddip3_out_ia_rdata[64], \cddip3_out_ia_rdata.r.part2 [0]);
tran (cddip3_out_ia_rdata[64], \cddip3_out_ia_rdata.f.tdata_hi [0]);
tran (cddip3_out_ia_rdata[63], \cddip3_out_ia_rdata.r.part1 [31]);
tran (cddip3_out_ia_rdata[63], \cddip3_out_ia_rdata.f.tdata_lo [31]);
tran (cddip3_out_ia_rdata[62], \cddip3_out_ia_rdata.r.part1 [30]);
tran (cddip3_out_ia_rdata[62], \cddip3_out_ia_rdata.f.tdata_lo [30]);
tran (cddip3_out_ia_rdata[61], \cddip3_out_ia_rdata.r.part1 [29]);
tran (cddip3_out_ia_rdata[61], \cddip3_out_ia_rdata.f.tdata_lo [29]);
tran (cddip3_out_ia_rdata[60], \cddip3_out_ia_rdata.r.part1 [28]);
tran (cddip3_out_ia_rdata[60], \cddip3_out_ia_rdata.f.tdata_lo [28]);
tran (cddip3_out_ia_rdata[59], \cddip3_out_ia_rdata.r.part1 [27]);
tran (cddip3_out_ia_rdata[59], \cddip3_out_ia_rdata.f.tdata_lo [27]);
tran (cddip3_out_ia_rdata[58], \cddip3_out_ia_rdata.r.part1 [26]);
tran (cddip3_out_ia_rdata[58], \cddip3_out_ia_rdata.f.tdata_lo [26]);
tran (cddip3_out_ia_rdata[57], \cddip3_out_ia_rdata.r.part1 [25]);
tran (cddip3_out_ia_rdata[57], \cddip3_out_ia_rdata.f.tdata_lo [25]);
tran (cddip3_out_ia_rdata[56], \cddip3_out_ia_rdata.r.part1 [24]);
tran (cddip3_out_ia_rdata[56], \cddip3_out_ia_rdata.f.tdata_lo [24]);
tran (cddip3_out_ia_rdata[55], \cddip3_out_ia_rdata.r.part1 [23]);
tran (cddip3_out_ia_rdata[55], \cddip3_out_ia_rdata.f.tdata_lo [23]);
tran (cddip3_out_ia_rdata[54], \cddip3_out_ia_rdata.r.part1 [22]);
tran (cddip3_out_ia_rdata[54], \cddip3_out_ia_rdata.f.tdata_lo [22]);
tran (cddip3_out_ia_rdata[53], \cddip3_out_ia_rdata.r.part1 [21]);
tran (cddip3_out_ia_rdata[53], \cddip3_out_ia_rdata.f.tdata_lo [21]);
tran (cddip3_out_ia_rdata[52], \cddip3_out_ia_rdata.r.part1 [20]);
tran (cddip3_out_ia_rdata[52], \cddip3_out_ia_rdata.f.tdata_lo [20]);
tran (cddip3_out_ia_rdata[51], \cddip3_out_ia_rdata.r.part1 [19]);
tran (cddip3_out_ia_rdata[51], \cddip3_out_ia_rdata.f.tdata_lo [19]);
tran (cddip3_out_ia_rdata[50], \cddip3_out_ia_rdata.r.part1 [18]);
tran (cddip3_out_ia_rdata[50], \cddip3_out_ia_rdata.f.tdata_lo [18]);
tran (cddip3_out_ia_rdata[49], \cddip3_out_ia_rdata.r.part1 [17]);
tran (cddip3_out_ia_rdata[49], \cddip3_out_ia_rdata.f.tdata_lo [17]);
tran (cddip3_out_ia_rdata[48], \cddip3_out_ia_rdata.r.part1 [16]);
tran (cddip3_out_ia_rdata[48], \cddip3_out_ia_rdata.f.tdata_lo [16]);
tran (cddip3_out_ia_rdata[47], \cddip3_out_ia_rdata.r.part1 [15]);
tran (cddip3_out_ia_rdata[47], \cddip3_out_ia_rdata.f.tdata_lo [15]);
tran (cddip3_out_ia_rdata[46], \cddip3_out_ia_rdata.r.part1 [14]);
tran (cddip3_out_ia_rdata[46], \cddip3_out_ia_rdata.f.tdata_lo [14]);
tran (cddip3_out_ia_rdata[45], \cddip3_out_ia_rdata.r.part1 [13]);
tran (cddip3_out_ia_rdata[45], \cddip3_out_ia_rdata.f.tdata_lo [13]);
tran (cddip3_out_ia_rdata[44], \cddip3_out_ia_rdata.r.part1 [12]);
tran (cddip3_out_ia_rdata[44], \cddip3_out_ia_rdata.f.tdata_lo [12]);
tran (cddip3_out_ia_rdata[43], \cddip3_out_ia_rdata.r.part1 [11]);
tran (cddip3_out_ia_rdata[43], \cddip3_out_ia_rdata.f.tdata_lo [11]);
tran (cddip3_out_ia_rdata[42], \cddip3_out_ia_rdata.r.part1 [10]);
tran (cddip3_out_ia_rdata[42], \cddip3_out_ia_rdata.f.tdata_lo [10]);
tran (cddip3_out_ia_rdata[41], \cddip3_out_ia_rdata.r.part1 [9]);
tran (cddip3_out_ia_rdata[41], \cddip3_out_ia_rdata.f.tdata_lo [9]);
tran (cddip3_out_ia_rdata[40], \cddip3_out_ia_rdata.r.part1 [8]);
tran (cddip3_out_ia_rdata[40], \cddip3_out_ia_rdata.f.tdata_lo [8]);
tran (cddip3_out_ia_rdata[39], \cddip3_out_ia_rdata.r.part1 [7]);
tran (cddip3_out_ia_rdata[39], \cddip3_out_ia_rdata.f.tdata_lo [7]);
tran (cddip3_out_ia_rdata[38], \cddip3_out_ia_rdata.r.part1 [6]);
tran (cddip3_out_ia_rdata[38], \cddip3_out_ia_rdata.f.tdata_lo [6]);
tran (cddip3_out_ia_rdata[37], \cddip3_out_ia_rdata.r.part1 [5]);
tran (cddip3_out_ia_rdata[37], \cddip3_out_ia_rdata.f.tdata_lo [5]);
tran (cddip3_out_ia_rdata[36], \cddip3_out_ia_rdata.r.part1 [4]);
tran (cddip3_out_ia_rdata[36], \cddip3_out_ia_rdata.f.tdata_lo [4]);
tran (cddip3_out_ia_rdata[35], \cddip3_out_ia_rdata.r.part1 [3]);
tran (cddip3_out_ia_rdata[35], \cddip3_out_ia_rdata.f.tdata_lo [3]);
tran (cddip3_out_ia_rdata[34], \cddip3_out_ia_rdata.r.part1 [2]);
tran (cddip3_out_ia_rdata[34], \cddip3_out_ia_rdata.f.tdata_lo [2]);
tran (cddip3_out_ia_rdata[33], \cddip3_out_ia_rdata.r.part1 [1]);
tran (cddip3_out_ia_rdata[33], \cddip3_out_ia_rdata.f.tdata_lo [1]);
tran (cddip3_out_ia_rdata[32], \cddip3_out_ia_rdata.r.part1 [0]);
tran (cddip3_out_ia_rdata[32], \cddip3_out_ia_rdata.f.tdata_lo [0]);
tran (cddip3_out_ia_rdata[31], \cddip3_out_ia_rdata.r.part0 [31]);
tran (cddip3_out_ia_rdata[31], \cddip3_out_ia_rdata.f.eob );
tran (cddip3_out_ia_rdata[30], \cddip3_out_ia_rdata.r.part0 [30]);
tran (cddip3_out_ia_rdata[30], \cddip3_out_ia_rdata.f.bytes_vld [7]);
tran (cddip3_out_ia_rdata[29], \cddip3_out_ia_rdata.r.part0 [29]);
tran (cddip3_out_ia_rdata[29], \cddip3_out_ia_rdata.f.bytes_vld [6]);
tran (cddip3_out_ia_rdata[28], \cddip3_out_ia_rdata.r.part0 [28]);
tran (cddip3_out_ia_rdata[28], \cddip3_out_ia_rdata.f.bytes_vld [5]);
tran (cddip3_out_ia_rdata[27], \cddip3_out_ia_rdata.r.part0 [27]);
tran (cddip3_out_ia_rdata[27], \cddip3_out_ia_rdata.f.bytes_vld [4]);
tran (cddip3_out_ia_rdata[26], \cddip3_out_ia_rdata.r.part0 [26]);
tran (cddip3_out_ia_rdata[26], \cddip3_out_ia_rdata.f.bytes_vld [3]);
tran (cddip3_out_ia_rdata[25], \cddip3_out_ia_rdata.r.part0 [25]);
tran (cddip3_out_ia_rdata[25], \cddip3_out_ia_rdata.f.bytes_vld [2]);
tran (cddip3_out_ia_rdata[24], \cddip3_out_ia_rdata.r.part0 [24]);
tran (cddip3_out_ia_rdata[24], \cddip3_out_ia_rdata.f.bytes_vld [1]);
tran (cddip3_out_ia_rdata[23], \cddip3_out_ia_rdata.r.part0 [23]);
tran (cddip3_out_ia_rdata[23], \cddip3_out_ia_rdata.f.bytes_vld [0]);
tran (cddip3_out_ia_rdata[22], \cddip3_out_ia_rdata.r.part0 [22]);
tran (cddip3_out_ia_rdata[22], \cddip3_out_ia_rdata.f.unused1 [7]);
tran (cddip3_out_ia_rdata[21], \cddip3_out_ia_rdata.r.part0 [21]);
tran (cddip3_out_ia_rdata[21], \cddip3_out_ia_rdata.f.unused1 [6]);
tran (cddip3_out_ia_rdata[20], \cddip3_out_ia_rdata.r.part0 [20]);
tran (cddip3_out_ia_rdata[20], \cddip3_out_ia_rdata.f.unused1 [5]);
tran (cddip3_out_ia_rdata[19], \cddip3_out_ia_rdata.r.part0 [19]);
tran (cddip3_out_ia_rdata[19], \cddip3_out_ia_rdata.f.unused1 [4]);
tran (cddip3_out_ia_rdata[18], \cddip3_out_ia_rdata.r.part0 [18]);
tran (cddip3_out_ia_rdata[18], \cddip3_out_ia_rdata.f.unused1 [3]);
tran (cddip3_out_ia_rdata[17], \cddip3_out_ia_rdata.r.part0 [17]);
tran (cddip3_out_ia_rdata[17], \cddip3_out_ia_rdata.f.unused1 [2]);
tran (cddip3_out_ia_rdata[16], \cddip3_out_ia_rdata.r.part0 [16]);
tran (cddip3_out_ia_rdata[16], \cddip3_out_ia_rdata.f.unused1 [1]);
tran (cddip3_out_ia_rdata[15], \cddip3_out_ia_rdata.r.part0 [15]);
tran (cddip3_out_ia_rdata[15], \cddip3_out_ia_rdata.f.unused1 [0]);
tran (cddip3_out_ia_rdata[14], \cddip3_out_ia_rdata.r.part0 [14]);
tran (cddip3_out_ia_rdata[14], \cddip3_out_ia_rdata.f.tid );
tran (cddip3_out_ia_rdata[13], \cddip3_out_ia_rdata.r.part0 [13]);
tran (cddip3_out_ia_rdata[13], \cddip3_out_ia_rdata.f.tuser [7]);
tran (cddip3_out_ia_rdata[12], \cddip3_out_ia_rdata.r.part0 [12]);
tran (cddip3_out_ia_rdata[12], \cddip3_out_ia_rdata.f.tuser [6]);
tran (cddip3_out_ia_rdata[11], \cddip3_out_ia_rdata.r.part0 [11]);
tran (cddip3_out_ia_rdata[11], \cddip3_out_ia_rdata.f.tuser [5]);
tran (cddip3_out_ia_rdata[10], \cddip3_out_ia_rdata.r.part0 [10]);
tran (cddip3_out_ia_rdata[10], \cddip3_out_ia_rdata.f.tuser [4]);
tran (cddip3_out_ia_rdata[9], \cddip3_out_ia_rdata.r.part0 [9]);
tran (cddip3_out_ia_rdata[9], \cddip3_out_ia_rdata.f.tuser [3]);
tran (cddip3_out_ia_rdata[8], \cddip3_out_ia_rdata.r.part0 [8]);
tran (cddip3_out_ia_rdata[8], \cddip3_out_ia_rdata.f.tuser [2]);
tran (cddip3_out_ia_rdata[7], \cddip3_out_ia_rdata.r.part0 [7]);
tran (cddip3_out_ia_rdata[7], \cddip3_out_ia_rdata.f.tuser [1]);
tran (cddip3_out_ia_rdata[6], \cddip3_out_ia_rdata.r.part0 [6]);
tran (cddip3_out_ia_rdata[6], \cddip3_out_ia_rdata.f.tuser [0]);
tran (cddip3_out_ia_rdata[5], \cddip3_out_ia_rdata.r.part0 [5]);
tran (cddip3_out_ia_rdata[5], \cddip3_out_ia_rdata.f.unused0 [5]);
tran (cddip3_out_ia_rdata[4], \cddip3_out_ia_rdata.r.part0 [4]);
tran (cddip3_out_ia_rdata[4], \cddip3_out_ia_rdata.f.unused0 [4]);
tran (cddip3_out_ia_rdata[3], \cddip3_out_ia_rdata.r.part0 [3]);
tran (cddip3_out_ia_rdata[3], \cddip3_out_ia_rdata.f.unused0 [3]);
tran (cddip3_out_ia_rdata[2], \cddip3_out_ia_rdata.r.part0 [2]);
tran (cddip3_out_ia_rdata[2], \cddip3_out_ia_rdata.f.unused0 [2]);
tran (cddip3_out_ia_rdata[1], \cddip3_out_ia_rdata.r.part0 [1]);
tran (cddip3_out_ia_rdata[1], \cddip3_out_ia_rdata.f.unused0 [1]);
tran (cddip3_out_ia_rdata[0], \cddip3_out_ia_rdata.r.part0 [0]);
tran (cddip3_out_ia_rdata[0], \cddip3_out_ia_rdata.f.unused0 [0]);
tran (cddip3_out_im_status[11], \cddip3_out_im_status.r.part0 [11]);
tran (cddip3_out_im_status[11], \cddip3_out_im_status.f.bank_hi );
tran (cddip3_out_im_status[10], \cddip3_out_im_status.r.part0 [10]);
tran (cddip3_out_im_status[10], \cddip3_out_im_status.f.bank_lo );
tran (cddip3_out_im_status[9], \cddip3_out_im_status.r.part0 [9]);
tran (cddip3_out_im_status[9], \cddip3_out_im_status.f.overflow );
tran (cddip3_out_im_status[8], \cddip3_out_im_status.r.part0 [8]);
tran (cddip3_out_im_status[8], \cddip3_out_im_status.f.wr_pointer [8]);
tran (cddip3_out_im_status[7], \cddip3_out_im_status.r.part0 [7]);
tran (cddip3_out_im_status[7], \cddip3_out_im_status.f.wr_pointer [7]);
tran (cddip3_out_im_status[6], \cddip3_out_im_status.r.part0 [6]);
tran (cddip3_out_im_status[6], \cddip3_out_im_status.f.wr_pointer [6]);
tran (cddip3_out_im_status[5], \cddip3_out_im_status.r.part0 [5]);
tran (cddip3_out_im_status[5], \cddip3_out_im_status.f.wr_pointer [5]);
tran (cddip3_out_im_status[4], \cddip3_out_im_status.r.part0 [4]);
tran (cddip3_out_im_status[4], \cddip3_out_im_status.f.wr_pointer [4]);
tran (cddip3_out_im_status[3], \cddip3_out_im_status.r.part0 [3]);
tran (cddip3_out_im_status[3], \cddip3_out_im_status.f.wr_pointer [3]);
tran (cddip3_out_im_status[2], \cddip3_out_im_status.r.part0 [2]);
tran (cddip3_out_im_status[2], \cddip3_out_im_status.f.wr_pointer [2]);
tran (cddip3_out_im_status[1], \cddip3_out_im_status.r.part0 [1]);
tran (cddip3_out_im_status[1], \cddip3_out_im_status.f.wr_pointer [1]);
tran (cddip3_out_im_status[0], \cddip3_out_im_status.r.part0 [0]);
tran (cddip3_out_im_status[0], \cddip3_out_im_status.f.wr_pointer [0]);
tran (ckv_ia_capability[19], \ckv_ia_capability.r.part0 [19]);
tran (ckv_ia_capability[19], \ckv_ia_capability.f.mem_type [3]);
tran (ckv_ia_capability[18], \ckv_ia_capability.r.part0 [18]);
tran (ckv_ia_capability[18], \ckv_ia_capability.f.mem_type [2]);
tran (ckv_ia_capability[17], \ckv_ia_capability.r.part0 [17]);
tran (ckv_ia_capability[17], \ckv_ia_capability.f.mem_type [1]);
tran (ckv_ia_capability[16], \ckv_ia_capability.r.part0 [16]);
tran (ckv_ia_capability[16], \ckv_ia_capability.f.mem_type [0]);
tran (ckv_ia_capability[15], \ckv_ia_capability.r.part0 [15]);
tran (ckv_ia_capability[15], \ckv_ia_capability.f.ack_error );
tran (ckv_ia_capability[14], \ckv_ia_capability.r.part0 [14]);
tran (ckv_ia_capability[14], \ckv_ia_capability.f.sim_tmo );
tran (ckv_ia_capability[13], \ckv_ia_capability.r.part0 [13]);
tran (ckv_ia_capability[13], \ckv_ia_capability.f.reserved_op [3]);
tran (ckv_ia_capability[12], \ckv_ia_capability.r.part0 [12]);
tran (ckv_ia_capability[12], \ckv_ia_capability.f.reserved_op [2]);
tran (ckv_ia_capability[11], \ckv_ia_capability.r.part0 [11]);
tran (ckv_ia_capability[11], \ckv_ia_capability.f.reserved_op [1]);
tran (ckv_ia_capability[10], \ckv_ia_capability.r.part0 [10]);
tran (ckv_ia_capability[10], \ckv_ia_capability.f.reserved_op [0]);
tran (ckv_ia_capability[9], \ckv_ia_capability.r.part0 [9]);
tran (ckv_ia_capability[9], \ckv_ia_capability.f.compare );
tran (ckv_ia_capability[8], \ckv_ia_capability.r.part0 [8]);
tran (ckv_ia_capability[8], \ckv_ia_capability.f.set_init_start );
tran (ckv_ia_capability[7], \ckv_ia_capability.r.part0 [7]);
tran (ckv_ia_capability[7], \ckv_ia_capability.f.initialize_inc );
tran (ckv_ia_capability[6], \ckv_ia_capability.r.part0 [6]);
tran (ckv_ia_capability[6], \ckv_ia_capability.f.initialize );
tran (ckv_ia_capability[5], \ckv_ia_capability.r.part0 [5]);
tran (ckv_ia_capability[5], \ckv_ia_capability.f.reset );
tran (ckv_ia_capability[4], \ckv_ia_capability.r.part0 [4]);
tran (ckv_ia_capability[4], \ckv_ia_capability.f.disabled );
tran (ckv_ia_capability[3], \ckv_ia_capability.r.part0 [3]);
tran (ckv_ia_capability[3], \ckv_ia_capability.f.enable );
tran (ckv_ia_capability[2], \ckv_ia_capability.r.part0 [2]);
tran (ckv_ia_capability[2], \ckv_ia_capability.f.write );
tran (ckv_ia_capability[1], \ckv_ia_capability.r.part0 [1]);
tran (ckv_ia_capability[1], \ckv_ia_capability.f.read );
tran (ckv_ia_capability[0], \ckv_ia_capability.r.part0 [0]);
tran (ckv_ia_capability[0], \ckv_ia_capability.f.nop );
tran (ckv_ia_status[22], \ckv_ia_status.r.part0 [22]);
tran (ckv_ia_status[22], \ckv_ia_status.f.code [2]);
tran (ckv_ia_status[21], \ckv_ia_status.r.part0 [21]);
tran (ckv_ia_status[21], \ckv_ia_status.f.code [1]);
tran (ckv_ia_status[20], \ckv_ia_status.r.part0 [20]);
tran (ckv_ia_status[20], \ckv_ia_status.f.code [0]);
tran (ckv_ia_status[19], \ckv_ia_status.r.part0 [19]);
tran (ckv_ia_status[19], \ckv_ia_status.f.datawords [4]);
tran (ckv_ia_status[18], \ckv_ia_status.r.part0 [18]);
tran (ckv_ia_status[18], \ckv_ia_status.f.datawords [3]);
tran (ckv_ia_status[17], \ckv_ia_status.r.part0 [17]);
tran (ckv_ia_status[17], \ckv_ia_status.f.datawords [2]);
tran (ckv_ia_status[16], \ckv_ia_status.r.part0 [16]);
tran (ckv_ia_status[16], \ckv_ia_status.f.datawords [1]);
tran (ckv_ia_status[15], \ckv_ia_status.r.part0 [15]);
tran (ckv_ia_status[15], \ckv_ia_status.f.datawords [0]);
tran (ckv_ia_status[14], \ckv_ia_status.r.part0 [14]);
tran (ckv_ia_status[14], \ckv_ia_status.f.addr [14]);
tran (ckv_ia_status[13], \ckv_ia_status.r.part0 [13]);
tran (ckv_ia_status[13], \ckv_ia_status.f.addr [13]);
tran (ckv_ia_status[12], \ckv_ia_status.r.part0 [12]);
tran (ckv_ia_status[12], \ckv_ia_status.f.addr [12]);
tran (ckv_ia_status[11], \ckv_ia_status.r.part0 [11]);
tran (ckv_ia_status[11], \ckv_ia_status.f.addr [11]);
tran (ckv_ia_status[10], \ckv_ia_status.r.part0 [10]);
tran (ckv_ia_status[10], \ckv_ia_status.f.addr [10]);
tran (ckv_ia_status[9], \ckv_ia_status.r.part0 [9]);
tran (ckv_ia_status[9], \ckv_ia_status.f.addr [9]);
tran (ckv_ia_status[8], \ckv_ia_status.r.part0 [8]);
tran (ckv_ia_status[8], \ckv_ia_status.f.addr [8]);
tran (ckv_ia_status[7], \ckv_ia_status.r.part0 [7]);
tran (ckv_ia_status[7], \ckv_ia_status.f.addr [7]);
tran (ckv_ia_status[6], \ckv_ia_status.r.part0 [6]);
tran (ckv_ia_status[6], \ckv_ia_status.f.addr [6]);
tran (ckv_ia_status[5], \ckv_ia_status.r.part0 [5]);
tran (ckv_ia_status[5], \ckv_ia_status.f.addr [5]);
tran (ckv_ia_status[4], \ckv_ia_status.r.part0 [4]);
tran (ckv_ia_status[4], \ckv_ia_status.f.addr [4]);
tran (ckv_ia_status[3], \ckv_ia_status.r.part0 [3]);
tran (ckv_ia_status[3], \ckv_ia_status.f.addr [3]);
tran (ckv_ia_status[2], \ckv_ia_status.r.part0 [2]);
tran (ckv_ia_status[2], \ckv_ia_status.f.addr [2]);
tran (ckv_ia_status[1], \ckv_ia_status.r.part0 [1]);
tran (ckv_ia_status[1], \ckv_ia_status.f.addr [1]);
tran (ckv_ia_status[0], \ckv_ia_status.r.part0 [0]);
tran (ckv_ia_status[0], \ckv_ia_status.f.addr [0]);
tran (kim_ia_capability[19], \kim_ia_capability.r.part0 [19]);
tran (kim_ia_capability[19], \kim_ia_capability.f.mem_type [3]);
tran (kim_ia_capability[18], \kim_ia_capability.r.part0 [18]);
tran (kim_ia_capability[18], \kim_ia_capability.f.mem_type [2]);
tran (kim_ia_capability[17], \kim_ia_capability.r.part0 [17]);
tran (kim_ia_capability[17], \kim_ia_capability.f.mem_type [1]);
tran (kim_ia_capability[16], \kim_ia_capability.r.part0 [16]);
tran (kim_ia_capability[16], \kim_ia_capability.f.mem_type [0]);
tran (kim_ia_capability[15], \kim_ia_capability.r.part0 [15]);
tran (kim_ia_capability[15], \kim_ia_capability.f.ack_error );
tran (kim_ia_capability[14], \kim_ia_capability.r.part0 [14]);
tran (kim_ia_capability[14], \kim_ia_capability.f.sim_tmo );
tran (kim_ia_capability[13], \kim_ia_capability.r.part0 [13]);
tran (kim_ia_capability[13], \kim_ia_capability.f.reserved_op [3]);
tran (kim_ia_capability[12], \kim_ia_capability.r.part0 [12]);
tran (kim_ia_capability[12], \kim_ia_capability.f.reserved_op [2]);
tran (kim_ia_capability[11], \kim_ia_capability.r.part0 [11]);
tran (kim_ia_capability[11], \kim_ia_capability.f.reserved_op [1]);
tran (kim_ia_capability[10], \kim_ia_capability.r.part0 [10]);
tran (kim_ia_capability[10], \kim_ia_capability.f.reserved_op [0]);
tran (kim_ia_capability[9], \kim_ia_capability.r.part0 [9]);
tran (kim_ia_capability[9], \kim_ia_capability.f.compare );
tran (kim_ia_capability[8], \kim_ia_capability.r.part0 [8]);
tran (kim_ia_capability[8], \kim_ia_capability.f.set_init_start );
tran (kim_ia_capability[7], \kim_ia_capability.r.part0 [7]);
tran (kim_ia_capability[7], \kim_ia_capability.f.initialize_inc );
tran (kim_ia_capability[6], \kim_ia_capability.r.part0 [6]);
tran (kim_ia_capability[6], \kim_ia_capability.f.initialize );
tran (kim_ia_capability[5], \kim_ia_capability.r.part0 [5]);
tran (kim_ia_capability[5], \kim_ia_capability.f.reset );
tran (kim_ia_capability[4], \kim_ia_capability.r.part0 [4]);
tran (kim_ia_capability[4], \kim_ia_capability.f.disabled );
tran (kim_ia_capability[3], \kim_ia_capability.r.part0 [3]);
tran (kim_ia_capability[3], \kim_ia_capability.f.enable );
tran (kim_ia_capability[2], \kim_ia_capability.r.part0 [2]);
tran (kim_ia_capability[2], \kim_ia_capability.f.write );
tran (kim_ia_capability[1], \kim_ia_capability.r.part0 [1]);
tran (kim_ia_capability[1], \kim_ia_capability.f.read );
tran (kim_ia_capability[0], \kim_ia_capability.r.part0 [0]);
tran (kim_ia_capability[0], \kim_ia_capability.f.nop );
tran (kim_ia_status[21], \kim_ia_status.r.part0 [21]);
tran (kim_ia_status[21], \kim_ia_status.f.code [2]);
tran (kim_ia_status[20], \kim_ia_status.r.part0 [20]);
tran (kim_ia_status[20], \kim_ia_status.f.code [1]);
tran (kim_ia_status[19], \kim_ia_status.r.part0 [19]);
tran (kim_ia_status[19], \kim_ia_status.f.code [0]);
tran (kim_ia_status[18], \kim_ia_status.r.part0 [18]);
tran (kim_ia_status[18], \kim_ia_status.f.datawords [4]);
tran (kim_ia_status[17], \kim_ia_status.r.part0 [17]);
tran (kim_ia_status[17], \kim_ia_status.f.datawords [3]);
tran (kim_ia_status[16], \kim_ia_status.r.part0 [16]);
tran (kim_ia_status[16], \kim_ia_status.f.datawords [2]);
tran (kim_ia_status[15], \kim_ia_status.r.part0 [15]);
tran (kim_ia_status[15], \kim_ia_status.f.datawords [1]);
tran (kim_ia_status[14], \kim_ia_status.r.part0 [14]);
tran (kim_ia_status[14], \kim_ia_status.f.datawords [0]);
tran (kim_ia_status[13], \kim_ia_status.r.part0 [13]);
tran (kim_ia_status[13], \kim_ia_status.f.addr [13]);
tran (kim_ia_status[12], \kim_ia_status.r.part0 [12]);
tran (kim_ia_status[12], \kim_ia_status.f.addr [12]);
tran (kim_ia_status[11], \kim_ia_status.r.part0 [11]);
tran (kim_ia_status[11], \kim_ia_status.f.addr [11]);
tran (kim_ia_status[10], \kim_ia_status.r.part0 [10]);
tran (kim_ia_status[10], \kim_ia_status.f.addr [10]);
tran (kim_ia_status[9], \kim_ia_status.r.part0 [9]);
tran (kim_ia_status[9], \kim_ia_status.f.addr [9]);
tran (kim_ia_status[8], \kim_ia_status.r.part0 [8]);
tran (kim_ia_status[8], \kim_ia_status.f.addr [8]);
tran (kim_ia_status[7], \kim_ia_status.r.part0 [7]);
tran (kim_ia_status[7], \kim_ia_status.f.addr [7]);
tran (kim_ia_status[6], \kim_ia_status.r.part0 [6]);
tran (kim_ia_status[6], \kim_ia_status.f.addr [6]);
tran (kim_ia_status[5], \kim_ia_status.r.part0 [5]);
tran (kim_ia_status[5], \kim_ia_status.f.addr [5]);
tran (kim_ia_status[4], \kim_ia_status.r.part0 [4]);
tran (kim_ia_status[4], \kim_ia_status.f.addr [4]);
tran (kim_ia_status[3], \kim_ia_status.r.part0 [3]);
tran (kim_ia_status[3], \kim_ia_status.f.addr [3]);
tran (kim_ia_status[2], \kim_ia_status.r.part0 [2]);
tran (kim_ia_status[2], \kim_ia_status.f.addr [2]);
tran (kim_ia_status[1], \kim_ia_status.r.part0 [1]);
tran (kim_ia_status[1], \kim_ia_status.f.addr [1]);
tran (kim_ia_status[0], \kim_ia_status.r.part0 [0]);
tran (kim_ia_status[0], \kim_ia_status.f.addr [0]);
tran (sa_snapshot_ia_status[12], \sa_snapshot_ia_status.r.part0 [12]);
tran (sa_snapshot_ia_status[12], \sa_snapshot_ia_status.f.code [2]);
tran (sa_snapshot_ia_status[11], \sa_snapshot_ia_status.r.part0 [11]);
tran (sa_snapshot_ia_status[11], \sa_snapshot_ia_status.f.code [1]);
tran (sa_snapshot_ia_status[10], \sa_snapshot_ia_status.r.part0 [10]);
tran (sa_snapshot_ia_status[10], \sa_snapshot_ia_status.f.code [0]);
tran (sa_snapshot_ia_status[9], \sa_snapshot_ia_status.r.part0 [9]);
tran (sa_snapshot_ia_status[9], \sa_snapshot_ia_status.f.datawords [4]);
tran (sa_snapshot_ia_status[8], \sa_snapshot_ia_status.r.part0 [8]);
tran (sa_snapshot_ia_status[8], \sa_snapshot_ia_status.f.datawords [3]);
tran (sa_snapshot_ia_status[7], \sa_snapshot_ia_status.r.part0 [7]);
tran (sa_snapshot_ia_status[7], \sa_snapshot_ia_status.f.datawords [2]);
tran (sa_snapshot_ia_status[6], \sa_snapshot_ia_status.r.part0 [6]);
tran (sa_snapshot_ia_status[6], \sa_snapshot_ia_status.f.datawords [1]);
tran (sa_snapshot_ia_status[5], \sa_snapshot_ia_status.r.part0 [5]);
tran (sa_snapshot_ia_status[5], \sa_snapshot_ia_status.f.datawords [0]);
tran (sa_snapshot_ia_status[4], \sa_snapshot_ia_status.r.part0 [4]);
tran (sa_snapshot_ia_status[4], \sa_snapshot_ia_status.f.addr [4]);
tran (sa_snapshot_ia_status[3], \sa_snapshot_ia_status.r.part0 [3]);
tran (sa_snapshot_ia_status[3], \sa_snapshot_ia_status.f.addr [3]);
tran (sa_snapshot_ia_status[2], \sa_snapshot_ia_status.r.part0 [2]);
tran (sa_snapshot_ia_status[2], \sa_snapshot_ia_status.f.addr [2]);
tran (sa_snapshot_ia_status[1], \sa_snapshot_ia_status.r.part0 [1]);
tran (sa_snapshot_ia_status[1], \sa_snapshot_ia_status.f.addr [1]);
tran (sa_snapshot_ia_status[0], \sa_snapshot_ia_status.r.part0 [0]);
tran (sa_snapshot_ia_status[0], \sa_snapshot_ia_status.f.addr [0]);
tran (sa_snapshot_ia_capability[15], \sa_snapshot_ia_capability.r.part0 [15]);
tran (sa_snapshot_ia_capability[15], \sa_snapshot_ia_capability.f.ack_error );
tran (sa_snapshot_ia_capability[14], \sa_snapshot_ia_capability.r.part0 [14]);
tran (sa_snapshot_ia_capability[14], \sa_snapshot_ia_capability.f.sim_tmo );
tran (sa_snapshot_ia_capability[13], \sa_snapshot_ia_capability.r.part0 [13]);
tran (sa_snapshot_ia_capability[13], \sa_snapshot_ia_capability.f.reserved_op [3]);
tran (sa_snapshot_ia_capability[12], \sa_snapshot_ia_capability.r.part0 [12]);
tran (sa_snapshot_ia_capability[12], \sa_snapshot_ia_capability.f.reserved_op [2]);
tran (sa_snapshot_ia_capability[11], \sa_snapshot_ia_capability.r.part0 [11]);
tran (sa_snapshot_ia_capability[11], \sa_snapshot_ia_capability.f.reserved_op [1]);
tran (sa_snapshot_ia_capability[10], \sa_snapshot_ia_capability.r.part0 [10]);
tran (sa_snapshot_ia_capability[10], \sa_snapshot_ia_capability.f.reserved_op [0]);
tran (sa_snapshot_ia_capability[9], \sa_snapshot_ia_capability.r.part0 [9]);
tran (sa_snapshot_ia_capability[9], \sa_snapshot_ia_capability.f.compare );
tran (sa_snapshot_ia_capability[8], \sa_snapshot_ia_capability.r.part0 [8]);
tran (sa_snapshot_ia_capability[8], \sa_snapshot_ia_capability.f.set_init_start );
tran (sa_snapshot_ia_capability[7], \sa_snapshot_ia_capability.r.part0 [7]);
tran (sa_snapshot_ia_capability[7], \sa_snapshot_ia_capability.f.initialize_inc );
tran (sa_snapshot_ia_capability[6], \sa_snapshot_ia_capability.r.part0 [6]);
tran (sa_snapshot_ia_capability[6], \sa_snapshot_ia_capability.f.initialize );
tran (sa_snapshot_ia_capability[5], \sa_snapshot_ia_capability.r.part0 [5]);
tran (sa_snapshot_ia_capability[5], \sa_snapshot_ia_capability.f.reset );
tran (sa_snapshot_ia_capability[4], \sa_snapshot_ia_capability.r.part0 [4]);
tran (sa_snapshot_ia_capability[4], \sa_snapshot_ia_capability.f.disabled );
tran (sa_snapshot_ia_capability[3], \sa_snapshot_ia_capability.r.part0 [3]);
tran (sa_snapshot_ia_capability[3], \sa_snapshot_ia_capability.f.enable );
tran (sa_snapshot_ia_capability[2], \sa_snapshot_ia_capability.r.part0 [2]);
tran (sa_snapshot_ia_capability[2], \sa_snapshot_ia_capability.f.write );
tran (sa_snapshot_ia_capability[1], \sa_snapshot_ia_capability.r.part0 [1]);
tran (sa_snapshot_ia_capability[1], \sa_snapshot_ia_capability.f.read );
tran (sa_snapshot_ia_capability[0], \sa_snapshot_ia_capability.r.part0 [0]);
tran (sa_snapshot_ia_capability[0], \sa_snapshot_ia_capability.f.nop );
tran (sa_snapshot_ia_capability[19], \sa_snapshot_ia_capability.r.part0 [19]);
tran (sa_snapshot_ia_capability[19], \sa_snapshot_ia_capability.f.mem_type [3]);
tran (sa_snapshot_ia_capability[18], \sa_snapshot_ia_capability.r.part0 [18]);
tran (sa_snapshot_ia_capability[18], \sa_snapshot_ia_capability.f.mem_type [2]);
tran (sa_snapshot_ia_capability[17], \sa_snapshot_ia_capability.r.part0 [17]);
tran (sa_snapshot_ia_capability[17], \sa_snapshot_ia_capability.f.mem_type [1]);
tran (sa_snapshot_ia_capability[16], \sa_snapshot_ia_capability.r.part0 [16]);
tran (sa_snapshot_ia_capability[16], \sa_snapshot_ia_capability.f.mem_type [0]);
tran (sa_snapshot_ia_rdata[63], \sa_snapshot_ia_rdata.r.part1 [31]);
tran (sa_snapshot_ia_rdata[63], \sa_snapshot_ia_rdata.f.unused [13]);
tran (sa_snapshot_ia_rdata[62], \sa_snapshot_ia_rdata.r.part1 [30]);
tran (sa_snapshot_ia_rdata[62], \sa_snapshot_ia_rdata.f.unused [12]);
tran (sa_snapshot_ia_rdata[61], \sa_snapshot_ia_rdata.r.part1 [29]);
tran (sa_snapshot_ia_rdata[61], \sa_snapshot_ia_rdata.f.unused [11]);
tran (sa_snapshot_ia_rdata[60], \sa_snapshot_ia_rdata.r.part1 [28]);
tran (sa_snapshot_ia_rdata[60], \sa_snapshot_ia_rdata.f.unused [10]);
tran (sa_snapshot_ia_rdata[59], \sa_snapshot_ia_rdata.r.part1 [27]);
tran (sa_snapshot_ia_rdata[59], \sa_snapshot_ia_rdata.f.unused [9]);
tran (sa_snapshot_ia_rdata[58], \sa_snapshot_ia_rdata.r.part1 [26]);
tran (sa_snapshot_ia_rdata[58], \sa_snapshot_ia_rdata.f.unused [8]);
tran (sa_snapshot_ia_rdata[57], \sa_snapshot_ia_rdata.r.part1 [25]);
tran (sa_snapshot_ia_rdata[57], \sa_snapshot_ia_rdata.f.unused [7]);
tran (sa_snapshot_ia_rdata[56], \sa_snapshot_ia_rdata.r.part1 [24]);
tran (sa_snapshot_ia_rdata[56], \sa_snapshot_ia_rdata.f.unused [6]);
tran (sa_snapshot_ia_rdata[55], \sa_snapshot_ia_rdata.r.part1 [23]);
tran (sa_snapshot_ia_rdata[55], \sa_snapshot_ia_rdata.f.unused [5]);
tran (sa_snapshot_ia_rdata[54], \sa_snapshot_ia_rdata.r.part1 [22]);
tran (sa_snapshot_ia_rdata[54], \sa_snapshot_ia_rdata.f.unused [4]);
tran (sa_snapshot_ia_rdata[53], \sa_snapshot_ia_rdata.r.part1 [21]);
tran (sa_snapshot_ia_rdata[53], \sa_snapshot_ia_rdata.f.unused [3]);
tran (sa_snapshot_ia_rdata[52], \sa_snapshot_ia_rdata.r.part1 [20]);
tran (sa_snapshot_ia_rdata[52], \sa_snapshot_ia_rdata.f.unused [2]);
tran (sa_snapshot_ia_rdata[51], \sa_snapshot_ia_rdata.r.part1 [19]);
tran (sa_snapshot_ia_rdata[51], \sa_snapshot_ia_rdata.f.unused [1]);
tran (sa_snapshot_ia_rdata[50], \sa_snapshot_ia_rdata.r.part1 [18]);
tran (sa_snapshot_ia_rdata[50], \sa_snapshot_ia_rdata.f.unused [0]);
tran (sa_snapshot_ia_rdata[49], \sa_snapshot_ia_rdata.r.part1 [17]);
tran (sa_snapshot_ia_rdata[49], \sa_snapshot_ia_rdata.f.upper [17]);
tran (sa_snapshot_ia_rdata[48], \sa_snapshot_ia_rdata.r.part1 [16]);
tran (sa_snapshot_ia_rdata[48], \sa_snapshot_ia_rdata.f.upper [16]);
tran (sa_snapshot_ia_rdata[47], \sa_snapshot_ia_rdata.r.part1 [15]);
tran (sa_snapshot_ia_rdata[47], \sa_snapshot_ia_rdata.f.upper [15]);
tran (sa_snapshot_ia_rdata[46], \sa_snapshot_ia_rdata.r.part1 [14]);
tran (sa_snapshot_ia_rdata[46], \sa_snapshot_ia_rdata.f.upper [14]);
tran (sa_snapshot_ia_rdata[45], \sa_snapshot_ia_rdata.r.part1 [13]);
tran (sa_snapshot_ia_rdata[45], \sa_snapshot_ia_rdata.f.upper [13]);
tran (sa_snapshot_ia_rdata[44], \sa_snapshot_ia_rdata.r.part1 [12]);
tran (sa_snapshot_ia_rdata[44], \sa_snapshot_ia_rdata.f.upper [12]);
tran (sa_snapshot_ia_rdata[43], \sa_snapshot_ia_rdata.r.part1 [11]);
tran (sa_snapshot_ia_rdata[43], \sa_snapshot_ia_rdata.f.upper [11]);
tran (sa_snapshot_ia_rdata[42], \sa_snapshot_ia_rdata.r.part1 [10]);
tran (sa_snapshot_ia_rdata[42], \sa_snapshot_ia_rdata.f.upper [10]);
tran (sa_snapshot_ia_rdata[41], \sa_snapshot_ia_rdata.r.part1 [9]);
tran (sa_snapshot_ia_rdata[41], \sa_snapshot_ia_rdata.f.upper [9]);
tran (sa_snapshot_ia_rdata[40], \sa_snapshot_ia_rdata.r.part1 [8]);
tran (sa_snapshot_ia_rdata[40], \sa_snapshot_ia_rdata.f.upper [8]);
tran (sa_snapshot_ia_rdata[39], \sa_snapshot_ia_rdata.r.part1 [7]);
tran (sa_snapshot_ia_rdata[39], \sa_snapshot_ia_rdata.f.upper [7]);
tran (sa_snapshot_ia_rdata[38], \sa_snapshot_ia_rdata.r.part1 [6]);
tran (sa_snapshot_ia_rdata[38], \sa_snapshot_ia_rdata.f.upper [6]);
tran (sa_snapshot_ia_rdata[37], \sa_snapshot_ia_rdata.r.part1 [5]);
tran (sa_snapshot_ia_rdata[37], \sa_snapshot_ia_rdata.f.upper [5]);
tran (sa_snapshot_ia_rdata[36], \sa_snapshot_ia_rdata.r.part1 [4]);
tran (sa_snapshot_ia_rdata[36], \sa_snapshot_ia_rdata.f.upper [4]);
tran (sa_snapshot_ia_rdata[35], \sa_snapshot_ia_rdata.r.part1 [3]);
tran (sa_snapshot_ia_rdata[35], \sa_snapshot_ia_rdata.f.upper [3]);
tran (sa_snapshot_ia_rdata[34], \sa_snapshot_ia_rdata.r.part1 [2]);
tran (sa_snapshot_ia_rdata[34], \sa_snapshot_ia_rdata.f.upper [2]);
tran (sa_snapshot_ia_rdata[33], \sa_snapshot_ia_rdata.r.part1 [1]);
tran (sa_snapshot_ia_rdata[33], \sa_snapshot_ia_rdata.f.upper [1]);
tran (sa_snapshot_ia_rdata[32], \sa_snapshot_ia_rdata.r.part1 [0]);
tran (sa_snapshot_ia_rdata[32], \sa_snapshot_ia_rdata.f.upper [0]);
tran (sa_snapshot_ia_rdata[31], \sa_snapshot_ia_rdata.r.part0 [31]);
tran (sa_snapshot_ia_rdata[31], \sa_snapshot_ia_rdata.f.lower [31]);
tran (sa_snapshot_ia_rdata[30], \sa_snapshot_ia_rdata.r.part0 [30]);
tran (sa_snapshot_ia_rdata[30], \sa_snapshot_ia_rdata.f.lower [30]);
tran (sa_snapshot_ia_rdata[29], \sa_snapshot_ia_rdata.r.part0 [29]);
tran (sa_snapshot_ia_rdata[29], \sa_snapshot_ia_rdata.f.lower [29]);
tran (sa_snapshot_ia_rdata[28], \sa_snapshot_ia_rdata.r.part0 [28]);
tran (sa_snapshot_ia_rdata[28], \sa_snapshot_ia_rdata.f.lower [28]);
tran (sa_snapshot_ia_rdata[27], \sa_snapshot_ia_rdata.r.part0 [27]);
tran (sa_snapshot_ia_rdata[27], \sa_snapshot_ia_rdata.f.lower [27]);
tran (sa_snapshot_ia_rdata[26], \sa_snapshot_ia_rdata.r.part0 [26]);
tran (sa_snapshot_ia_rdata[26], \sa_snapshot_ia_rdata.f.lower [26]);
tran (sa_snapshot_ia_rdata[25], \sa_snapshot_ia_rdata.r.part0 [25]);
tran (sa_snapshot_ia_rdata[25], \sa_snapshot_ia_rdata.f.lower [25]);
tran (sa_snapshot_ia_rdata[24], \sa_snapshot_ia_rdata.r.part0 [24]);
tran (sa_snapshot_ia_rdata[24], \sa_snapshot_ia_rdata.f.lower [24]);
tran (sa_snapshot_ia_rdata[23], \sa_snapshot_ia_rdata.r.part0 [23]);
tran (sa_snapshot_ia_rdata[23], \sa_snapshot_ia_rdata.f.lower [23]);
tran (sa_snapshot_ia_rdata[22], \sa_snapshot_ia_rdata.r.part0 [22]);
tran (sa_snapshot_ia_rdata[22], \sa_snapshot_ia_rdata.f.lower [22]);
tran (sa_snapshot_ia_rdata[21], \sa_snapshot_ia_rdata.r.part0 [21]);
tran (sa_snapshot_ia_rdata[21], \sa_snapshot_ia_rdata.f.lower [21]);
tran (sa_snapshot_ia_rdata[20], \sa_snapshot_ia_rdata.r.part0 [20]);
tran (sa_snapshot_ia_rdata[20], \sa_snapshot_ia_rdata.f.lower [20]);
tran (sa_snapshot_ia_rdata[19], \sa_snapshot_ia_rdata.r.part0 [19]);
tran (sa_snapshot_ia_rdata[19], \sa_snapshot_ia_rdata.f.lower [19]);
tran (sa_snapshot_ia_rdata[18], \sa_snapshot_ia_rdata.r.part0 [18]);
tran (sa_snapshot_ia_rdata[18], \sa_snapshot_ia_rdata.f.lower [18]);
tran (sa_snapshot_ia_rdata[17], \sa_snapshot_ia_rdata.r.part0 [17]);
tran (sa_snapshot_ia_rdata[17], \sa_snapshot_ia_rdata.f.lower [17]);
tran (sa_snapshot_ia_rdata[16], \sa_snapshot_ia_rdata.r.part0 [16]);
tran (sa_snapshot_ia_rdata[16], \sa_snapshot_ia_rdata.f.lower [16]);
tran (sa_snapshot_ia_rdata[15], \sa_snapshot_ia_rdata.r.part0 [15]);
tran (sa_snapshot_ia_rdata[15], \sa_snapshot_ia_rdata.f.lower [15]);
tran (sa_snapshot_ia_rdata[14], \sa_snapshot_ia_rdata.r.part0 [14]);
tran (sa_snapshot_ia_rdata[14], \sa_snapshot_ia_rdata.f.lower [14]);
tran (sa_snapshot_ia_rdata[13], \sa_snapshot_ia_rdata.r.part0 [13]);
tran (sa_snapshot_ia_rdata[13], \sa_snapshot_ia_rdata.f.lower [13]);
tran (sa_snapshot_ia_rdata[12], \sa_snapshot_ia_rdata.r.part0 [12]);
tran (sa_snapshot_ia_rdata[12], \sa_snapshot_ia_rdata.f.lower [12]);
tran (sa_snapshot_ia_rdata[11], \sa_snapshot_ia_rdata.r.part0 [11]);
tran (sa_snapshot_ia_rdata[11], \sa_snapshot_ia_rdata.f.lower [11]);
tran (sa_snapshot_ia_rdata[10], \sa_snapshot_ia_rdata.r.part0 [10]);
tran (sa_snapshot_ia_rdata[10], \sa_snapshot_ia_rdata.f.lower [10]);
tran (sa_snapshot_ia_rdata[9], \sa_snapshot_ia_rdata.r.part0 [9]);
tran (sa_snapshot_ia_rdata[9], \sa_snapshot_ia_rdata.f.lower [9]);
tran (sa_snapshot_ia_rdata[8], \sa_snapshot_ia_rdata.r.part0 [8]);
tran (sa_snapshot_ia_rdata[8], \sa_snapshot_ia_rdata.f.lower [8]);
tran (sa_snapshot_ia_rdata[7], \sa_snapshot_ia_rdata.r.part0 [7]);
tran (sa_snapshot_ia_rdata[7], \sa_snapshot_ia_rdata.f.lower [7]);
tran (sa_snapshot_ia_rdata[6], \sa_snapshot_ia_rdata.r.part0 [6]);
tran (sa_snapshot_ia_rdata[6], \sa_snapshot_ia_rdata.f.lower [6]);
tran (sa_snapshot_ia_rdata[5], \sa_snapshot_ia_rdata.r.part0 [5]);
tran (sa_snapshot_ia_rdata[5], \sa_snapshot_ia_rdata.f.lower [5]);
tran (sa_snapshot_ia_rdata[4], \sa_snapshot_ia_rdata.r.part0 [4]);
tran (sa_snapshot_ia_rdata[4], \sa_snapshot_ia_rdata.f.lower [4]);
tran (sa_snapshot_ia_rdata[3], \sa_snapshot_ia_rdata.r.part0 [3]);
tran (sa_snapshot_ia_rdata[3], \sa_snapshot_ia_rdata.f.lower [3]);
tran (sa_snapshot_ia_rdata[2], \sa_snapshot_ia_rdata.r.part0 [2]);
tran (sa_snapshot_ia_rdata[2], \sa_snapshot_ia_rdata.f.lower [2]);
tran (sa_snapshot_ia_rdata[1], \sa_snapshot_ia_rdata.r.part0 [1]);
tran (sa_snapshot_ia_rdata[1], \sa_snapshot_ia_rdata.f.lower [1]);
tran (sa_snapshot_ia_rdata[0], \sa_snapshot_ia_rdata.r.part0 [0]);
tran (sa_snapshot_ia_rdata[0], \sa_snapshot_ia_rdata.f.lower [0]);
tran (sa_count_ia_status[12], \sa_count_ia_status.r.part0 [12]);
tran (sa_count_ia_status[12], \sa_count_ia_status.f.code [2]);
tran (sa_count_ia_status[11], \sa_count_ia_status.r.part0 [11]);
tran (sa_count_ia_status[11], \sa_count_ia_status.f.code [1]);
tran (sa_count_ia_status[10], \sa_count_ia_status.r.part0 [10]);
tran (sa_count_ia_status[10], \sa_count_ia_status.f.code [0]);
tran (sa_count_ia_status[9], \sa_count_ia_status.r.part0 [9]);
tran (sa_count_ia_status[9], \sa_count_ia_status.f.datawords [4]);
tran (sa_count_ia_status[8], \sa_count_ia_status.r.part0 [8]);
tran (sa_count_ia_status[8], \sa_count_ia_status.f.datawords [3]);
tran (sa_count_ia_status[7], \sa_count_ia_status.r.part0 [7]);
tran (sa_count_ia_status[7], \sa_count_ia_status.f.datawords [2]);
tran (sa_count_ia_status[6], \sa_count_ia_status.r.part0 [6]);
tran (sa_count_ia_status[6], \sa_count_ia_status.f.datawords [1]);
tran (sa_count_ia_status[5], \sa_count_ia_status.r.part0 [5]);
tran (sa_count_ia_status[5], \sa_count_ia_status.f.datawords [0]);
tran (sa_count_ia_status[4], \sa_count_ia_status.r.part0 [4]);
tran (sa_count_ia_status[4], \sa_count_ia_status.f.addr [4]);
tran (sa_count_ia_status[3], \sa_count_ia_status.r.part0 [3]);
tran (sa_count_ia_status[3], \sa_count_ia_status.f.addr [3]);
tran (sa_count_ia_status[2], \sa_count_ia_status.r.part0 [2]);
tran (sa_count_ia_status[2], \sa_count_ia_status.f.addr [2]);
tran (sa_count_ia_status[1], \sa_count_ia_status.r.part0 [1]);
tran (sa_count_ia_status[1], \sa_count_ia_status.f.addr [1]);
tran (sa_count_ia_status[0], \sa_count_ia_status.r.part0 [0]);
tran (sa_count_ia_status[0], \sa_count_ia_status.f.addr [0]);
tran (sa_count_ia_capability[15], \sa_count_ia_capability.r.part0 [15]);
tran (sa_count_ia_capability[15], \sa_count_ia_capability.f.ack_error );
tran (sa_count_ia_capability[14], \sa_count_ia_capability.r.part0 [14]);
tran (sa_count_ia_capability[14], \sa_count_ia_capability.f.sim_tmo );
tran (sa_count_ia_capability[13], \sa_count_ia_capability.r.part0 [13]);
tran (sa_count_ia_capability[13], \sa_count_ia_capability.f.reserved_op [3]);
tran (sa_count_ia_capability[12], \sa_count_ia_capability.r.part0 [12]);
tran (sa_count_ia_capability[12], \sa_count_ia_capability.f.reserved_op [2]);
tran (sa_count_ia_capability[11], \sa_count_ia_capability.r.part0 [11]);
tran (sa_count_ia_capability[11], \sa_count_ia_capability.f.reserved_op [1]);
tran (sa_count_ia_capability[10], \sa_count_ia_capability.r.part0 [10]);
tran (sa_count_ia_capability[10], \sa_count_ia_capability.f.reserved_op [0]);
tran (sa_count_ia_capability[9], \sa_count_ia_capability.r.part0 [9]);
tran (sa_count_ia_capability[9], \sa_count_ia_capability.f.compare );
tran (sa_count_ia_capability[8], \sa_count_ia_capability.r.part0 [8]);
tran (sa_count_ia_capability[8], \sa_count_ia_capability.f.set_init_start );
tran (sa_count_ia_capability[7], \sa_count_ia_capability.r.part0 [7]);
tran (sa_count_ia_capability[7], \sa_count_ia_capability.f.initialize_inc );
tran (sa_count_ia_capability[6], \sa_count_ia_capability.r.part0 [6]);
tran (sa_count_ia_capability[6], \sa_count_ia_capability.f.initialize );
tran (sa_count_ia_capability[5], \sa_count_ia_capability.r.part0 [5]);
tran (sa_count_ia_capability[5], \sa_count_ia_capability.f.reset );
tran (sa_count_ia_capability[4], \sa_count_ia_capability.r.part0 [4]);
tran (sa_count_ia_capability[4], \sa_count_ia_capability.f.disabled );
tran (sa_count_ia_capability[3], \sa_count_ia_capability.r.part0 [3]);
tran (sa_count_ia_capability[3], \sa_count_ia_capability.f.enable );
tran (sa_count_ia_capability[2], \sa_count_ia_capability.r.part0 [2]);
tran (sa_count_ia_capability[2], \sa_count_ia_capability.f.write );
tran (sa_count_ia_capability[1], \sa_count_ia_capability.r.part0 [1]);
tran (sa_count_ia_capability[1], \sa_count_ia_capability.f.read );
tran (sa_count_ia_capability[0], \sa_count_ia_capability.r.part0 [0]);
tran (sa_count_ia_capability[0], \sa_count_ia_capability.f.nop );
tran (sa_count_ia_capability[19], \sa_count_ia_capability.r.part0 [19]);
tran (sa_count_ia_capability[19], \sa_count_ia_capability.f.mem_type [3]);
tran (sa_count_ia_capability[18], \sa_count_ia_capability.r.part0 [18]);
tran (sa_count_ia_capability[18], \sa_count_ia_capability.f.mem_type [2]);
tran (sa_count_ia_capability[17], \sa_count_ia_capability.r.part0 [17]);
tran (sa_count_ia_capability[17], \sa_count_ia_capability.f.mem_type [1]);
tran (sa_count_ia_capability[16], \sa_count_ia_capability.r.part0 [16]);
tran (sa_count_ia_capability[16], \sa_count_ia_capability.f.mem_type [0]);
tran (sa_count_ia_rdata[63], \sa_count_ia_rdata.r.part1 [31]);
tran (sa_count_ia_rdata[63], \sa_count_ia_rdata.f.unused [13]);
tran (sa_count_ia_rdata[62], \sa_count_ia_rdata.r.part1 [30]);
tran (sa_count_ia_rdata[62], \sa_count_ia_rdata.f.unused [12]);
tran (sa_count_ia_rdata[61], \sa_count_ia_rdata.r.part1 [29]);
tran (sa_count_ia_rdata[61], \sa_count_ia_rdata.f.unused [11]);
tran (sa_count_ia_rdata[60], \sa_count_ia_rdata.r.part1 [28]);
tran (sa_count_ia_rdata[60], \sa_count_ia_rdata.f.unused [10]);
tran (sa_count_ia_rdata[59], \sa_count_ia_rdata.r.part1 [27]);
tran (sa_count_ia_rdata[59], \sa_count_ia_rdata.f.unused [9]);
tran (sa_count_ia_rdata[58], \sa_count_ia_rdata.r.part1 [26]);
tran (sa_count_ia_rdata[58], \sa_count_ia_rdata.f.unused [8]);
tran (sa_count_ia_rdata[57], \sa_count_ia_rdata.r.part1 [25]);
tran (sa_count_ia_rdata[57], \sa_count_ia_rdata.f.unused [7]);
tran (sa_count_ia_rdata[56], \sa_count_ia_rdata.r.part1 [24]);
tran (sa_count_ia_rdata[56], \sa_count_ia_rdata.f.unused [6]);
tran (sa_count_ia_rdata[55], \sa_count_ia_rdata.r.part1 [23]);
tran (sa_count_ia_rdata[55], \sa_count_ia_rdata.f.unused [5]);
tran (sa_count_ia_rdata[54], \sa_count_ia_rdata.r.part1 [22]);
tran (sa_count_ia_rdata[54], \sa_count_ia_rdata.f.unused [4]);
tran (sa_count_ia_rdata[53], \sa_count_ia_rdata.r.part1 [21]);
tran (sa_count_ia_rdata[53], \sa_count_ia_rdata.f.unused [3]);
tran (sa_count_ia_rdata[52], \sa_count_ia_rdata.r.part1 [20]);
tran (sa_count_ia_rdata[52], \sa_count_ia_rdata.f.unused [2]);
tran (sa_count_ia_rdata[51], \sa_count_ia_rdata.r.part1 [19]);
tran (sa_count_ia_rdata[51], \sa_count_ia_rdata.f.unused [1]);
tran (sa_count_ia_rdata[50], \sa_count_ia_rdata.r.part1 [18]);
tran (sa_count_ia_rdata[50], \sa_count_ia_rdata.f.unused [0]);
tran (sa_count_ia_rdata[49], \sa_count_ia_rdata.r.part1 [17]);
tran (sa_count_ia_rdata[49], \sa_count_ia_rdata.f.upper [17]);
tran (sa_count_ia_rdata[48], \sa_count_ia_rdata.r.part1 [16]);
tran (sa_count_ia_rdata[48], \sa_count_ia_rdata.f.upper [16]);
tran (sa_count_ia_rdata[47], \sa_count_ia_rdata.r.part1 [15]);
tran (sa_count_ia_rdata[47], \sa_count_ia_rdata.f.upper [15]);
tran (sa_count_ia_rdata[46], \sa_count_ia_rdata.r.part1 [14]);
tran (sa_count_ia_rdata[46], \sa_count_ia_rdata.f.upper [14]);
tran (sa_count_ia_rdata[45], \sa_count_ia_rdata.r.part1 [13]);
tran (sa_count_ia_rdata[45], \sa_count_ia_rdata.f.upper [13]);
tran (sa_count_ia_rdata[44], \sa_count_ia_rdata.r.part1 [12]);
tran (sa_count_ia_rdata[44], \sa_count_ia_rdata.f.upper [12]);
tran (sa_count_ia_rdata[43], \sa_count_ia_rdata.r.part1 [11]);
tran (sa_count_ia_rdata[43], \sa_count_ia_rdata.f.upper [11]);
tran (sa_count_ia_rdata[42], \sa_count_ia_rdata.r.part1 [10]);
tran (sa_count_ia_rdata[42], \sa_count_ia_rdata.f.upper [10]);
tran (sa_count_ia_rdata[41], \sa_count_ia_rdata.r.part1 [9]);
tran (sa_count_ia_rdata[41], \sa_count_ia_rdata.f.upper [9]);
tran (sa_count_ia_rdata[40], \sa_count_ia_rdata.r.part1 [8]);
tran (sa_count_ia_rdata[40], \sa_count_ia_rdata.f.upper [8]);
tran (sa_count_ia_rdata[39], \sa_count_ia_rdata.r.part1 [7]);
tran (sa_count_ia_rdata[39], \sa_count_ia_rdata.f.upper [7]);
tran (sa_count_ia_rdata[38], \sa_count_ia_rdata.r.part1 [6]);
tran (sa_count_ia_rdata[38], \sa_count_ia_rdata.f.upper [6]);
tran (sa_count_ia_rdata[37], \sa_count_ia_rdata.r.part1 [5]);
tran (sa_count_ia_rdata[37], \sa_count_ia_rdata.f.upper [5]);
tran (sa_count_ia_rdata[36], \sa_count_ia_rdata.r.part1 [4]);
tran (sa_count_ia_rdata[36], \sa_count_ia_rdata.f.upper [4]);
tran (sa_count_ia_rdata[35], \sa_count_ia_rdata.r.part1 [3]);
tran (sa_count_ia_rdata[35], \sa_count_ia_rdata.f.upper [3]);
tran (sa_count_ia_rdata[34], \sa_count_ia_rdata.r.part1 [2]);
tran (sa_count_ia_rdata[34], \sa_count_ia_rdata.f.upper [2]);
tran (sa_count_ia_rdata[33], \sa_count_ia_rdata.r.part1 [1]);
tran (sa_count_ia_rdata[33], \sa_count_ia_rdata.f.upper [1]);
tran (sa_count_ia_rdata[32], \sa_count_ia_rdata.r.part1 [0]);
tran (sa_count_ia_rdata[32], \sa_count_ia_rdata.f.upper [0]);
tran (sa_count_ia_rdata[31], \sa_count_ia_rdata.r.part0 [31]);
tran (sa_count_ia_rdata[31], \sa_count_ia_rdata.f.lower [31]);
tran (sa_count_ia_rdata[30], \sa_count_ia_rdata.r.part0 [30]);
tran (sa_count_ia_rdata[30], \sa_count_ia_rdata.f.lower [30]);
tran (sa_count_ia_rdata[29], \sa_count_ia_rdata.r.part0 [29]);
tran (sa_count_ia_rdata[29], \sa_count_ia_rdata.f.lower [29]);
tran (sa_count_ia_rdata[28], \sa_count_ia_rdata.r.part0 [28]);
tran (sa_count_ia_rdata[28], \sa_count_ia_rdata.f.lower [28]);
tran (sa_count_ia_rdata[27], \sa_count_ia_rdata.r.part0 [27]);
tran (sa_count_ia_rdata[27], \sa_count_ia_rdata.f.lower [27]);
tran (sa_count_ia_rdata[26], \sa_count_ia_rdata.r.part0 [26]);
tran (sa_count_ia_rdata[26], \sa_count_ia_rdata.f.lower [26]);
tran (sa_count_ia_rdata[25], \sa_count_ia_rdata.r.part0 [25]);
tran (sa_count_ia_rdata[25], \sa_count_ia_rdata.f.lower [25]);
tran (sa_count_ia_rdata[24], \sa_count_ia_rdata.r.part0 [24]);
tran (sa_count_ia_rdata[24], \sa_count_ia_rdata.f.lower [24]);
tran (sa_count_ia_rdata[23], \sa_count_ia_rdata.r.part0 [23]);
tran (sa_count_ia_rdata[23], \sa_count_ia_rdata.f.lower [23]);
tran (sa_count_ia_rdata[22], \sa_count_ia_rdata.r.part0 [22]);
tran (sa_count_ia_rdata[22], \sa_count_ia_rdata.f.lower [22]);
tran (sa_count_ia_rdata[21], \sa_count_ia_rdata.r.part0 [21]);
tran (sa_count_ia_rdata[21], \sa_count_ia_rdata.f.lower [21]);
tran (sa_count_ia_rdata[20], \sa_count_ia_rdata.r.part0 [20]);
tran (sa_count_ia_rdata[20], \sa_count_ia_rdata.f.lower [20]);
tran (sa_count_ia_rdata[19], \sa_count_ia_rdata.r.part0 [19]);
tran (sa_count_ia_rdata[19], \sa_count_ia_rdata.f.lower [19]);
tran (sa_count_ia_rdata[18], \sa_count_ia_rdata.r.part0 [18]);
tran (sa_count_ia_rdata[18], \sa_count_ia_rdata.f.lower [18]);
tran (sa_count_ia_rdata[17], \sa_count_ia_rdata.r.part0 [17]);
tran (sa_count_ia_rdata[17], \sa_count_ia_rdata.f.lower [17]);
tran (sa_count_ia_rdata[16], \sa_count_ia_rdata.r.part0 [16]);
tran (sa_count_ia_rdata[16], \sa_count_ia_rdata.f.lower [16]);
tran (sa_count_ia_rdata[15], \sa_count_ia_rdata.r.part0 [15]);
tran (sa_count_ia_rdata[15], \sa_count_ia_rdata.f.lower [15]);
tran (sa_count_ia_rdata[14], \sa_count_ia_rdata.r.part0 [14]);
tran (sa_count_ia_rdata[14], \sa_count_ia_rdata.f.lower [14]);
tran (sa_count_ia_rdata[13], \sa_count_ia_rdata.r.part0 [13]);
tran (sa_count_ia_rdata[13], \sa_count_ia_rdata.f.lower [13]);
tran (sa_count_ia_rdata[12], \sa_count_ia_rdata.r.part0 [12]);
tran (sa_count_ia_rdata[12], \sa_count_ia_rdata.f.lower [12]);
tran (sa_count_ia_rdata[11], \sa_count_ia_rdata.r.part0 [11]);
tran (sa_count_ia_rdata[11], \sa_count_ia_rdata.f.lower [11]);
tran (sa_count_ia_rdata[10], \sa_count_ia_rdata.r.part0 [10]);
tran (sa_count_ia_rdata[10], \sa_count_ia_rdata.f.lower [10]);
tran (sa_count_ia_rdata[9], \sa_count_ia_rdata.r.part0 [9]);
tran (sa_count_ia_rdata[9], \sa_count_ia_rdata.f.lower [9]);
tran (sa_count_ia_rdata[8], \sa_count_ia_rdata.r.part0 [8]);
tran (sa_count_ia_rdata[8], \sa_count_ia_rdata.f.lower [8]);
tran (sa_count_ia_rdata[7], \sa_count_ia_rdata.r.part0 [7]);
tran (sa_count_ia_rdata[7], \sa_count_ia_rdata.f.lower [7]);
tran (sa_count_ia_rdata[6], \sa_count_ia_rdata.r.part0 [6]);
tran (sa_count_ia_rdata[6], \sa_count_ia_rdata.f.lower [6]);
tran (sa_count_ia_rdata[5], \sa_count_ia_rdata.r.part0 [5]);
tran (sa_count_ia_rdata[5], \sa_count_ia_rdata.f.lower [5]);
tran (sa_count_ia_rdata[4], \sa_count_ia_rdata.r.part0 [4]);
tran (sa_count_ia_rdata[4], \sa_count_ia_rdata.f.lower [4]);
tran (sa_count_ia_rdata[3], \sa_count_ia_rdata.r.part0 [3]);
tran (sa_count_ia_rdata[3], \sa_count_ia_rdata.f.lower [3]);
tran (sa_count_ia_rdata[2], \sa_count_ia_rdata.r.part0 [2]);
tran (sa_count_ia_rdata[2], \sa_count_ia_rdata.f.lower [2]);
tran (sa_count_ia_rdata[1], \sa_count_ia_rdata.r.part0 [1]);
tran (sa_count_ia_rdata[1], \sa_count_ia_rdata.f.lower [1]);
tran (sa_count_ia_rdata[0], \sa_count_ia_rdata.r.part0 [0]);
tran (sa_count_ia_rdata[0], \sa_count_ia_rdata.f.lower [0]);
tran (sa_ctrl_ia_status[12], \sa_ctrl_ia_status.r.part0 [12]);
tran (sa_ctrl_ia_status[12], \sa_ctrl_ia_status.f.code [2]);
tran (sa_ctrl_ia_status[11], \sa_ctrl_ia_status.r.part0 [11]);
tran (sa_ctrl_ia_status[11], \sa_ctrl_ia_status.f.code [1]);
tran (sa_ctrl_ia_status[10], \sa_ctrl_ia_status.r.part0 [10]);
tran (sa_ctrl_ia_status[10], \sa_ctrl_ia_status.f.code [0]);
tran (sa_ctrl_ia_status[9], \sa_ctrl_ia_status.r.part0 [9]);
tran (sa_ctrl_ia_status[9], \sa_ctrl_ia_status.f.datawords [4]);
tran (sa_ctrl_ia_status[8], \sa_ctrl_ia_status.r.part0 [8]);
tran (sa_ctrl_ia_status[8], \sa_ctrl_ia_status.f.datawords [3]);
tran (sa_ctrl_ia_status[7], \sa_ctrl_ia_status.r.part0 [7]);
tran (sa_ctrl_ia_status[7], \sa_ctrl_ia_status.f.datawords [2]);
tran (sa_ctrl_ia_status[6], \sa_ctrl_ia_status.r.part0 [6]);
tran (sa_ctrl_ia_status[6], \sa_ctrl_ia_status.f.datawords [1]);
tran (sa_ctrl_ia_status[5], \sa_ctrl_ia_status.r.part0 [5]);
tran (sa_ctrl_ia_status[5], \sa_ctrl_ia_status.f.datawords [0]);
tran (sa_ctrl_ia_status[4], \sa_ctrl_ia_status.r.part0 [4]);
tran (sa_ctrl_ia_status[4], \sa_ctrl_ia_status.f.addr [4]);
tran (sa_ctrl_ia_status[3], \sa_ctrl_ia_status.r.part0 [3]);
tran (sa_ctrl_ia_status[3], \sa_ctrl_ia_status.f.addr [3]);
tran (sa_ctrl_ia_status[2], \sa_ctrl_ia_status.r.part0 [2]);
tran (sa_ctrl_ia_status[2], \sa_ctrl_ia_status.f.addr [2]);
tran (sa_ctrl_ia_status[1], \sa_ctrl_ia_status.r.part0 [1]);
tran (sa_ctrl_ia_status[1], \sa_ctrl_ia_status.f.addr [1]);
tran (sa_ctrl_ia_status[0], \sa_ctrl_ia_status.r.part0 [0]);
tran (sa_ctrl_ia_status[0], \sa_ctrl_ia_status.f.addr [0]);
tran (sa_ctrl_ia_capability[15], \sa_ctrl_ia_capability.r.part0 [15]);
tran (sa_ctrl_ia_capability[15], \sa_ctrl_ia_capability.f.ack_error );
tran (sa_ctrl_ia_capability[14], \sa_ctrl_ia_capability.r.part0 [14]);
tran (sa_ctrl_ia_capability[14], \sa_ctrl_ia_capability.f.sim_tmo );
tran (sa_ctrl_ia_capability[13], \sa_ctrl_ia_capability.r.part0 [13]);
tran (sa_ctrl_ia_capability[13], \sa_ctrl_ia_capability.f.reserved_op [3]);
tran (sa_ctrl_ia_capability[12], \sa_ctrl_ia_capability.r.part0 [12]);
tran (sa_ctrl_ia_capability[12], \sa_ctrl_ia_capability.f.reserved_op [2]);
tran (sa_ctrl_ia_capability[11], \sa_ctrl_ia_capability.r.part0 [11]);
tran (sa_ctrl_ia_capability[11], \sa_ctrl_ia_capability.f.reserved_op [1]);
tran (sa_ctrl_ia_capability[10], \sa_ctrl_ia_capability.r.part0 [10]);
tran (sa_ctrl_ia_capability[10], \sa_ctrl_ia_capability.f.reserved_op [0]);
tran (sa_ctrl_ia_capability[9], \sa_ctrl_ia_capability.r.part0 [9]);
tran (sa_ctrl_ia_capability[9], \sa_ctrl_ia_capability.f.compare );
tran (sa_ctrl_ia_capability[8], \sa_ctrl_ia_capability.r.part0 [8]);
tran (sa_ctrl_ia_capability[8], \sa_ctrl_ia_capability.f.set_init_start );
tran (sa_ctrl_ia_capability[7], \sa_ctrl_ia_capability.r.part0 [7]);
tran (sa_ctrl_ia_capability[7], \sa_ctrl_ia_capability.f.initialize_inc );
tran (sa_ctrl_ia_capability[6], \sa_ctrl_ia_capability.r.part0 [6]);
tran (sa_ctrl_ia_capability[6], \sa_ctrl_ia_capability.f.initialize );
tran (sa_ctrl_ia_capability[5], \sa_ctrl_ia_capability.r.part0 [5]);
tran (sa_ctrl_ia_capability[5], \sa_ctrl_ia_capability.f.reset );
tran (sa_ctrl_ia_capability[4], \sa_ctrl_ia_capability.r.part0 [4]);
tran (sa_ctrl_ia_capability[4], \sa_ctrl_ia_capability.f.disabled );
tran (sa_ctrl_ia_capability[3], \sa_ctrl_ia_capability.r.part0 [3]);
tran (sa_ctrl_ia_capability[3], \sa_ctrl_ia_capability.f.enable );
tran (sa_ctrl_ia_capability[2], \sa_ctrl_ia_capability.r.part0 [2]);
tran (sa_ctrl_ia_capability[2], \sa_ctrl_ia_capability.f.write );
tran (sa_ctrl_ia_capability[1], \sa_ctrl_ia_capability.r.part0 [1]);
tran (sa_ctrl_ia_capability[1], \sa_ctrl_ia_capability.f.read );
tran (sa_ctrl_ia_capability[0], \sa_ctrl_ia_capability.r.part0 [0]);
tran (sa_ctrl_ia_capability[0], \sa_ctrl_ia_capability.f.nop );
tran (sa_ctrl_ia_capability[19], \sa_ctrl_ia_capability.r.part0 [19]);
tran (sa_ctrl_ia_capability[19], \sa_ctrl_ia_capability.f.mem_type [3]);
tran (sa_ctrl_ia_capability[18], \sa_ctrl_ia_capability.r.part0 [18]);
tran (sa_ctrl_ia_capability[18], \sa_ctrl_ia_capability.f.mem_type [2]);
tran (sa_ctrl_ia_capability[17], \sa_ctrl_ia_capability.r.part0 [17]);
tran (sa_ctrl_ia_capability[17], \sa_ctrl_ia_capability.f.mem_type [1]);
tran (sa_ctrl_ia_capability[16], \sa_ctrl_ia_capability.r.part0 [16]);
tran (sa_ctrl_ia_capability[16], \sa_ctrl_ia_capability.f.mem_type [0]);
tran (sa_ctrl_ia_rdata[31], \sa_ctrl_ia_rdata.r.part0 [31]);
tran (sa_ctrl_ia_rdata[31], \sa_ctrl_ia_rdata.f.spare [26]);
tran (sa_ctrl_ia_rdata[30], \sa_ctrl_ia_rdata.r.part0 [30]);
tran (sa_ctrl_ia_rdata[30], \sa_ctrl_ia_rdata.f.spare [25]);
tran (sa_ctrl_ia_rdata[29], \sa_ctrl_ia_rdata.r.part0 [29]);
tran (sa_ctrl_ia_rdata[29], \sa_ctrl_ia_rdata.f.spare [24]);
tran (sa_ctrl_ia_rdata[28], \sa_ctrl_ia_rdata.r.part0 [28]);
tran (sa_ctrl_ia_rdata[28], \sa_ctrl_ia_rdata.f.spare [23]);
tran (sa_ctrl_ia_rdata[27], \sa_ctrl_ia_rdata.r.part0 [27]);
tran (sa_ctrl_ia_rdata[27], \sa_ctrl_ia_rdata.f.spare [22]);
tran (sa_ctrl_ia_rdata[26], \sa_ctrl_ia_rdata.r.part0 [26]);
tran (sa_ctrl_ia_rdata[26], \sa_ctrl_ia_rdata.f.spare [21]);
tran (sa_ctrl_ia_rdata[25], \sa_ctrl_ia_rdata.r.part0 [25]);
tran (sa_ctrl_ia_rdata[25], \sa_ctrl_ia_rdata.f.spare [20]);
tran (sa_ctrl_ia_rdata[24], \sa_ctrl_ia_rdata.r.part0 [24]);
tran (sa_ctrl_ia_rdata[24], \sa_ctrl_ia_rdata.f.spare [19]);
tran (sa_ctrl_ia_rdata[23], \sa_ctrl_ia_rdata.r.part0 [23]);
tran (sa_ctrl_ia_rdata[23], \sa_ctrl_ia_rdata.f.spare [18]);
tran (sa_ctrl_ia_rdata[22], \sa_ctrl_ia_rdata.r.part0 [22]);
tran (sa_ctrl_ia_rdata[22], \sa_ctrl_ia_rdata.f.spare [17]);
tran (sa_ctrl_ia_rdata[21], \sa_ctrl_ia_rdata.r.part0 [21]);
tran (sa_ctrl_ia_rdata[21], \sa_ctrl_ia_rdata.f.spare [16]);
tran (sa_ctrl_ia_rdata[20], \sa_ctrl_ia_rdata.r.part0 [20]);
tran (sa_ctrl_ia_rdata[20], \sa_ctrl_ia_rdata.f.spare [15]);
tran (sa_ctrl_ia_rdata[19], \sa_ctrl_ia_rdata.r.part0 [19]);
tran (sa_ctrl_ia_rdata[19], \sa_ctrl_ia_rdata.f.spare [14]);
tran (sa_ctrl_ia_rdata[18], \sa_ctrl_ia_rdata.r.part0 [18]);
tran (sa_ctrl_ia_rdata[18], \sa_ctrl_ia_rdata.f.spare [13]);
tran (sa_ctrl_ia_rdata[17], \sa_ctrl_ia_rdata.r.part0 [17]);
tran (sa_ctrl_ia_rdata[17], \sa_ctrl_ia_rdata.f.spare [12]);
tran (sa_ctrl_ia_rdata[16], \sa_ctrl_ia_rdata.r.part0 [16]);
tran (sa_ctrl_ia_rdata[16], \sa_ctrl_ia_rdata.f.spare [11]);
tran (sa_ctrl_ia_rdata[15], \sa_ctrl_ia_rdata.r.part0 [15]);
tran (sa_ctrl_ia_rdata[15], \sa_ctrl_ia_rdata.f.spare [10]);
tran (sa_ctrl_ia_rdata[14], \sa_ctrl_ia_rdata.r.part0 [14]);
tran (sa_ctrl_ia_rdata[14], \sa_ctrl_ia_rdata.f.spare [9]);
tran (sa_ctrl_ia_rdata[13], \sa_ctrl_ia_rdata.r.part0 [13]);
tran (sa_ctrl_ia_rdata[13], \sa_ctrl_ia_rdata.f.spare [8]);
tran (sa_ctrl_ia_rdata[12], \sa_ctrl_ia_rdata.r.part0 [12]);
tran (sa_ctrl_ia_rdata[12], \sa_ctrl_ia_rdata.f.spare [7]);
tran (sa_ctrl_ia_rdata[11], \sa_ctrl_ia_rdata.r.part0 [11]);
tran (sa_ctrl_ia_rdata[11], \sa_ctrl_ia_rdata.f.spare [6]);
tran (sa_ctrl_ia_rdata[10], \sa_ctrl_ia_rdata.r.part0 [10]);
tran (sa_ctrl_ia_rdata[10], \sa_ctrl_ia_rdata.f.spare [5]);
tran (sa_ctrl_ia_rdata[9], \sa_ctrl_ia_rdata.r.part0 [9]);
tran (sa_ctrl_ia_rdata[9], \sa_ctrl_ia_rdata.f.spare [4]);
tran (sa_ctrl_ia_rdata[8], \sa_ctrl_ia_rdata.r.part0 [8]);
tran (sa_ctrl_ia_rdata[8], \sa_ctrl_ia_rdata.f.spare [3]);
tran (sa_ctrl_ia_rdata[7], \sa_ctrl_ia_rdata.r.part0 [7]);
tran (sa_ctrl_ia_rdata[7], \sa_ctrl_ia_rdata.f.spare [2]);
tran (sa_ctrl_ia_rdata[6], \sa_ctrl_ia_rdata.r.part0 [6]);
tran (sa_ctrl_ia_rdata[6], \sa_ctrl_ia_rdata.f.spare [1]);
tran (sa_ctrl_ia_rdata[5], \sa_ctrl_ia_rdata.r.part0 [5]);
tran (sa_ctrl_ia_rdata[5], \sa_ctrl_ia_rdata.f.spare [0]);
tran (sa_ctrl_ia_rdata[4], \sa_ctrl_ia_rdata.r.part0 [4]);
tran (sa_ctrl_ia_rdata[4], \sa_ctrl_ia_rdata.f.sa_event_sel [4]);
tran (sa_ctrl_ia_rdata[3], \sa_ctrl_ia_rdata.r.part0 [3]);
tran (sa_ctrl_ia_rdata[3], \sa_ctrl_ia_rdata.f.sa_event_sel [3]);
tran (sa_ctrl_ia_rdata[2], \sa_ctrl_ia_rdata.r.part0 [2]);
tran (sa_ctrl_ia_rdata[2], \sa_ctrl_ia_rdata.f.sa_event_sel [2]);
tran (sa_ctrl_ia_rdata[1], \sa_ctrl_ia_rdata.r.part0 [1]);
tran (sa_ctrl_ia_rdata[1], \sa_ctrl_ia_rdata.f.sa_event_sel [1]);
tran (sa_ctrl_ia_rdata[0], \sa_ctrl_ia_rdata.r.part0 [0]);
tran (sa_ctrl_ia_rdata[0], \sa_ctrl_ia_rdata.f.sa_event_sel [0]);
tran (cceip0_im_din[22], \cceip0_im_din.desc.im_meta [22]);
tran (cceip0_im_din[21], \cceip0_im_din.desc.im_meta [21]);
tran (cceip0_im_din[20], \cceip0_im_din.desc.im_meta [20]);
tran (cceip0_im_din[19], \cceip0_im_din.desc.im_meta [19]);
tran (cceip0_im_din[18], \cceip0_im_din.desc.im_meta [18]);
tran (cceip0_im_din[17], \cceip0_im_din.desc.im_meta [17]);
tran (cceip0_im_din[16], \cceip0_im_din.desc.im_meta [16]);
tran (cceip0_im_din[15], \cceip0_im_din.desc.im_meta [15]);
tran (cceip0_im_din[5], \cceip0_im_din.desc.im_meta [5]);
tran (cceip0_im_din[4], \cceip0_im_din.desc.im_meta [4]);
tran (cceip0_im_din[3], \cceip0_im_din.desc.im_meta [3]);
tran (cceip0_im_din[2], \cceip0_im_din.desc.im_meta [2]);
tran (cceip0_im_din[1], \cceip0_im_din.desc.im_meta [1]);
tran (cceip0_im_din[0], \cceip0_im_din.desc.im_meta [0]);
tran (cddip0_im_din[22], \cddip0_im_din.desc.im_meta [22]);
tran (cddip0_im_din[21], \cddip0_im_din.desc.im_meta [21]);
tran (cddip0_im_din[20], \cddip0_im_din.desc.im_meta [20]);
tran (cddip0_im_din[19], \cddip0_im_din.desc.im_meta [19]);
tran (cddip0_im_din[18], \cddip0_im_din.desc.im_meta [18]);
tran (cddip0_im_din[17], \cddip0_im_din.desc.im_meta [17]);
tran (cddip0_im_din[16], \cddip0_im_din.desc.im_meta [16]);
tran (cddip0_im_din[15], \cddip0_im_din.desc.im_meta [15]);
tran (cddip0_im_din[5], \cddip0_im_din.desc.im_meta [5]);
tran (cddip0_im_din[4], \cddip0_im_din.desc.im_meta [4]);
tran (cddip0_im_din[3], \cddip0_im_din.desc.im_meta [3]);
tran (cddip0_im_din[2], \cddip0_im_din.desc.im_meta [2]);
tran (cddip0_im_din[1], \cddip0_im_din.desc.im_meta [1]);
tran (cddip0_im_din[0], \cddip0_im_din.desc.im_meta [0]);
tran (cceip1_im_din[22], \cceip1_im_din.desc.im_meta [22]);
tran (cceip1_im_din[21], \cceip1_im_din.desc.im_meta [21]);
tran (cceip1_im_din[20], \cceip1_im_din.desc.im_meta [20]);
tran (cceip1_im_din[19], \cceip1_im_din.desc.im_meta [19]);
tran (cceip1_im_din[18], \cceip1_im_din.desc.im_meta [18]);
tran (cceip1_im_din[17], \cceip1_im_din.desc.im_meta [17]);
tran (cceip1_im_din[16], \cceip1_im_din.desc.im_meta [16]);
tran (cceip1_im_din[15], \cceip1_im_din.desc.im_meta [15]);
tran (cceip1_im_din[5], \cceip1_im_din.desc.im_meta [5]);
tran (cceip1_im_din[4], \cceip1_im_din.desc.im_meta [4]);
tran (cceip1_im_din[3], \cceip1_im_din.desc.im_meta [3]);
tran (cceip1_im_din[2], \cceip1_im_din.desc.im_meta [2]);
tran (cceip1_im_din[1], \cceip1_im_din.desc.im_meta [1]);
tran (cceip1_im_din[0], \cceip1_im_din.desc.im_meta [0]);
tran (cddip1_im_din[22], \cddip1_im_din.desc.im_meta [22]);
tran (cddip1_im_din[21], \cddip1_im_din.desc.im_meta [21]);
tran (cddip1_im_din[20], \cddip1_im_din.desc.im_meta [20]);
tran (cddip1_im_din[19], \cddip1_im_din.desc.im_meta [19]);
tran (cddip1_im_din[18], \cddip1_im_din.desc.im_meta [18]);
tran (cddip1_im_din[17], \cddip1_im_din.desc.im_meta [17]);
tran (cddip1_im_din[16], \cddip1_im_din.desc.im_meta [16]);
tran (cddip1_im_din[15], \cddip1_im_din.desc.im_meta [15]);
tran (cddip1_im_din[5], \cddip1_im_din.desc.im_meta [5]);
tran (cddip1_im_din[4], \cddip1_im_din.desc.im_meta [4]);
tran (cddip1_im_din[3], \cddip1_im_din.desc.im_meta [3]);
tran (cddip1_im_din[2], \cddip1_im_din.desc.im_meta [2]);
tran (cddip1_im_din[1], \cddip1_im_din.desc.im_meta [1]);
tran (cddip1_im_din[0], \cddip1_im_din.desc.im_meta [0]);
tran (cceip2_im_din[22], \cceip2_im_din.desc.im_meta [22]);
tran (cceip2_im_din[21], \cceip2_im_din.desc.im_meta [21]);
tran (cceip2_im_din[20], \cceip2_im_din.desc.im_meta [20]);
tran (cceip2_im_din[19], \cceip2_im_din.desc.im_meta [19]);
tran (cceip2_im_din[18], \cceip2_im_din.desc.im_meta [18]);
tran (cceip2_im_din[17], \cceip2_im_din.desc.im_meta [17]);
tran (cceip2_im_din[16], \cceip2_im_din.desc.im_meta [16]);
tran (cceip2_im_din[15], \cceip2_im_din.desc.im_meta [15]);
tran (cceip2_im_din[5], \cceip2_im_din.desc.im_meta [5]);
tran (cceip2_im_din[4], \cceip2_im_din.desc.im_meta [4]);
tran (cceip2_im_din[3], \cceip2_im_din.desc.im_meta [3]);
tran (cceip2_im_din[2], \cceip2_im_din.desc.im_meta [2]);
tran (cceip2_im_din[1], \cceip2_im_din.desc.im_meta [1]);
tran (cceip2_im_din[0], \cceip2_im_din.desc.im_meta [0]);
tran (cddip2_im_din[22], \cddip2_im_din.desc.im_meta [22]);
tran (cddip2_im_din[21], \cddip2_im_din.desc.im_meta [21]);
tran (cddip2_im_din[20], \cddip2_im_din.desc.im_meta [20]);
tran (cddip2_im_din[19], \cddip2_im_din.desc.im_meta [19]);
tran (cddip2_im_din[18], \cddip2_im_din.desc.im_meta [18]);
tran (cddip2_im_din[17], \cddip2_im_din.desc.im_meta [17]);
tran (cddip2_im_din[16], \cddip2_im_din.desc.im_meta [16]);
tran (cddip2_im_din[15], \cddip2_im_din.desc.im_meta [15]);
tran (cddip2_im_din[5], \cddip2_im_din.desc.im_meta [5]);
tran (cddip2_im_din[4], \cddip2_im_din.desc.im_meta [4]);
tran (cddip2_im_din[3], \cddip2_im_din.desc.im_meta [3]);
tran (cddip2_im_din[2], \cddip2_im_din.desc.im_meta [2]);
tran (cddip2_im_din[1], \cddip2_im_din.desc.im_meta [1]);
tran (cddip2_im_din[0], \cddip2_im_din.desc.im_meta [0]);
tran (cceip3_im_din[22], \cceip3_im_din.desc.im_meta [22]);
tran (cceip3_im_din[21], \cceip3_im_din.desc.im_meta [21]);
tran (cceip3_im_din[20], \cceip3_im_din.desc.im_meta [20]);
tran (cceip3_im_din[19], \cceip3_im_din.desc.im_meta [19]);
tran (cceip3_im_din[18], \cceip3_im_din.desc.im_meta [18]);
tran (cceip3_im_din[17], \cceip3_im_din.desc.im_meta [17]);
tran (cceip3_im_din[16], \cceip3_im_din.desc.im_meta [16]);
tran (cceip3_im_din[15], \cceip3_im_din.desc.im_meta [15]);
tran (cceip3_im_din[5], \cceip3_im_din.desc.im_meta [5]);
tran (cceip3_im_din[4], \cceip3_im_din.desc.im_meta [4]);
tran (cceip3_im_din[3], \cceip3_im_din.desc.im_meta [3]);
tran (cceip3_im_din[2], \cceip3_im_din.desc.im_meta [2]);
tran (cceip3_im_din[1], \cceip3_im_din.desc.im_meta [1]);
tran (cceip3_im_din[0], \cceip3_im_din.desc.im_meta [0]);
tran (cddip3_im_din[22], \cddip3_im_din.desc.im_meta [22]);
tran (cddip3_im_din[21], \cddip3_im_din.desc.im_meta [21]);
tran (cddip3_im_din[20], \cddip3_im_din.desc.im_meta [20]);
tran (cddip3_im_din[19], \cddip3_im_din.desc.im_meta [19]);
tran (cddip3_im_din[18], \cddip3_im_din.desc.im_meta [18]);
tran (cddip3_im_din[17], \cddip3_im_din.desc.im_meta [17]);
tran (cddip3_im_din[16], \cddip3_im_din.desc.im_meta [16]);
tran (cddip3_im_din[15], \cddip3_im_din.desc.im_meta [15]);
tran (cddip3_im_din[5], \cddip3_im_din.desc.im_meta [5]);
tran (cddip3_im_din[4], \cddip3_im_din.desc.im_meta [4]);
tran (cddip3_im_din[3], \cddip3_im_din.desc.im_meta [3]);
tran (cddip3_im_din[2], \cddip3_im_din.desc.im_meta [2]);
tran (cddip3_im_din[1], \cddip3_im_din.desc.im_meta [1]);
tran (cddip3_im_din[0], \cddip3_im_din.desc.im_meta [0]);
tran (revid_wire[7], \revid_wire.r.part0 [7]);
tran (revid_wire[7], \revid_wire.f.revid [7]);
tran (revid_wire[6], \revid_wire.r.part0 [6]);
tran (revid_wire[6], \revid_wire.f.revid [6]);
tran (revid_wire[5], \revid_wire.r.part0 [5]);
tran (revid_wire[5], \revid_wire.f.revid [5]);
tran (revid_wire[4], \revid_wire.r.part0 [4]);
tran (revid_wire[4], \revid_wire.f.revid [4]);
tran (revid_wire[3], \revid_wire.r.part0 [3]);
tran (revid_wire[3], \revid_wire.f.revid [3]);
tran (revid_wire[2], \revid_wire.r.part0 [2]);
tran (revid_wire[2], \revid_wire.f.revid [2]);
tran (revid_wire[1], \revid_wire.r.part0 [1]);
tran (revid_wire[1], \revid_wire.f.revid [1]);
tran (revid_wire[0], \revid_wire.r.part0 [0]);
tran (revid_wire[0], \revid_wire.f.revid [0]);
tran (im_available_kme_cddip3[1], \im_available_kme_cddip3.bank_hi );
tran (im_available_kme_cddip3[0], \im_available_kme_cddip3.bank_lo );
tran (im_available_kme_cddip2[1], \im_available_kme_cddip2.bank_hi );
tran (im_available_kme_cddip2[0], \im_available_kme_cddip2.bank_lo );
tran (im_available_kme_cddip1[1], \im_available_kme_cddip1.bank_hi );
tran (im_available_kme_cddip1[0], \im_available_kme_cddip1.bank_lo );
tran (im_available_kme_cddip0[1], \im_available_kme_cddip0.bank_hi );
tran (im_available_kme_cddip0[0], \im_available_kme_cddip0.bank_lo );
tran (im_available_kme_cceip3[1], \im_available_kme_cceip3.bank_hi );
tran (im_available_kme_cceip3[0], \im_available_kme_cceip3.bank_lo );
tran (im_available_kme_cceip2[1], \im_available_kme_cceip2.bank_hi );
tran (im_available_kme_cceip2[0], \im_available_kme_cceip2.bank_lo );
tran (im_available_kme_cceip1[1], \im_available_kme_cceip1.bank_hi );
tran (im_available_kme_cceip1[0], \im_available_kme_cceip1.bank_lo );
tran (im_available_kme_cceip0[1], \im_available_kme_cceip0.bank_hi );
tran (im_available_kme_cceip0[0], \im_available_kme_cceip0.bank_lo );
tran (im_consumed_kme_cceip0[1], \im_consumed_kme_cceip0.bank_hi );
tran (im_consumed_kme_cceip0[0], \im_consumed_kme_cceip0.bank_lo );
tran (im_consumed_kme_cddip0[1], \im_consumed_kme_cddip0.bank_hi );
tran (im_consumed_kme_cddip0[0], \im_consumed_kme_cddip0.bank_lo );
tran (im_consumed_kme_cceip1[1], \im_consumed_kme_cceip1.bank_hi );
tran (im_consumed_kme_cceip1[0], \im_consumed_kme_cceip1.bank_lo );
tran (im_consumed_kme_cddip1[1], \im_consumed_kme_cddip1.bank_hi );
tran (im_consumed_kme_cddip1[0], \im_consumed_kme_cddip1.bank_lo );
tran (im_consumed_kme_cceip2[1], \im_consumed_kme_cceip2.bank_hi );
tran (im_consumed_kme_cceip2[0], \im_consumed_kme_cceip2.bank_lo );
tran (im_consumed_kme_cddip2[1], \im_consumed_kme_cddip2.bank_hi );
tran (im_consumed_kme_cddip2[0], \im_consumed_kme_cddip2.bank_lo );
tran (im_consumed_kme_cceip3[1], \im_consumed_kme_cceip3.bank_hi );
tran (im_consumed_kme_cceip3[0], \im_consumed_kme_cceip3.bank_lo );
tran (im_consumed_kme_cddip3[1], \im_consumed_kme_cddip3.bank_hi );
tran (im_consumed_kme_cddip3[0], \im_consumed_kme_cddip3.bank_lo );
tran (\sa_ctrl_rst_dat[0][0] , \sa_ctrl_rst_dat[0].r.part0[0] );
tran (\sa_ctrl_rst_dat[0][0] , \sa_ctrl_rst_dat[0].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[0][1] , \sa_ctrl_rst_dat[0].r.part0[1] );
tran (\sa_ctrl_rst_dat[0][1] , \sa_ctrl_rst_dat[0].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[0][2] , \sa_ctrl_rst_dat[0].r.part0[2] );
tran (\sa_ctrl_rst_dat[0][2] , \sa_ctrl_rst_dat[0].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[0][3] , \sa_ctrl_rst_dat[0].r.part0[3] );
tran (\sa_ctrl_rst_dat[0][3] , \sa_ctrl_rst_dat[0].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[0][4] , \sa_ctrl_rst_dat[0].r.part0[4] );
tran (\sa_ctrl_rst_dat[0][4] , \sa_ctrl_rst_dat[0].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[0][5] , \sa_ctrl_rst_dat[0].r.part0[5] );
tran (\sa_ctrl_rst_dat[0][5] , \sa_ctrl_rst_dat[0].f.spare[0] );
tran (\sa_ctrl_rst_dat[0][6] , \sa_ctrl_rst_dat[0].r.part0[6] );
tran (\sa_ctrl_rst_dat[0][6] , \sa_ctrl_rst_dat[0].f.spare[1] );
tran (\sa_ctrl_rst_dat[0][7] , \sa_ctrl_rst_dat[0].r.part0[7] );
tran (\sa_ctrl_rst_dat[0][7] , \sa_ctrl_rst_dat[0].f.spare[2] );
tran (\sa_ctrl_rst_dat[0][8] , \sa_ctrl_rst_dat[0].r.part0[8] );
tran (\sa_ctrl_rst_dat[0][8] , \sa_ctrl_rst_dat[0].f.spare[3] );
tran (\sa_ctrl_rst_dat[0][9] , \sa_ctrl_rst_dat[0].r.part0[9] );
tran (\sa_ctrl_rst_dat[0][9] , \sa_ctrl_rst_dat[0].f.spare[4] );
tran (\sa_ctrl_rst_dat[0][10] , \sa_ctrl_rst_dat[0].r.part0[10] );
tran (\sa_ctrl_rst_dat[0][10] , \sa_ctrl_rst_dat[0].f.spare[5] );
tran (\sa_ctrl_rst_dat[0][11] , \sa_ctrl_rst_dat[0].r.part0[11] );
tran (\sa_ctrl_rst_dat[0][11] , \sa_ctrl_rst_dat[0].f.spare[6] );
tran (\sa_ctrl_rst_dat[0][12] , \sa_ctrl_rst_dat[0].r.part0[12] );
tran (\sa_ctrl_rst_dat[0][12] , \sa_ctrl_rst_dat[0].f.spare[7] );
tran (\sa_ctrl_rst_dat[0][13] , \sa_ctrl_rst_dat[0].r.part0[13] );
tran (\sa_ctrl_rst_dat[0][13] , \sa_ctrl_rst_dat[0].f.spare[8] );
tran (\sa_ctrl_rst_dat[0][14] , \sa_ctrl_rst_dat[0].r.part0[14] );
tran (\sa_ctrl_rst_dat[0][14] , \sa_ctrl_rst_dat[0].f.spare[9] );
tran (\sa_ctrl_rst_dat[0][15] , \sa_ctrl_rst_dat[0].r.part0[15] );
tran (\sa_ctrl_rst_dat[0][15] , \sa_ctrl_rst_dat[0].f.spare[10] );
tran (\sa_ctrl_rst_dat[0][16] , \sa_ctrl_rst_dat[0].r.part0[16] );
tran (\sa_ctrl_rst_dat[0][16] , \sa_ctrl_rst_dat[0].f.spare[11] );
tran (\sa_ctrl_rst_dat[0][17] , \sa_ctrl_rst_dat[0].r.part0[17] );
tran (\sa_ctrl_rst_dat[0][17] , \sa_ctrl_rst_dat[0].f.spare[12] );
tran (\sa_ctrl_rst_dat[0][18] , \sa_ctrl_rst_dat[0].r.part0[18] );
tran (\sa_ctrl_rst_dat[0][18] , \sa_ctrl_rst_dat[0].f.spare[13] );
tran (\sa_ctrl_rst_dat[0][19] , \sa_ctrl_rst_dat[0].r.part0[19] );
tran (\sa_ctrl_rst_dat[0][19] , \sa_ctrl_rst_dat[0].f.spare[14] );
tran (\sa_ctrl_rst_dat[0][20] , \sa_ctrl_rst_dat[0].r.part0[20] );
tran (\sa_ctrl_rst_dat[0][20] , \sa_ctrl_rst_dat[0].f.spare[15] );
tran (\sa_ctrl_rst_dat[0][21] , \sa_ctrl_rst_dat[0].r.part0[21] );
tran (\sa_ctrl_rst_dat[0][21] , \sa_ctrl_rst_dat[0].f.spare[16] );
tran (\sa_ctrl_rst_dat[0][22] , \sa_ctrl_rst_dat[0].r.part0[22] );
tran (\sa_ctrl_rst_dat[0][22] , \sa_ctrl_rst_dat[0].f.spare[17] );
tran (\sa_ctrl_rst_dat[0][23] , \sa_ctrl_rst_dat[0].r.part0[23] );
tran (\sa_ctrl_rst_dat[0][23] , \sa_ctrl_rst_dat[0].f.spare[18] );
tran (\sa_ctrl_rst_dat[0][24] , \sa_ctrl_rst_dat[0].r.part0[24] );
tran (\sa_ctrl_rst_dat[0][24] , \sa_ctrl_rst_dat[0].f.spare[19] );
tran (\sa_ctrl_rst_dat[0][25] , \sa_ctrl_rst_dat[0].r.part0[25] );
tran (\sa_ctrl_rst_dat[0][25] , \sa_ctrl_rst_dat[0].f.spare[20] );
tran (\sa_ctrl_rst_dat[0][26] , \sa_ctrl_rst_dat[0].r.part0[26] );
tran (\sa_ctrl_rst_dat[0][26] , \sa_ctrl_rst_dat[0].f.spare[21] );
tran (\sa_ctrl_rst_dat[0][27] , \sa_ctrl_rst_dat[0].r.part0[27] );
tran (\sa_ctrl_rst_dat[0][27] , \sa_ctrl_rst_dat[0].f.spare[22] );
tran (\sa_ctrl_rst_dat[0][28] , \sa_ctrl_rst_dat[0].r.part0[28] );
tran (\sa_ctrl_rst_dat[0][28] , \sa_ctrl_rst_dat[0].f.spare[23] );
tran (\sa_ctrl_rst_dat[0][29] , \sa_ctrl_rst_dat[0].r.part0[29] );
tran (\sa_ctrl_rst_dat[0][29] , \sa_ctrl_rst_dat[0].f.spare[24] );
tran (\sa_ctrl_rst_dat[0][30] , \sa_ctrl_rst_dat[0].r.part0[30] );
tran (\sa_ctrl_rst_dat[0][30] , \sa_ctrl_rst_dat[0].f.spare[25] );
tran (\sa_ctrl_rst_dat[0][31] , \sa_ctrl_rst_dat[0].r.part0[31] );
tran (\sa_ctrl_rst_dat[0][31] , \sa_ctrl_rst_dat[0].f.spare[26] );
tran (\sa_ctrl_rst_dat[1][0] , \sa_ctrl_rst_dat[1].r.part0[0] );
tran (\sa_ctrl_rst_dat[1][0] , \sa_ctrl_rst_dat[1].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[1][1] , \sa_ctrl_rst_dat[1].r.part0[1] );
tran (\sa_ctrl_rst_dat[1][1] , \sa_ctrl_rst_dat[1].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[1][2] , \sa_ctrl_rst_dat[1].r.part0[2] );
tran (\sa_ctrl_rst_dat[1][2] , \sa_ctrl_rst_dat[1].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[1][3] , \sa_ctrl_rst_dat[1].r.part0[3] );
tran (\sa_ctrl_rst_dat[1][3] , \sa_ctrl_rst_dat[1].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[1][4] , \sa_ctrl_rst_dat[1].r.part0[4] );
tran (\sa_ctrl_rst_dat[1][4] , \sa_ctrl_rst_dat[1].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[1][5] , \sa_ctrl_rst_dat[1].r.part0[5] );
tran (\sa_ctrl_rst_dat[1][5] , \sa_ctrl_rst_dat[1].f.spare[0] );
tran (\sa_ctrl_rst_dat[1][6] , \sa_ctrl_rst_dat[1].r.part0[6] );
tran (\sa_ctrl_rst_dat[1][6] , \sa_ctrl_rst_dat[1].f.spare[1] );
tran (\sa_ctrl_rst_dat[1][7] , \sa_ctrl_rst_dat[1].r.part0[7] );
tran (\sa_ctrl_rst_dat[1][7] , \sa_ctrl_rst_dat[1].f.spare[2] );
tran (\sa_ctrl_rst_dat[1][8] , \sa_ctrl_rst_dat[1].r.part0[8] );
tran (\sa_ctrl_rst_dat[1][8] , \sa_ctrl_rst_dat[1].f.spare[3] );
tran (\sa_ctrl_rst_dat[1][9] , \sa_ctrl_rst_dat[1].r.part0[9] );
tran (\sa_ctrl_rst_dat[1][9] , \sa_ctrl_rst_dat[1].f.spare[4] );
tran (\sa_ctrl_rst_dat[1][10] , \sa_ctrl_rst_dat[1].r.part0[10] );
tran (\sa_ctrl_rst_dat[1][10] , \sa_ctrl_rst_dat[1].f.spare[5] );
tran (\sa_ctrl_rst_dat[1][11] , \sa_ctrl_rst_dat[1].r.part0[11] );
tran (\sa_ctrl_rst_dat[1][11] , \sa_ctrl_rst_dat[1].f.spare[6] );
tran (\sa_ctrl_rst_dat[1][12] , \sa_ctrl_rst_dat[1].r.part0[12] );
tran (\sa_ctrl_rst_dat[1][12] , \sa_ctrl_rst_dat[1].f.spare[7] );
tran (\sa_ctrl_rst_dat[1][13] , \sa_ctrl_rst_dat[1].r.part0[13] );
tran (\sa_ctrl_rst_dat[1][13] , \sa_ctrl_rst_dat[1].f.spare[8] );
tran (\sa_ctrl_rst_dat[1][14] , \sa_ctrl_rst_dat[1].r.part0[14] );
tran (\sa_ctrl_rst_dat[1][14] , \sa_ctrl_rst_dat[1].f.spare[9] );
tran (\sa_ctrl_rst_dat[1][15] , \sa_ctrl_rst_dat[1].r.part0[15] );
tran (\sa_ctrl_rst_dat[1][15] , \sa_ctrl_rst_dat[1].f.spare[10] );
tran (\sa_ctrl_rst_dat[1][16] , \sa_ctrl_rst_dat[1].r.part0[16] );
tran (\sa_ctrl_rst_dat[1][16] , \sa_ctrl_rst_dat[1].f.spare[11] );
tran (\sa_ctrl_rst_dat[1][17] , \sa_ctrl_rst_dat[1].r.part0[17] );
tran (\sa_ctrl_rst_dat[1][17] , \sa_ctrl_rst_dat[1].f.spare[12] );
tran (\sa_ctrl_rst_dat[1][18] , \sa_ctrl_rst_dat[1].r.part0[18] );
tran (\sa_ctrl_rst_dat[1][18] , \sa_ctrl_rst_dat[1].f.spare[13] );
tran (\sa_ctrl_rst_dat[1][19] , \sa_ctrl_rst_dat[1].r.part0[19] );
tran (\sa_ctrl_rst_dat[1][19] , \sa_ctrl_rst_dat[1].f.spare[14] );
tran (\sa_ctrl_rst_dat[1][20] , \sa_ctrl_rst_dat[1].r.part0[20] );
tran (\sa_ctrl_rst_dat[1][20] , \sa_ctrl_rst_dat[1].f.spare[15] );
tran (\sa_ctrl_rst_dat[1][21] , \sa_ctrl_rst_dat[1].r.part0[21] );
tran (\sa_ctrl_rst_dat[1][21] , \sa_ctrl_rst_dat[1].f.spare[16] );
tran (\sa_ctrl_rst_dat[1][22] , \sa_ctrl_rst_dat[1].r.part0[22] );
tran (\sa_ctrl_rst_dat[1][22] , \sa_ctrl_rst_dat[1].f.spare[17] );
tran (\sa_ctrl_rst_dat[1][23] , \sa_ctrl_rst_dat[1].r.part0[23] );
tran (\sa_ctrl_rst_dat[1][23] , \sa_ctrl_rst_dat[1].f.spare[18] );
tran (\sa_ctrl_rst_dat[1][24] , \sa_ctrl_rst_dat[1].r.part0[24] );
tran (\sa_ctrl_rst_dat[1][24] , \sa_ctrl_rst_dat[1].f.spare[19] );
tran (\sa_ctrl_rst_dat[1][25] , \sa_ctrl_rst_dat[1].r.part0[25] );
tran (\sa_ctrl_rst_dat[1][25] , \sa_ctrl_rst_dat[1].f.spare[20] );
tran (\sa_ctrl_rst_dat[1][26] , \sa_ctrl_rst_dat[1].r.part0[26] );
tran (\sa_ctrl_rst_dat[1][26] , \sa_ctrl_rst_dat[1].f.spare[21] );
tran (\sa_ctrl_rst_dat[1][27] , \sa_ctrl_rst_dat[1].r.part0[27] );
tran (\sa_ctrl_rst_dat[1][27] , \sa_ctrl_rst_dat[1].f.spare[22] );
tran (\sa_ctrl_rst_dat[1][28] , \sa_ctrl_rst_dat[1].r.part0[28] );
tran (\sa_ctrl_rst_dat[1][28] , \sa_ctrl_rst_dat[1].f.spare[23] );
tran (\sa_ctrl_rst_dat[1][29] , \sa_ctrl_rst_dat[1].r.part0[29] );
tran (\sa_ctrl_rst_dat[1][29] , \sa_ctrl_rst_dat[1].f.spare[24] );
tran (\sa_ctrl_rst_dat[1][30] , \sa_ctrl_rst_dat[1].r.part0[30] );
tran (\sa_ctrl_rst_dat[1][30] , \sa_ctrl_rst_dat[1].f.spare[25] );
tran (\sa_ctrl_rst_dat[1][31] , \sa_ctrl_rst_dat[1].r.part0[31] );
tran (\sa_ctrl_rst_dat[1][31] , \sa_ctrl_rst_dat[1].f.spare[26] );
tran (\sa_ctrl_rst_dat[2][0] , \sa_ctrl_rst_dat[2].r.part0[0] );
tran (\sa_ctrl_rst_dat[2][0] , \sa_ctrl_rst_dat[2].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[2][1] , \sa_ctrl_rst_dat[2].r.part0[1] );
tran (\sa_ctrl_rst_dat[2][1] , \sa_ctrl_rst_dat[2].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[2][2] , \sa_ctrl_rst_dat[2].r.part0[2] );
tran (\sa_ctrl_rst_dat[2][2] , \sa_ctrl_rst_dat[2].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[2][3] , \sa_ctrl_rst_dat[2].r.part0[3] );
tran (\sa_ctrl_rst_dat[2][3] , \sa_ctrl_rst_dat[2].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[2][4] , \sa_ctrl_rst_dat[2].r.part0[4] );
tran (\sa_ctrl_rst_dat[2][4] , \sa_ctrl_rst_dat[2].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[2][5] , \sa_ctrl_rst_dat[2].r.part0[5] );
tran (\sa_ctrl_rst_dat[2][5] , \sa_ctrl_rst_dat[2].f.spare[0] );
tran (\sa_ctrl_rst_dat[2][6] , \sa_ctrl_rst_dat[2].r.part0[6] );
tran (\sa_ctrl_rst_dat[2][6] , \sa_ctrl_rst_dat[2].f.spare[1] );
tran (\sa_ctrl_rst_dat[2][7] , \sa_ctrl_rst_dat[2].r.part0[7] );
tran (\sa_ctrl_rst_dat[2][7] , \sa_ctrl_rst_dat[2].f.spare[2] );
tran (\sa_ctrl_rst_dat[2][8] , \sa_ctrl_rst_dat[2].r.part0[8] );
tran (\sa_ctrl_rst_dat[2][8] , \sa_ctrl_rst_dat[2].f.spare[3] );
tran (\sa_ctrl_rst_dat[2][9] , \sa_ctrl_rst_dat[2].r.part0[9] );
tran (\sa_ctrl_rst_dat[2][9] , \sa_ctrl_rst_dat[2].f.spare[4] );
tran (\sa_ctrl_rst_dat[2][10] , \sa_ctrl_rst_dat[2].r.part0[10] );
tran (\sa_ctrl_rst_dat[2][10] , \sa_ctrl_rst_dat[2].f.spare[5] );
tran (\sa_ctrl_rst_dat[2][11] , \sa_ctrl_rst_dat[2].r.part0[11] );
tran (\sa_ctrl_rst_dat[2][11] , \sa_ctrl_rst_dat[2].f.spare[6] );
tran (\sa_ctrl_rst_dat[2][12] , \sa_ctrl_rst_dat[2].r.part0[12] );
tran (\sa_ctrl_rst_dat[2][12] , \sa_ctrl_rst_dat[2].f.spare[7] );
tran (\sa_ctrl_rst_dat[2][13] , \sa_ctrl_rst_dat[2].r.part0[13] );
tran (\sa_ctrl_rst_dat[2][13] , \sa_ctrl_rst_dat[2].f.spare[8] );
tran (\sa_ctrl_rst_dat[2][14] , \sa_ctrl_rst_dat[2].r.part0[14] );
tran (\sa_ctrl_rst_dat[2][14] , \sa_ctrl_rst_dat[2].f.spare[9] );
tran (\sa_ctrl_rst_dat[2][15] , \sa_ctrl_rst_dat[2].r.part0[15] );
tran (\sa_ctrl_rst_dat[2][15] , \sa_ctrl_rst_dat[2].f.spare[10] );
tran (\sa_ctrl_rst_dat[2][16] , \sa_ctrl_rst_dat[2].r.part0[16] );
tran (\sa_ctrl_rst_dat[2][16] , \sa_ctrl_rst_dat[2].f.spare[11] );
tran (\sa_ctrl_rst_dat[2][17] , \sa_ctrl_rst_dat[2].r.part0[17] );
tran (\sa_ctrl_rst_dat[2][17] , \sa_ctrl_rst_dat[2].f.spare[12] );
tran (\sa_ctrl_rst_dat[2][18] , \sa_ctrl_rst_dat[2].r.part0[18] );
tran (\sa_ctrl_rst_dat[2][18] , \sa_ctrl_rst_dat[2].f.spare[13] );
tran (\sa_ctrl_rst_dat[2][19] , \sa_ctrl_rst_dat[2].r.part0[19] );
tran (\sa_ctrl_rst_dat[2][19] , \sa_ctrl_rst_dat[2].f.spare[14] );
tran (\sa_ctrl_rst_dat[2][20] , \sa_ctrl_rst_dat[2].r.part0[20] );
tran (\sa_ctrl_rst_dat[2][20] , \sa_ctrl_rst_dat[2].f.spare[15] );
tran (\sa_ctrl_rst_dat[2][21] , \sa_ctrl_rst_dat[2].r.part0[21] );
tran (\sa_ctrl_rst_dat[2][21] , \sa_ctrl_rst_dat[2].f.spare[16] );
tran (\sa_ctrl_rst_dat[2][22] , \sa_ctrl_rst_dat[2].r.part0[22] );
tran (\sa_ctrl_rst_dat[2][22] , \sa_ctrl_rst_dat[2].f.spare[17] );
tran (\sa_ctrl_rst_dat[2][23] , \sa_ctrl_rst_dat[2].r.part0[23] );
tran (\sa_ctrl_rst_dat[2][23] , \sa_ctrl_rst_dat[2].f.spare[18] );
tran (\sa_ctrl_rst_dat[2][24] , \sa_ctrl_rst_dat[2].r.part0[24] );
tran (\sa_ctrl_rst_dat[2][24] , \sa_ctrl_rst_dat[2].f.spare[19] );
tran (\sa_ctrl_rst_dat[2][25] , \sa_ctrl_rst_dat[2].r.part0[25] );
tran (\sa_ctrl_rst_dat[2][25] , \sa_ctrl_rst_dat[2].f.spare[20] );
tran (\sa_ctrl_rst_dat[2][26] , \sa_ctrl_rst_dat[2].r.part0[26] );
tran (\sa_ctrl_rst_dat[2][26] , \sa_ctrl_rst_dat[2].f.spare[21] );
tran (\sa_ctrl_rst_dat[2][27] , \sa_ctrl_rst_dat[2].r.part0[27] );
tran (\sa_ctrl_rst_dat[2][27] , \sa_ctrl_rst_dat[2].f.spare[22] );
tran (\sa_ctrl_rst_dat[2][28] , \sa_ctrl_rst_dat[2].r.part0[28] );
tran (\sa_ctrl_rst_dat[2][28] , \sa_ctrl_rst_dat[2].f.spare[23] );
tran (\sa_ctrl_rst_dat[2][29] , \sa_ctrl_rst_dat[2].r.part0[29] );
tran (\sa_ctrl_rst_dat[2][29] , \sa_ctrl_rst_dat[2].f.spare[24] );
tran (\sa_ctrl_rst_dat[2][30] , \sa_ctrl_rst_dat[2].r.part0[30] );
tran (\sa_ctrl_rst_dat[2][30] , \sa_ctrl_rst_dat[2].f.spare[25] );
tran (\sa_ctrl_rst_dat[2][31] , \sa_ctrl_rst_dat[2].r.part0[31] );
tran (\sa_ctrl_rst_dat[2][31] , \sa_ctrl_rst_dat[2].f.spare[26] );
tran (\sa_ctrl_rst_dat[3][0] , \sa_ctrl_rst_dat[3].r.part0[0] );
tran (\sa_ctrl_rst_dat[3][0] , \sa_ctrl_rst_dat[3].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[3][1] , \sa_ctrl_rst_dat[3].r.part0[1] );
tran (\sa_ctrl_rst_dat[3][1] , \sa_ctrl_rst_dat[3].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[3][2] , \sa_ctrl_rst_dat[3].r.part0[2] );
tran (\sa_ctrl_rst_dat[3][2] , \sa_ctrl_rst_dat[3].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[3][3] , \sa_ctrl_rst_dat[3].r.part0[3] );
tran (\sa_ctrl_rst_dat[3][3] , \sa_ctrl_rst_dat[3].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[3][4] , \sa_ctrl_rst_dat[3].r.part0[4] );
tran (\sa_ctrl_rst_dat[3][4] , \sa_ctrl_rst_dat[3].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[3][5] , \sa_ctrl_rst_dat[3].r.part0[5] );
tran (\sa_ctrl_rst_dat[3][5] , \sa_ctrl_rst_dat[3].f.spare[0] );
tran (\sa_ctrl_rst_dat[3][6] , \sa_ctrl_rst_dat[3].r.part0[6] );
tran (\sa_ctrl_rst_dat[3][6] , \sa_ctrl_rst_dat[3].f.spare[1] );
tran (\sa_ctrl_rst_dat[3][7] , \sa_ctrl_rst_dat[3].r.part0[7] );
tran (\sa_ctrl_rst_dat[3][7] , \sa_ctrl_rst_dat[3].f.spare[2] );
tran (\sa_ctrl_rst_dat[3][8] , \sa_ctrl_rst_dat[3].r.part0[8] );
tran (\sa_ctrl_rst_dat[3][8] , \sa_ctrl_rst_dat[3].f.spare[3] );
tran (\sa_ctrl_rst_dat[3][9] , \sa_ctrl_rst_dat[3].r.part0[9] );
tran (\sa_ctrl_rst_dat[3][9] , \sa_ctrl_rst_dat[3].f.spare[4] );
tran (\sa_ctrl_rst_dat[3][10] , \sa_ctrl_rst_dat[3].r.part0[10] );
tran (\sa_ctrl_rst_dat[3][10] , \sa_ctrl_rst_dat[3].f.spare[5] );
tran (\sa_ctrl_rst_dat[3][11] , \sa_ctrl_rst_dat[3].r.part0[11] );
tran (\sa_ctrl_rst_dat[3][11] , \sa_ctrl_rst_dat[3].f.spare[6] );
tran (\sa_ctrl_rst_dat[3][12] , \sa_ctrl_rst_dat[3].r.part0[12] );
tran (\sa_ctrl_rst_dat[3][12] , \sa_ctrl_rst_dat[3].f.spare[7] );
tran (\sa_ctrl_rst_dat[3][13] , \sa_ctrl_rst_dat[3].r.part0[13] );
tran (\sa_ctrl_rst_dat[3][13] , \sa_ctrl_rst_dat[3].f.spare[8] );
tran (\sa_ctrl_rst_dat[3][14] , \sa_ctrl_rst_dat[3].r.part0[14] );
tran (\sa_ctrl_rst_dat[3][14] , \sa_ctrl_rst_dat[3].f.spare[9] );
tran (\sa_ctrl_rst_dat[3][15] , \sa_ctrl_rst_dat[3].r.part0[15] );
tran (\sa_ctrl_rst_dat[3][15] , \sa_ctrl_rst_dat[3].f.spare[10] );
tran (\sa_ctrl_rst_dat[3][16] , \sa_ctrl_rst_dat[3].r.part0[16] );
tran (\sa_ctrl_rst_dat[3][16] , \sa_ctrl_rst_dat[3].f.spare[11] );
tran (\sa_ctrl_rst_dat[3][17] , \sa_ctrl_rst_dat[3].r.part0[17] );
tran (\sa_ctrl_rst_dat[3][17] , \sa_ctrl_rst_dat[3].f.spare[12] );
tran (\sa_ctrl_rst_dat[3][18] , \sa_ctrl_rst_dat[3].r.part0[18] );
tran (\sa_ctrl_rst_dat[3][18] , \sa_ctrl_rst_dat[3].f.spare[13] );
tran (\sa_ctrl_rst_dat[3][19] , \sa_ctrl_rst_dat[3].r.part0[19] );
tran (\sa_ctrl_rst_dat[3][19] , \sa_ctrl_rst_dat[3].f.spare[14] );
tran (\sa_ctrl_rst_dat[3][20] , \sa_ctrl_rst_dat[3].r.part0[20] );
tran (\sa_ctrl_rst_dat[3][20] , \sa_ctrl_rst_dat[3].f.spare[15] );
tran (\sa_ctrl_rst_dat[3][21] , \sa_ctrl_rst_dat[3].r.part0[21] );
tran (\sa_ctrl_rst_dat[3][21] , \sa_ctrl_rst_dat[3].f.spare[16] );
tran (\sa_ctrl_rst_dat[3][22] , \sa_ctrl_rst_dat[3].r.part0[22] );
tran (\sa_ctrl_rst_dat[3][22] , \sa_ctrl_rst_dat[3].f.spare[17] );
tran (\sa_ctrl_rst_dat[3][23] , \sa_ctrl_rst_dat[3].r.part0[23] );
tran (\sa_ctrl_rst_dat[3][23] , \sa_ctrl_rst_dat[3].f.spare[18] );
tran (\sa_ctrl_rst_dat[3][24] , \sa_ctrl_rst_dat[3].r.part0[24] );
tran (\sa_ctrl_rst_dat[3][24] , \sa_ctrl_rst_dat[3].f.spare[19] );
tran (\sa_ctrl_rst_dat[3][25] , \sa_ctrl_rst_dat[3].r.part0[25] );
tran (\sa_ctrl_rst_dat[3][25] , \sa_ctrl_rst_dat[3].f.spare[20] );
tran (\sa_ctrl_rst_dat[3][26] , \sa_ctrl_rst_dat[3].r.part0[26] );
tran (\sa_ctrl_rst_dat[3][26] , \sa_ctrl_rst_dat[3].f.spare[21] );
tran (\sa_ctrl_rst_dat[3][27] , \sa_ctrl_rst_dat[3].r.part0[27] );
tran (\sa_ctrl_rst_dat[3][27] , \sa_ctrl_rst_dat[3].f.spare[22] );
tran (\sa_ctrl_rst_dat[3][28] , \sa_ctrl_rst_dat[3].r.part0[28] );
tran (\sa_ctrl_rst_dat[3][28] , \sa_ctrl_rst_dat[3].f.spare[23] );
tran (\sa_ctrl_rst_dat[3][29] , \sa_ctrl_rst_dat[3].r.part0[29] );
tran (\sa_ctrl_rst_dat[3][29] , \sa_ctrl_rst_dat[3].f.spare[24] );
tran (\sa_ctrl_rst_dat[3][30] , \sa_ctrl_rst_dat[3].r.part0[30] );
tran (\sa_ctrl_rst_dat[3][30] , \sa_ctrl_rst_dat[3].f.spare[25] );
tran (\sa_ctrl_rst_dat[3][31] , \sa_ctrl_rst_dat[3].r.part0[31] );
tran (\sa_ctrl_rst_dat[3][31] , \sa_ctrl_rst_dat[3].f.spare[26] );
tran (\sa_ctrl_rst_dat[4][0] , \sa_ctrl_rst_dat[4].r.part0[0] );
tran (\sa_ctrl_rst_dat[4][0] , \sa_ctrl_rst_dat[4].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[4][1] , \sa_ctrl_rst_dat[4].r.part0[1] );
tran (\sa_ctrl_rst_dat[4][1] , \sa_ctrl_rst_dat[4].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[4][2] , \sa_ctrl_rst_dat[4].r.part0[2] );
tran (\sa_ctrl_rst_dat[4][2] , \sa_ctrl_rst_dat[4].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[4][3] , \sa_ctrl_rst_dat[4].r.part0[3] );
tran (\sa_ctrl_rst_dat[4][3] , \sa_ctrl_rst_dat[4].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[4][4] , \sa_ctrl_rst_dat[4].r.part0[4] );
tran (\sa_ctrl_rst_dat[4][4] , \sa_ctrl_rst_dat[4].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[4][5] , \sa_ctrl_rst_dat[4].r.part0[5] );
tran (\sa_ctrl_rst_dat[4][5] , \sa_ctrl_rst_dat[4].f.spare[0] );
tran (\sa_ctrl_rst_dat[4][6] , \sa_ctrl_rst_dat[4].r.part0[6] );
tran (\sa_ctrl_rst_dat[4][6] , \sa_ctrl_rst_dat[4].f.spare[1] );
tran (\sa_ctrl_rst_dat[4][7] , \sa_ctrl_rst_dat[4].r.part0[7] );
tran (\sa_ctrl_rst_dat[4][7] , \sa_ctrl_rst_dat[4].f.spare[2] );
tran (\sa_ctrl_rst_dat[4][8] , \sa_ctrl_rst_dat[4].r.part0[8] );
tran (\sa_ctrl_rst_dat[4][8] , \sa_ctrl_rst_dat[4].f.spare[3] );
tran (\sa_ctrl_rst_dat[4][9] , \sa_ctrl_rst_dat[4].r.part0[9] );
tran (\sa_ctrl_rst_dat[4][9] , \sa_ctrl_rst_dat[4].f.spare[4] );
tran (\sa_ctrl_rst_dat[4][10] , \sa_ctrl_rst_dat[4].r.part0[10] );
tran (\sa_ctrl_rst_dat[4][10] , \sa_ctrl_rst_dat[4].f.spare[5] );
tran (\sa_ctrl_rst_dat[4][11] , \sa_ctrl_rst_dat[4].r.part0[11] );
tran (\sa_ctrl_rst_dat[4][11] , \sa_ctrl_rst_dat[4].f.spare[6] );
tran (\sa_ctrl_rst_dat[4][12] , \sa_ctrl_rst_dat[4].r.part0[12] );
tran (\sa_ctrl_rst_dat[4][12] , \sa_ctrl_rst_dat[4].f.spare[7] );
tran (\sa_ctrl_rst_dat[4][13] , \sa_ctrl_rst_dat[4].r.part0[13] );
tran (\sa_ctrl_rst_dat[4][13] , \sa_ctrl_rst_dat[4].f.spare[8] );
tran (\sa_ctrl_rst_dat[4][14] , \sa_ctrl_rst_dat[4].r.part0[14] );
tran (\sa_ctrl_rst_dat[4][14] , \sa_ctrl_rst_dat[4].f.spare[9] );
tran (\sa_ctrl_rst_dat[4][15] , \sa_ctrl_rst_dat[4].r.part0[15] );
tran (\sa_ctrl_rst_dat[4][15] , \sa_ctrl_rst_dat[4].f.spare[10] );
tran (\sa_ctrl_rst_dat[4][16] , \sa_ctrl_rst_dat[4].r.part0[16] );
tran (\sa_ctrl_rst_dat[4][16] , \sa_ctrl_rst_dat[4].f.spare[11] );
tran (\sa_ctrl_rst_dat[4][17] , \sa_ctrl_rst_dat[4].r.part0[17] );
tran (\sa_ctrl_rst_dat[4][17] , \sa_ctrl_rst_dat[4].f.spare[12] );
tran (\sa_ctrl_rst_dat[4][18] , \sa_ctrl_rst_dat[4].r.part0[18] );
tran (\sa_ctrl_rst_dat[4][18] , \sa_ctrl_rst_dat[4].f.spare[13] );
tran (\sa_ctrl_rst_dat[4][19] , \sa_ctrl_rst_dat[4].r.part0[19] );
tran (\sa_ctrl_rst_dat[4][19] , \sa_ctrl_rst_dat[4].f.spare[14] );
tran (\sa_ctrl_rst_dat[4][20] , \sa_ctrl_rst_dat[4].r.part0[20] );
tran (\sa_ctrl_rst_dat[4][20] , \sa_ctrl_rst_dat[4].f.spare[15] );
tran (\sa_ctrl_rst_dat[4][21] , \sa_ctrl_rst_dat[4].r.part0[21] );
tran (\sa_ctrl_rst_dat[4][21] , \sa_ctrl_rst_dat[4].f.spare[16] );
tran (\sa_ctrl_rst_dat[4][22] , \sa_ctrl_rst_dat[4].r.part0[22] );
tran (\sa_ctrl_rst_dat[4][22] , \sa_ctrl_rst_dat[4].f.spare[17] );
tran (\sa_ctrl_rst_dat[4][23] , \sa_ctrl_rst_dat[4].r.part0[23] );
tran (\sa_ctrl_rst_dat[4][23] , \sa_ctrl_rst_dat[4].f.spare[18] );
tran (\sa_ctrl_rst_dat[4][24] , \sa_ctrl_rst_dat[4].r.part0[24] );
tran (\sa_ctrl_rst_dat[4][24] , \sa_ctrl_rst_dat[4].f.spare[19] );
tran (\sa_ctrl_rst_dat[4][25] , \sa_ctrl_rst_dat[4].r.part0[25] );
tran (\sa_ctrl_rst_dat[4][25] , \sa_ctrl_rst_dat[4].f.spare[20] );
tran (\sa_ctrl_rst_dat[4][26] , \sa_ctrl_rst_dat[4].r.part0[26] );
tran (\sa_ctrl_rst_dat[4][26] , \sa_ctrl_rst_dat[4].f.spare[21] );
tran (\sa_ctrl_rst_dat[4][27] , \sa_ctrl_rst_dat[4].r.part0[27] );
tran (\sa_ctrl_rst_dat[4][27] , \sa_ctrl_rst_dat[4].f.spare[22] );
tran (\sa_ctrl_rst_dat[4][28] , \sa_ctrl_rst_dat[4].r.part0[28] );
tran (\sa_ctrl_rst_dat[4][28] , \sa_ctrl_rst_dat[4].f.spare[23] );
tran (\sa_ctrl_rst_dat[4][29] , \sa_ctrl_rst_dat[4].r.part0[29] );
tran (\sa_ctrl_rst_dat[4][29] , \sa_ctrl_rst_dat[4].f.spare[24] );
tran (\sa_ctrl_rst_dat[4][30] , \sa_ctrl_rst_dat[4].r.part0[30] );
tran (\sa_ctrl_rst_dat[4][30] , \sa_ctrl_rst_dat[4].f.spare[25] );
tran (\sa_ctrl_rst_dat[4][31] , \sa_ctrl_rst_dat[4].r.part0[31] );
tran (\sa_ctrl_rst_dat[4][31] , \sa_ctrl_rst_dat[4].f.spare[26] );
tran (\sa_ctrl_rst_dat[5][0] , \sa_ctrl_rst_dat[5].r.part0[0] );
tran (\sa_ctrl_rst_dat[5][0] , \sa_ctrl_rst_dat[5].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[5][1] , \sa_ctrl_rst_dat[5].r.part0[1] );
tran (\sa_ctrl_rst_dat[5][1] , \sa_ctrl_rst_dat[5].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[5][2] , \sa_ctrl_rst_dat[5].r.part0[2] );
tran (\sa_ctrl_rst_dat[5][2] , \sa_ctrl_rst_dat[5].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[5][3] , \sa_ctrl_rst_dat[5].r.part0[3] );
tran (\sa_ctrl_rst_dat[5][3] , \sa_ctrl_rst_dat[5].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[5][4] , \sa_ctrl_rst_dat[5].r.part0[4] );
tran (\sa_ctrl_rst_dat[5][4] , \sa_ctrl_rst_dat[5].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[5][5] , \sa_ctrl_rst_dat[5].r.part0[5] );
tran (\sa_ctrl_rst_dat[5][5] , \sa_ctrl_rst_dat[5].f.spare[0] );
tran (\sa_ctrl_rst_dat[5][6] , \sa_ctrl_rst_dat[5].r.part0[6] );
tran (\sa_ctrl_rst_dat[5][6] , \sa_ctrl_rst_dat[5].f.spare[1] );
tran (\sa_ctrl_rst_dat[5][7] , \sa_ctrl_rst_dat[5].r.part0[7] );
tran (\sa_ctrl_rst_dat[5][7] , \sa_ctrl_rst_dat[5].f.spare[2] );
tran (\sa_ctrl_rst_dat[5][8] , \sa_ctrl_rst_dat[5].r.part0[8] );
tran (\sa_ctrl_rst_dat[5][8] , \sa_ctrl_rst_dat[5].f.spare[3] );
tran (\sa_ctrl_rst_dat[5][9] , \sa_ctrl_rst_dat[5].r.part0[9] );
tran (\sa_ctrl_rst_dat[5][9] , \sa_ctrl_rst_dat[5].f.spare[4] );
tran (\sa_ctrl_rst_dat[5][10] , \sa_ctrl_rst_dat[5].r.part0[10] );
tran (\sa_ctrl_rst_dat[5][10] , \sa_ctrl_rst_dat[5].f.spare[5] );
tran (\sa_ctrl_rst_dat[5][11] , \sa_ctrl_rst_dat[5].r.part0[11] );
tran (\sa_ctrl_rst_dat[5][11] , \sa_ctrl_rst_dat[5].f.spare[6] );
tran (\sa_ctrl_rst_dat[5][12] , \sa_ctrl_rst_dat[5].r.part0[12] );
tran (\sa_ctrl_rst_dat[5][12] , \sa_ctrl_rst_dat[5].f.spare[7] );
tran (\sa_ctrl_rst_dat[5][13] , \sa_ctrl_rst_dat[5].r.part0[13] );
tran (\sa_ctrl_rst_dat[5][13] , \sa_ctrl_rst_dat[5].f.spare[8] );
tran (\sa_ctrl_rst_dat[5][14] , \sa_ctrl_rst_dat[5].r.part0[14] );
tran (\sa_ctrl_rst_dat[5][14] , \sa_ctrl_rst_dat[5].f.spare[9] );
tran (\sa_ctrl_rst_dat[5][15] , \sa_ctrl_rst_dat[5].r.part0[15] );
tran (\sa_ctrl_rst_dat[5][15] , \sa_ctrl_rst_dat[5].f.spare[10] );
tran (\sa_ctrl_rst_dat[5][16] , \sa_ctrl_rst_dat[5].r.part0[16] );
tran (\sa_ctrl_rst_dat[5][16] , \sa_ctrl_rst_dat[5].f.spare[11] );
tran (\sa_ctrl_rst_dat[5][17] , \sa_ctrl_rst_dat[5].r.part0[17] );
tran (\sa_ctrl_rst_dat[5][17] , \sa_ctrl_rst_dat[5].f.spare[12] );
tran (\sa_ctrl_rst_dat[5][18] , \sa_ctrl_rst_dat[5].r.part0[18] );
tran (\sa_ctrl_rst_dat[5][18] , \sa_ctrl_rst_dat[5].f.spare[13] );
tran (\sa_ctrl_rst_dat[5][19] , \sa_ctrl_rst_dat[5].r.part0[19] );
tran (\sa_ctrl_rst_dat[5][19] , \sa_ctrl_rst_dat[5].f.spare[14] );
tran (\sa_ctrl_rst_dat[5][20] , \sa_ctrl_rst_dat[5].r.part0[20] );
tran (\sa_ctrl_rst_dat[5][20] , \sa_ctrl_rst_dat[5].f.spare[15] );
tran (\sa_ctrl_rst_dat[5][21] , \sa_ctrl_rst_dat[5].r.part0[21] );
tran (\sa_ctrl_rst_dat[5][21] , \sa_ctrl_rst_dat[5].f.spare[16] );
tran (\sa_ctrl_rst_dat[5][22] , \sa_ctrl_rst_dat[5].r.part0[22] );
tran (\sa_ctrl_rst_dat[5][22] , \sa_ctrl_rst_dat[5].f.spare[17] );
tran (\sa_ctrl_rst_dat[5][23] , \sa_ctrl_rst_dat[5].r.part0[23] );
tran (\sa_ctrl_rst_dat[5][23] , \sa_ctrl_rst_dat[5].f.spare[18] );
tran (\sa_ctrl_rst_dat[5][24] , \sa_ctrl_rst_dat[5].r.part0[24] );
tran (\sa_ctrl_rst_dat[5][24] , \sa_ctrl_rst_dat[5].f.spare[19] );
tran (\sa_ctrl_rst_dat[5][25] , \sa_ctrl_rst_dat[5].r.part0[25] );
tran (\sa_ctrl_rst_dat[5][25] , \sa_ctrl_rst_dat[5].f.spare[20] );
tran (\sa_ctrl_rst_dat[5][26] , \sa_ctrl_rst_dat[5].r.part0[26] );
tran (\sa_ctrl_rst_dat[5][26] , \sa_ctrl_rst_dat[5].f.spare[21] );
tran (\sa_ctrl_rst_dat[5][27] , \sa_ctrl_rst_dat[5].r.part0[27] );
tran (\sa_ctrl_rst_dat[5][27] , \sa_ctrl_rst_dat[5].f.spare[22] );
tran (\sa_ctrl_rst_dat[5][28] , \sa_ctrl_rst_dat[5].r.part0[28] );
tran (\sa_ctrl_rst_dat[5][28] , \sa_ctrl_rst_dat[5].f.spare[23] );
tran (\sa_ctrl_rst_dat[5][29] , \sa_ctrl_rst_dat[5].r.part0[29] );
tran (\sa_ctrl_rst_dat[5][29] , \sa_ctrl_rst_dat[5].f.spare[24] );
tran (\sa_ctrl_rst_dat[5][30] , \sa_ctrl_rst_dat[5].r.part0[30] );
tran (\sa_ctrl_rst_dat[5][30] , \sa_ctrl_rst_dat[5].f.spare[25] );
tran (\sa_ctrl_rst_dat[5][31] , \sa_ctrl_rst_dat[5].r.part0[31] );
tran (\sa_ctrl_rst_dat[5][31] , \sa_ctrl_rst_dat[5].f.spare[26] );
tran (\sa_ctrl_rst_dat[6][0] , \sa_ctrl_rst_dat[6].r.part0[0] );
tran (\sa_ctrl_rst_dat[6][0] , \sa_ctrl_rst_dat[6].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[6][1] , \sa_ctrl_rst_dat[6].r.part0[1] );
tran (\sa_ctrl_rst_dat[6][1] , \sa_ctrl_rst_dat[6].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[6][2] , \sa_ctrl_rst_dat[6].r.part0[2] );
tran (\sa_ctrl_rst_dat[6][2] , \sa_ctrl_rst_dat[6].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[6][3] , \sa_ctrl_rst_dat[6].r.part0[3] );
tran (\sa_ctrl_rst_dat[6][3] , \sa_ctrl_rst_dat[6].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[6][4] , \sa_ctrl_rst_dat[6].r.part0[4] );
tran (\sa_ctrl_rst_dat[6][4] , \sa_ctrl_rst_dat[6].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[6][5] , \sa_ctrl_rst_dat[6].r.part0[5] );
tran (\sa_ctrl_rst_dat[6][5] , \sa_ctrl_rst_dat[6].f.spare[0] );
tran (\sa_ctrl_rst_dat[6][6] , \sa_ctrl_rst_dat[6].r.part0[6] );
tran (\sa_ctrl_rst_dat[6][6] , \sa_ctrl_rst_dat[6].f.spare[1] );
tran (\sa_ctrl_rst_dat[6][7] , \sa_ctrl_rst_dat[6].r.part0[7] );
tran (\sa_ctrl_rst_dat[6][7] , \sa_ctrl_rst_dat[6].f.spare[2] );
tran (\sa_ctrl_rst_dat[6][8] , \sa_ctrl_rst_dat[6].r.part0[8] );
tran (\sa_ctrl_rst_dat[6][8] , \sa_ctrl_rst_dat[6].f.spare[3] );
tran (\sa_ctrl_rst_dat[6][9] , \sa_ctrl_rst_dat[6].r.part0[9] );
tran (\sa_ctrl_rst_dat[6][9] , \sa_ctrl_rst_dat[6].f.spare[4] );
tran (\sa_ctrl_rst_dat[6][10] , \sa_ctrl_rst_dat[6].r.part0[10] );
tran (\sa_ctrl_rst_dat[6][10] , \sa_ctrl_rst_dat[6].f.spare[5] );
tran (\sa_ctrl_rst_dat[6][11] , \sa_ctrl_rst_dat[6].r.part0[11] );
tran (\sa_ctrl_rst_dat[6][11] , \sa_ctrl_rst_dat[6].f.spare[6] );
tran (\sa_ctrl_rst_dat[6][12] , \sa_ctrl_rst_dat[6].r.part0[12] );
tran (\sa_ctrl_rst_dat[6][12] , \sa_ctrl_rst_dat[6].f.spare[7] );
tran (\sa_ctrl_rst_dat[6][13] , \sa_ctrl_rst_dat[6].r.part0[13] );
tran (\sa_ctrl_rst_dat[6][13] , \sa_ctrl_rst_dat[6].f.spare[8] );
tran (\sa_ctrl_rst_dat[6][14] , \sa_ctrl_rst_dat[6].r.part0[14] );
tran (\sa_ctrl_rst_dat[6][14] , \sa_ctrl_rst_dat[6].f.spare[9] );
tran (\sa_ctrl_rst_dat[6][15] , \sa_ctrl_rst_dat[6].r.part0[15] );
tran (\sa_ctrl_rst_dat[6][15] , \sa_ctrl_rst_dat[6].f.spare[10] );
tran (\sa_ctrl_rst_dat[6][16] , \sa_ctrl_rst_dat[6].r.part0[16] );
tran (\sa_ctrl_rst_dat[6][16] , \sa_ctrl_rst_dat[6].f.spare[11] );
tran (\sa_ctrl_rst_dat[6][17] , \sa_ctrl_rst_dat[6].r.part0[17] );
tran (\sa_ctrl_rst_dat[6][17] , \sa_ctrl_rst_dat[6].f.spare[12] );
tran (\sa_ctrl_rst_dat[6][18] , \sa_ctrl_rst_dat[6].r.part0[18] );
tran (\sa_ctrl_rst_dat[6][18] , \sa_ctrl_rst_dat[6].f.spare[13] );
tran (\sa_ctrl_rst_dat[6][19] , \sa_ctrl_rst_dat[6].r.part0[19] );
tran (\sa_ctrl_rst_dat[6][19] , \sa_ctrl_rst_dat[6].f.spare[14] );
tran (\sa_ctrl_rst_dat[6][20] , \sa_ctrl_rst_dat[6].r.part0[20] );
tran (\sa_ctrl_rst_dat[6][20] , \sa_ctrl_rst_dat[6].f.spare[15] );
tran (\sa_ctrl_rst_dat[6][21] , \sa_ctrl_rst_dat[6].r.part0[21] );
tran (\sa_ctrl_rst_dat[6][21] , \sa_ctrl_rst_dat[6].f.spare[16] );
tran (\sa_ctrl_rst_dat[6][22] , \sa_ctrl_rst_dat[6].r.part0[22] );
tran (\sa_ctrl_rst_dat[6][22] , \sa_ctrl_rst_dat[6].f.spare[17] );
tran (\sa_ctrl_rst_dat[6][23] , \sa_ctrl_rst_dat[6].r.part0[23] );
tran (\sa_ctrl_rst_dat[6][23] , \sa_ctrl_rst_dat[6].f.spare[18] );
tran (\sa_ctrl_rst_dat[6][24] , \sa_ctrl_rst_dat[6].r.part0[24] );
tran (\sa_ctrl_rst_dat[6][24] , \sa_ctrl_rst_dat[6].f.spare[19] );
tran (\sa_ctrl_rst_dat[6][25] , \sa_ctrl_rst_dat[6].r.part0[25] );
tran (\sa_ctrl_rst_dat[6][25] , \sa_ctrl_rst_dat[6].f.spare[20] );
tran (\sa_ctrl_rst_dat[6][26] , \sa_ctrl_rst_dat[6].r.part0[26] );
tran (\sa_ctrl_rst_dat[6][26] , \sa_ctrl_rst_dat[6].f.spare[21] );
tran (\sa_ctrl_rst_dat[6][27] , \sa_ctrl_rst_dat[6].r.part0[27] );
tran (\sa_ctrl_rst_dat[6][27] , \sa_ctrl_rst_dat[6].f.spare[22] );
tran (\sa_ctrl_rst_dat[6][28] , \sa_ctrl_rst_dat[6].r.part0[28] );
tran (\sa_ctrl_rst_dat[6][28] , \sa_ctrl_rst_dat[6].f.spare[23] );
tran (\sa_ctrl_rst_dat[6][29] , \sa_ctrl_rst_dat[6].r.part0[29] );
tran (\sa_ctrl_rst_dat[6][29] , \sa_ctrl_rst_dat[6].f.spare[24] );
tran (\sa_ctrl_rst_dat[6][30] , \sa_ctrl_rst_dat[6].r.part0[30] );
tran (\sa_ctrl_rst_dat[6][30] , \sa_ctrl_rst_dat[6].f.spare[25] );
tran (\sa_ctrl_rst_dat[6][31] , \sa_ctrl_rst_dat[6].r.part0[31] );
tran (\sa_ctrl_rst_dat[6][31] , \sa_ctrl_rst_dat[6].f.spare[26] );
tran (\sa_ctrl_rst_dat[7][0] , \sa_ctrl_rst_dat[7].r.part0[0] );
tran (\sa_ctrl_rst_dat[7][0] , \sa_ctrl_rst_dat[7].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[7][1] , \sa_ctrl_rst_dat[7].r.part0[1] );
tran (\sa_ctrl_rst_dat[7][1] , \sa_ctrl_rst_dat[7].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[7][2] , \sa_ctrl_rst_dat[7].r.part0[2] );
tran (\sa_ctrl_rst_dat[7][2] , \sa_ctrl_rst_dat[7].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[7][3] , \sa_ctrl_rst_dat[7].r.part0[3] );
tran (\sa_ctrl_rst_dat[7][3] , \sa_ctrl_rst_dat[7].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[7][4] , \sa_ctrl_rst_dat[7].r.part0[4] );
tran (\sa_ctrl_rst_dat[7][4] , \sa_ctrl_rst_dat[7].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[7][5] , \sa_ctrl_rst_dat[7].r.part0[5] );
tran (\sa_ctrl_rst_dat[7][5] , \sa_ctrl_rst_dat[7].f.spare[0] );
tran (\sa_ctrl_rst_dat[7][6] , \sa_ctrl_rst_dat[7].r.part0[6] );
tran (\sa_ctrl_rst_dat[7][6] , \sa_ctrl_rst_dat[7].f.spare[1] );
tran (\sa_ctrl_rst_dat[7][7] , \sa_ctrl_rst_dat[7].r.part0[7] );
tran (\sa_ctrl_rst_dat[7][7] , \sa_ctrl_rst_dat[7].f.spare[2] );
tran (\sa_ctrl_rst_dat[7][8] , \sa_ctrl_rst_dat[7].r.part0[8] );
tran (\sa_ctrl_rst_dat[7][8] , \sa_ctrl_rst_dat[7].f.spare[3] );
tran (\sa_ctrl_rst_dat[7][9] , \sa_ctrl_rst_dat[7].r.part0[9] );
tran (\sa_ctrl_rst_dat[7][9] , \sa_ctrl_rst_dat[7].f.spare[4] );
tran (\sa_ctrl_rst_dat[7][10] , \sa_ctrl_rst_dat[7].r.part0[10] );
tran (\sa_ctrl_rst_dat[7][10] , \sa_ctrl_rst_dat[7].f.spare[5] );
tran (\sa_ctrl_rst_dat[7][11] , \sa_ctrl_rst_dat[7].r.part0[11] );
tran (\sa_ctrl_rst_dat[7][11] , \sa_ctrl_rst_dat[7].f.spare[6] );
tran (\sa_ctrl_rst_dat[7][12] , \sa_ctrl_rst_dat[7].r.part0[12] );
tran (\sa_ctrl_rst_dat[7][12] , \sa_ctrl_rst_dat[7].f.spare[7] );
tran (\sa_ctrl_rst_dat[7][13] , \sa_ctrl_rst_dat[7].r.part0[13] );
tran (\sa_ctrl_rst_dat[7][13] , \sa_ctrl_rst_dat[7].f.spare[8] );
tran (\sa_ctrl_rst_dat[7][14] , \sa_ctrl_rst_dat[7].r.part0[14] );
tran (\sa_ctrl_rst_dat[7][14] , \sa_ctrl_rst_dat[7].f.spare[9] );
tran (\sa_ctrl_rst_dat[7][15] , \sa_ctrl_rst_dat[7].r.part0[15] );
tran (\sa_ctrl_rst_dat[7][15] , \sa_ctrl_rst_dat[7].f.spare[10] );
tran (\sa_ctrl_rst_dat[7][16] , \sa_ctrl_rst_dat[7].r.part0[16] );
tran (\sa_ctrl_rst_dat[7][16] , \sa_ctrl_rst_dat[7].f.spare[11] );
tran (\sa_ctrl_rst_dat[7][17] , \sa_ctrl_rst_dat[7].r.part0[17] );
tran (\sa_ctrl_rst_dat[7][17] , \sa_ctrl_rst_dat[7].f.spare[12] );
tran (\sa_ctrl_rst_dat[7][18] , \sa_ctrl_rst_dat[7].r.part0[18] );
tran (\sa_ctrl_rst_dat[7][18] , \sa_ctrl_rst_dat[7].f.spare[13] );
tran (\sa_ctrl_rst_dat[7][19] , \sa_ctrl_rst_dat[7].r.part0[19] );
tran (\sa_ctrl_rst_dat[7][19] , \sa_ctrl_rst_dat[7].f.spare[14] );
tran (\sa_ctrl_rst_dat[7][20] , \sa_ctrl_rst_dat[7].r.part0[20] );
tran (\sa_ctrl_rst_dat[7][20] , \sa_ctrl_rst_dat[7].f.spare[15] );
tran (\sa_ctrl_rst_dat[7][21] , \sa_ctrl_rst_dat[7].r.part0[21] );
tran (\sa_ctrl_rst_dat[7][21] , \sa_ctrl_rst_dat[7].f.spare[16] );
tran (\sa_ctrl_rst_dat[7][22] , \sa_ctrl_rst_dat[7].r.part0[22] );
tran (\sa_ctrl_rst_dat[7][22] , \sa_ctrl_rst_dat[7].f.spare[17] );
tran (\sa_ctrl_rst_dat[7][23] , \sa_ctrl_rst_dat[7].r.part0[23] );
tran (\sa_ctrl_rst_dat[7][23] , \sa_ctrl_rst_dat[7].f.spare[18] );
tran (\sa_ctrl_rst_dat[7][24] , \sa_ctrl_rst_dat[7].r.part0[24] );
tran (\sa_ctrl_rst_dat[7][24] , \sa_ctrl_rst_dat[7].f.spare[19] );
tran (\sa_ctrl_rst_dat[7][25] , \sa_ctrl_rst_dat[7].r.part0[25] );
tran (\sa_ctrl_rst_dat[7][25] , \sa_ctrl_rst_dat[7].f.spare[20] );
tran (\sa_ctrl_rst_dat[7][26] , \sa_ctrl_rst_dat[7].r.part0[26] );
tran (\sa_ctrl_rst_dat[7][26] , \sa_ctrl_rst_dat[7].f.spare[21] );
tran (\sa_ctrl_rst_dat[7][27] , \sa_ctrl_rst_dat[7].r.part0[27] );
tran (\sa_ctrl_rst_dat[7][27] , \sa_ctrl_rst_dat[7].f.spare[22] );
tran (\sa_ctrl_rst_dat[7][28] , \sa_ctrl_rst_dat[7].r.part0[28] );
tran (\sa_ctrl_rst_dat[7][28] , \sa_ctrl_rst_dat[7].f.spare[23] );
tran (\sa_ctrl_rst_dat[7][29] , \sa_ctrl_rst_dat[7].r.part0[29] );
tran (\sa_ctrl_rst_dat[7][29] , \sa_ctrl_rst_dat[7].f.spare[24] );
tran (\sa_ctrl_rst_dat[7][30] , \sa_ctrl_rst_dat[7].r.part0[30] );
tran (\sa_ctrl_rst_dat[7][30] , \sa_ctrl_rst_dat[7].f.spare[25] );
tran (\sa_ctrl_rst_dat[7][31] , \sa_ctrl_rst_dat[7].r.part0[31] );
tran (\sa_ctrl_rst_dat[7][31] , \sa_ctrl_rst_dat[7].f.spare[26] );
tran (\sa_ctrl_rst_dat[8][0] , \sa_ctrl_rst_dat[8].r.part0[0] );
tran (\sa_ctrl_rst_dat[8][0] , \sa_ctrl_rst_dat[8].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[8][1] , \sa_ctrl_rst_dat[8].r.part0[1] );
tran (\sa_ctrl_rst_dat[8][1] , \sa_ctrl_rst_dat[8].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[8][2] , \sa_ctrl_rst_dat[8].r.part0[2] );
tran (\sa_ctrl_rst_dat[8][2] , \sa_ctrl_rst_dat[8].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[8][3] , \sa_ctrl_rst_dat[8].r.part0[3] );
tran (\sa_ctrl_rst_dat[8][3] , \sa_ctrl_rst_dat[8].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[8][4] , \sa_ctrl_rst_dat[8].r.part0[4] );
tran (\sa_ctrl_rst_dat[8][4] , \sa_ctrl_rst_dat[8].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[8][5] , \sa_ctrl_rst_dat[8].r.part0[5] );
tran (\sa_ctrl_rst_dat[8][5] , \sa_ctrl_rst_dat[8].f.spare[0] );
tran (\sa_ctrl_rst_dat[8][6] , \sa_ctrl_rst_dat[8].r.part0[6] );
tran (\sa_ctrl_rst_dat[8][6] , \sa_ctrl_rst_dat[8].f.spare[1] );
tran (\sa_ctrl_rst_dat[8][7] , \sa_ctrl_rst_dat[8].r.part0[7] );
tran (\sa_ctrl_rst_dat[8][7] , \sa_ctrl_rst_dat[8].f.spare[2] );
tran (\sa_ctrl_rst_dat[8][8] , \sa_ctrl_rst_dat[8].r.part0[8] );
tran (\sa_ctrl_rst_dat[8][8] , \sa_ctrl_rst_dat[8].f.spare[3] );
tran (\sa_ctrl_rst_dat[8][9] , \sa_ctrl_rst_dat[8].r.part0[9] );
tran (\sa_ctrl_rst_dat[8][9] , \sa_ctrl_rst_dat[8].f.spare[4] );
tran (\sa_ctrl_rst_dat[8][10] , \sa_ctrl_rst_dat[8].r.part0[10] );
tran (\sa_ctrl_rst_dat[8][10] , \sa_ctrl_rst_dat[8].f.spare[5] );
tran (\sa_ctrl_rst_dat[8][11] , \sa_ctrl_rst_dat[8].r.part0[11] );
tran (\sa_ctrl_rst_dat[8][11] , \sa_ctrl_rst_dat[8].f.spare[6] );
tran (\sa_ctrl_rst_dat[8][12] , \sa_ctrl_rst_dat[8].r.part0[12] );
tran (\sa_ctrl_rst_dat[8][12] , \sa_ctrl_rst_dat[8].f.spare[7] );
tran (\sa_ctrl_rst_dat[8][13] , \sa_ctrl_rst_dat[8].r.part0[13] );
tran (\sa_ctrl_rst_dat[8][13] , \sa_ctrl_rst_dat[8].f.spare[8] );
tran (\sa_ctrl_rst_dat[8][14] , \sa_ctrl_rst_dat[8].r.part0[14] );
tran (\sa_ctrl_rst_dat[8][14] , \sa_ctrl_rst_dat[8].f.spare[9] );
tran (\sa_ctrl_rst_dat[8][15] , \sa_ctrl_rst_dat[8].r.part0[15] );
tran (\sa_ctrl_rst_dat[8][15] , \sa_ctrl_rst_dat[8].f.spare[10] );
tran (\sa_ctrl_rst_dat[8][16] , \sa_ctrl_rst_dat[8].r.part0[16] );
tran (\sa_ctrl_rst_dat[8][16] , \sa_ctrl_rst_dat[8].f.spare[11] );
tran (\sa_ctrl_rst_dat[8][17] , \sa_ctrl_rst_dat[8].r.part0[17] );
tran (\sa_ctrl_rst_dat[8][17] , \sa_ctrl_rst_dat[8].f.spare[12] );
tran (\sa_ctrl_rst_dat[8][18] , \sa_ctrl_rst_dat[8].r.part0[18] );
tran (\sa_ctrl_rst_dat[8][18] , \sa_ctrl_rst_dat[8].f.spare[13] );
tran (\sa_ctrl_rst_dat[8][19] , \sa_ctrl_rst_dat[8].r.part0[19] );
tran (\sa_ctrl_rst_dat[8][19] , \sa_ctrl_rst_dat[8].f.spare[14] );
tran (\sa_ctrl_rst_dat[8][20] , \sa_ctrl_rst_dat[8].r.part0[20] );
tran (\sa_ctrl_rst_dat[8][20] , \sa_ctrl_rst_dat[8].f.spare[15] );
tran (\sa_ctrl_rst_dat[8][21] , \sa_ctrl_rst_dat[8].r.part0[21] );
tran (\sa_ctrl_rst_dat[8][21] , \sa_ctrl_rst_dat[8].f.spare[16] );
tran (\sa_ctrl_rst_dat[8][22] , \sa_ctrl_rst_dat[8].r.part0[22] );
tran (\sa_ctrl_rst_dat[8][22] , \sa_ctrl_rst_dat[8].f.spare[17] );
tran (\sa_ctrl_rst_dat[8][23] , \sa_ctrl_rst_dat[8].r.part0[23] );
tran (\sa_ctrl_rst_dat[8][23] , \sa_ctrl_rst_dat[8].f.spare[18] );
tran (\sa_ctrl_rst_dat[8][24] , \sa_ctrl_rst_dat[8].r.part0[24] );
tran (\sa_ctrl_rst_dat[8][24] , \sa_ctrl_rst_dat[8].f.spare[19] );
tran (\sa_ctrl_rst_dat[8][25] , \sa_ctrl_rst_dat[8].r.part0[25] );
tran (\sa_ctrl_rst_dat[8][25] , \sa_ctrl_rst_dat[8].f.spare[20] );
tran (\sa_ctrl_rst_dat[8][26] , \sa_ctrl_rst_dat[8].r.part0[26] );
tran (\sa_ctrl_rst_dat[8][26] , \sa_ctrl_rst_dat[8].f.spare[21] );
tran (\sa_ctrl_rst_dat[8][27] , \sa_ctrl_rst_dat[8].r.part0[27] );
tran (\sa_ctrl_rst_dat[8][27] , \sa_ctrl_rst_dat[8].f.spare[22] );
tran (\sa_ctrl_rst_dat[8][28] , \sa_ctrl_rst_dat[8].r.part0[28] );
tran (\sa_ctrl_rst_dat[8][28] , \sa_ctrl_rst_dat[8].f.spare[23] );
tran (\sa_ctrl_rst_dat[8][29] , \sa_ctrl_rst_dat[8].r.part0[29] );
tran (\sa_ctrl_rst_dat[8][29] , \sa_ctrl_rst_dat[8].f.spare[24] );
tran (\sa_ctrl_rst_dat[8][30] , \sa_ctrl_rst_dat[8].r.part0[30] );
tran (\sa_ctrl_rst_dat[8][30] , \sa_ctrl_rst_dat[8].f.spare[25] );
tran (\sa_ctrl_rst_dat[8][31] , \sa_ctrl_rst_dat[8].r.part0[31] );
tran (\sa_ctrl_rst_dat[8][31] , \sa_ctrl_rst_dat[8].f.spare[26] );
tran (\sa_ctrl_rst_dat[9][0] , \sa_ctrl_rst_dat[9].r.part0[0] );
tran (\sa_ctrl_rst_dat[9][0] , \sa_ctrl_rst_dat[9].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[9][1] , \sa_ctrl_rst_dat[9].r.part0[1] );
tran (\sa_ctrl_rst_dat[9][1] , \sa_ctrl_rst_dat[9].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[9][2] , \sa_ctrl_rst_dat[9].r.part0[2] );
tran (\sa_ctrl_rst_dat[9][2] , \sa_ctrl_rst_dat[9].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[9][3] , \sa_ctrl_rst_dat[9].r.part0[3] );
tran (\sa_ctrl_rst_dat[9][3] , \sa_ctrl_rst_dat[9].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[9][4] , \sa_ctrl_rst_dat[9].r.part0[4] );
tran (\sa_ctrl_rst_dat[9][4] , \sa_ctrl_rst_dat[9].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[9][5] , \sa_ctrl_rst_dat[9].r.part0[5] );
tran (\sa_ctrl_rst_dat[9][5] , \sa_ctrl_rst_dat[9].f.spare[0] );
tran (\sa_ctrl_rst_dat[9][6] , \sa_ctrl_rst_dat[9].r.part0[6] );
tran (\sa_ctrl_rst_dat[9][6] , \sa_ctrl_rst_dat[9].f.spare[1] );
tran (\sa_ctrl_rst_dat[9][7] , \sa_ctrl_rst_dat[9].r.part0[7] );
tran (\sa_ctrl_rst_dat[9][7] , \sa_ctrl_rst_dat[9].f.spare[2] );
tran (\sa_ctrl_rst_dat[9][8] , \sa_ctrl_rst_dat[9].r.part0[8] );
tran (\sa_ctrl_rst_dat[9][8] , \sa_ctrl_rst_dat[9].f.spare[3] );
tran (\sa_ctrl_rst_dat[9][9] , \sa_ctrl_rst_dat[9].r.part0[9] );
tran (\sa_ctrl_rst_dat[9][9] , \sa_ctrl_rst_dat[9].f.spare[4] );
tran (\sa_ctrl_rst_dat[9][10] , \sa_ctrl_rst_dat[9].r.part0[10] );
tran (\sa_ctrl_rst_dat[9][10] , \sa_ctrl_rst_dat[9].f.spare[5] );
tran (\sa_ctrl_rst_dat[9][11] , \sa_ctrl_rst_dat[9].r.part0[11] );
tran (\sa_ctrl_rst_dat[9][11] , \sa_ctrl_rst_dat[9].f.spare[6] );
tran (\sa_ctrl_rst_dat[9][12] , \sa_ctrl_rst_dat[9].r.part0[12] );
tran (\sa_ctrl_rst_dat[9][12] , \sa_ctrl_rst_dat[9].f.spare[7] );
tran (\sa_ctrl_rst_dat[9][13] , \sa_ctrl_rst_dat[9].r.part0[13] );
tran (\sa_ctrl_rst_dat[9][13] , \sa_ctrl_rst_dat[9].f.spare[8] );
tran (\sa_ctrl_rst_dat[9][14] , \sa_ctrl_rst_dat[9].r.part0[14] );
tran (\sa_ctrl_rst_dat[9][14] , \sa_ctrl_rst_dat[9].f.spare[9] );
tran (\sa_ctrl_rst_dat[9][15] , \sa_ctrl_rst_dat[9].r.part0[15] );
tran (\sa_ctrl_rst_dat[9][15] , \sa_ctrl_rst_dat[9].f.spare[10] );
tran (\sa_ctrl_rst_dat[9][16] , \sa_ctrl_rst_dat[9].r.part0[16] );
tran (\sa_ctrl_rst_dat[9][16] , \sa_ctrl_rst_dat[9].f.spare[11] );
tran (\sa_ctrl_rst_dat[9][17] , \sa_ctrl_rst_dat[9].r.part0[17] );
tran (\sa_ctrl_rst_dat[9][17] , \sa_ctrl_rst_dat[9].f.spare[12] );
tran (\sa_ctrl_rst_dat[9][18] , \sa_ctrl_rst_dat[9].r.part0[18] );
tran (\sa_ctrl_rst_dat[9][18] , \sa_ctrl_rst_dat[9].f.spare[13] );
tran (\sa_ctrl_rst_dat[9][19] , \sa_ctrl_rst_dat[9].r.part0[19] );
tran (\sa_ctrl_rst_dat[9][19] , \sa_ctrl_rst_dat[9].f.spare[14] );
tran (\sa_ctrl_rst_dat[9][20] , \sa_ctrl_rst_dat[9].r.part0[20] );
tran (\sa_ctrl_rst_dat[9][20] , \sa_ctrl_rst_dat[9].f.spare[15] );
tran (\sa_ctrl_rst_dat[9][21] , \sa_ctrl_rst_dat[9].r.part0[21] );
tran (\sa_ctrl_rst_dat[9][21] , \sa_ctrl_rst_dat[9].f.spare[16] );
tran (\sa_ctrl_rst_dat[9][22] , \sa_ctrl_rst_dat[9].r.part0[22] );
tran (\sa_ctrl_rst_dat[9][22] , \sa_ctrl_rst_dat[9].f.spare[17] );
tran (\sa_ctrl_rst_dat[9][23] , \sa_ctrl_rst_dat[9].r.part0[23] );
tran (\sa_ctrl_rst_dat[9][23] , \sa_ctrl_rst_dat[9].f.spare[18] );
tran (\sa_ctrl_rst_dat[9][24] , \sa_ctrl_rst_dat[9].r.part0[24] );
tran (\sa_ctrl_rst_dat[9][24] , \sa_ctrl_rst_dat[9].f.spare[19] );
tran (\sa_ctrl_rst_dat[9][25] , \sa_ctrl_rst_dat[9].r.part0[25] );
tran (\sa_ctrl_rst_dat[9][25] , \sa_ctrl_rst_dat[9].f.spare[20] );
tran (\sa_ctrl_rst_dat[9][26] , \sa_ctrl_rst_dat[9].r.part0[26] );
tran (\sa_ctrl_rst_dat[9][26] , \sa_ctrl_rst_dat[9].f.spare[21] );
tran (\sa_ctrl_rst_dat[9][27] , \sa_ctrl_rst_dat[9].r.part0[27] );
tran (\sa_ctrl_rst_dat[9][27] , \sa_ctrl_rst_dat[9].f.spare[22] );
tran (\sa_ctrl_rst_dat[9][28] , \sa_ctrl_rst_dat[9].r.part0[28] );
tran (\sa_ctrl_rst_dat[9][28] , \sa_ctrl_rst_dat[9].f.spare[23] );
tran (\sa_ctrl_rst_dat[9][29] , \sa_ctrl_rst_dat[9].r.part0[29] );
tran (\sa_ctrl_rst_dat[9][29] , \sa_ctrl_rst_dat[9].f.spare[24] );
tran (\sa_ctrl_rst_dat[9][30] , \sa_ctrl_rst_dat[9].r.part0[30] );
tran (\sa_ctrl_rst_dat[9][30] , \sa_ctrl_rst_dat[9].f.spare[25] );
tran (\sa_ctrl_rst_dat[9][31] , \sa_ctrl_rst_dat[9].r.part0[31] );
tran (\sa_ctrl_rst_dat[9][31] , \sa_ctrl_rst_dat[9].f.spare[26] );
tran (\sa_ctrl_rst_dat[10][0] , \sa_ctrl_rst_dat[10].r.part0[0] );
tran (\sa_ctrl_rst_dat[10][0] , \sa_ctrl_rst_dat[10].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[10][1] , \sa_ctrl_rst_dat[10].r.part0[1] );
tran (\sa_ctrl_rst_dat[10][1] , \sa_ctrl_rst_dat[10].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[10][2] , \sa_ctrl_rst_dat[10].r.part0[2] );
tran (\sa_ctrl_rst_dat[10][2] , \sa_ctrl_rst_dat[10].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[10][3] , \sa_ctrl_rst_dat[10].r.part0[3] );
tran (\sa_ctrl_rst_dat[10][3] , \sa_ctrl_rst_dat[10].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[10][4] , \sa_ctrl_rst_dat[10].r.part0[4] );
tran (\sa_ctrl_rst_dat[10][4] , \sa_ctrl_rst_dat[10].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[10][5] , \sa_ctrl_rst_dat[10].r.part0[5] );
tran (\sa_ctrl_rst_dat[10][5] , \sa_ctrl_rst_dat[10].f.spare[0] );
tran (\sa_ctrl_rst_dat[10][6] , \sa_ctrl_rst_dat[10].r.part0[6] );
tran (\sa_ctrl_rst_dat[10][6] , \sa_ctrl_rst_dat[10].f.spare[1] );
tran (\sa_ctrl_rst_dat[10][7] , \sa_ctrl_rst_dat[10].r.part0[7] );
tran (\sa_ctrl_rst_dat[10][7] , \sa_ctrl_rst_dat[10].f.spare[2] );
tran (\sa_ctrl_rst_dat[10][8] , \sa_ctrl_rst_dat[10].r.part0[8] );
tran (\sa_ctrl_rst_dat[10][8] , \sa_ctrl_rst_dat[10].f.spare[3] );
tran (\sa_ctrl_rst_dat[10][9] , \sa_ctrl_rst_dat[10].r.part0[9] );
tran (\sa_ctrl_rst_dat[10][9] , \sa_ctrl_rst_dat[10].f.spare[4] );
tran (\sa_ctrl_rst_dat[10][10] , \sa_ctrl_rst_dat[10].r.part0[10] );
tran (\sa_ctrl_rst_dat[10][10] , \sa_ctrl_rst_dat[10].f.spare[5] );
tran (\sa_ctrl_rst_dat[10][11] , \sa_ctrl_rst_dat[10].r.part0[11] );
tran (\sa_ctrl_rst_dat[10][11] , \sa_ctrl_rst_dat[10].f.spare[6] );
tran (\sa_ctrl_rst_dat[10][12] , \sa_ctrl_rst_dat[10].r.part0[12] );
tran (\sa_ctrl_rst_dat[10][12] , \sa_ctrl_rst_dat[10].f.spare[7] );
tran (\sa_ctrl_rst_dat[10][13] , \sa_ctrl_rst_dat[10].r.part0[13] );
tran (\sa_ctrl_rst_dat[10][13] , \sa_ctrl_rst_dat[10].f.spare[8] );
tran (\sa_ctrl_rst_dat[10][14] , \sa_ctrl_rst_dat[10].r.part0[14] );
tran (\sa_ctrl_rst_dat[10][14] , \sa_ctrl_rst_dat[10].f.spare[9] );
tran (\sa_ctrl_rst_dat[10][15] , \sa_ctrl_rst_dat[10].r.part0[15] );
tran (\sa_ctrl_rst_dat[10][15] , \sa_ctrl_rst_dat[10].f.spare[10] );
tran (\sa_ctrl_rst_dat[10][16] , \sa_ctrl_rst_dat[10].r.part0[16] );
tran (\sa_ctrl_rst_dat[10][16] , \sa_ctrl_rst_dat[10].f.spare[11] );
tran (\sa_ctrl_rst_dat[10][17] , \sa_ctrl_rst_dat[10].r.part0[17] );
tran (\sa_ctrl_rst_dat[10][17] , \sa_ctrl_rst_dat[10].f.spare[12] );
tran (\sa_ctrl_rst_dat[10][18] , \sa_ctrl_rst_dat[10].r.part0[18] );
tran (\sa_ctrl_rst_dat[10][18] , \sa_ctrl_rst_dat[10].f.spare[13] );
tran (\sa_ctrl_rst_dat[10][19] , \sa_ctrl_rst_dat[10].r.part0[19] );
tran (\sa_ctrl_rst_dat[10][19] , \sa_ctrl_rst_dat[10].f.spare[14] );
tran (\sa_ctrl_rst_dat[10][20] , \sa_ctrl_rst_dat[10].r.part0[20] );
tran (\sa_ctrl_rst_dat[10][20] , \sa_ctrl_rst_dat[10].f.spare[15] );
tran (\sa_ctrl_rst_dat[10][21] , \sa_ctrl_rst_dat[10].r.part0[21] );
tran (\sa_ctrl_rst_dat[10][21] , \sa_ctrl_rst_dat[10].f.spare[16] );
tran (\sa_ctrl_rst_dat[10][22] , \sa_ctrl_rst_dat[10].r.part0[22] );
tran (\sa_ctrl_rst_dat[10][22] , \sa_ctrl_rst_dat[10].f.spare[17] );
tran (\sa_ctrl_rst_dat[10][23] , \sa_ctrl_rst_dat[10].r.part0[23] );
tran (\sa_ctrl_rst_dat[10][23] , \sa_ctrl_rst_dat[10].f.spare[18] );
tran (\sa_ctrl_rst_dat[10][24] , \sa_ctrl_rst_dat[10].r.part0[24] );
tran (\sa_ctrl_rst_dat[10][24] , \sa_ctrl_rst_dat[10].f.spare[19] );
tran (\sa_ctrl_rst_dat[10][25] , \sa_ctrl_rst_dat[10].r.part0[25] );
tran (\sa_ctrl_rst_dat[10][25] , \sa_ctrl_rst_dat[10].f.spare[20] );
tran (\sa_ctrl_rst_dat[10][26] , \sa_ctrl_rst_dat[10].r.part0[26] );
tran (\sa_ctrl_rst_dat[10][26] , \sa_ctrl_rst_dat[10].f.spare[21] );
tran (\sa_ctrl_rst_dat[10][27] , \sa_ctrl_rst_dat[10].r.part0[27] );
tran (\sa_ctrl_rst_dat[10][27] , \sa_ctrl_rst_dat[10].f.spare[22] );
tran (\sa_ctrl_rst_dat[10][28] , \sa_ctrl_rst_dat[10].r.part0[28] );
tran (\sa_ctrl_rst_dat[10][28] , \sa_ctrl_rst_dat[10].f.spare[23] );
tran (\sa_ctrl_rst_dat[10][29] , \sa_ctrl_rst_dat[10].r.part0[29] );
tran (\sa_ctrl_rst_dat[10][29] , \sa_ctrl_rst_dat[10].f.spare[24] );
tran (\sa_ctrl_rst_dat[10][30] , \sa_ctrl_rst_dat[10].r.part0[30] );
tran (\sa_ctrl_rst_dat[10][30] , \sa_ctrl_rst_dat[10].f.spare[25] );
tran (\sa_ctrl_rst_dat[10][31] , \sa_ctrl_rst_dat[10].r.part0[31] );
tran (\sa_ctrl_rst_dat[10][31] , \sa_ctrl_rst_dat[10].f.spare[26] );
tran (\sa_ctrl_rst_dat[11][0] , \sa_ctrl_rst_dat[11].r.part0[0] );
tran (\sa_ctrl_rst_dat[11][0] , \sa_ctrl_rst_dat[11].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[11][1] , \sa_ctrl_rst_dat[11].r.part0[1] );
tran (\sa_ctrl_rst_dat[11][1] , \sa_ctrl_rst_dat[11].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[11][2] , \sa_ctrl_rst_dat[11].r.part0[2] );
tran (\sa_ctrl_rst_dat[11][2] , \sa_ctrl_rst_dat[11].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[11][3] , \sa_ctrl_rst_dat[11].r.part0[3] );
tran (\sa_ctrl_rst_dat[11][3] , \sa_ctrl_rst_dat[11].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[11][4] , \sa_ctrl_rst_dat[11].r.part0[4] );
tran (\sa_ctrl_rst_dat[11][4] , \sa_ctrl_rst_dat[11].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[11][5] , \sa_ctrl_rst_dat[11].r.part0[5] );
tran (\sa_ctrl_rst_dat[11][5] , \sa_ctrl_rst_dat[11].f.spare[0] );
tran (\sa_ctrl_rst_dat[11][6] , \sa_ctrl_rst_dat[11].r.part0[6] );
tran (\sa_ctrl_rst_dat[11][6] , \sa_ctrl_rst_dat[11].f.spare[1] );
tran (\sa_ctrl_rst_dat[11][7] , \sa_ctrl_rst_dat[11].r.part0[7] );
tran (\sa_ctrl_rst_dat[11][7] , \sa_ctrl_rst_dat[11].f.spare[2] );
tran (\sa_ctrl_rst_dat[11][8] , \sa_ctrl_rst_dat[11].r.part0[8] );
tran (\sa_ctrl_rst_dat[11][8] , \sa_ctrl_rst_dat[11].f.spare[3] );
tran (\sa_ctrl_rst_dat[11][9] , \sa_ctrl_rst_dat[11].r.part0[9] );
tran (\sa_ctrl_rst_dat[11][9] , \sa_ctrl_rst_dat[11].f.spare[4] );
tran (\sa_ctrl_rst_dat[11][10] , \sa_ctrl_rst_dat[11].r.part0[10] );
tran (\sa_ctrl_rst_dat[11][10] , \sa_ctrl_rst_dat[11].f.spare[5] );
tran (\sa_ctrl_rst_dat[11][11] , \sa_ctrl_rst_dat[11].r.part0[11] );
tran (\sa_ctrl_rst_dat[11][11] , \sa_ctrl_rst_dat[11].f.spare[6] );
tran (\sa_ctrl_rst_dat[11][12] , \sa_ctrl_rst_dat[11].r.part0[12] );
tran (\sa_ctrl_rst_dat[11][12] , \sa_ctrl_rst_dat[11].f.spare[7] );
tran (\sa_ctrl_rst_dat[11][13] , \sa_ctrl_rst_dat[11].r.part0[13] );
tran (\sa_ctrl_rst_dat[11][13] , \sa_ctrl_rst_dat[11].f.spare[8] );
tran (\sa_ctrl_rst_dat[11][14] , \sa_ctrl_rst_dat[11].r.part0[14] );
tran (\sa_ctrl_rst_dat[11][14] , \sa_ctrl_rst_dat[11].f.spare[9] );
tran (\sa_ctrl_rst_dat[11][15] , \sa_ctrl_rst_dat[11].r.part0[15] );
tran (\sa_ctrl_rst_dat[11][15] , \sa_ctrl_rst_dat[11].f.spare[10] );
tran (\sa_ctrl_rst_dat[11][16] , \sa_ctrl_rst_dat[11].r.part0[16] );
tran (\sa_ctrl_rst_dat[11][16] , \sa_ctrl_rst_dat[11].f.spare[11] );
tran (\sa_ctrl_rst_dat[11][17] , \sa_ctrl_rst_dat[11].r.part0[17] );
tran (\sa_ctrl_rst_dat[11][17] , \sa_ctrl_rst_dat[11].f.spare[12] );
tran (\sa_ctrl_rst_dat[11][18] , \sa_ctrl_rst_dat[11].r.part0[18] );
tran (\sa_ctrl_rst_dat[11][18] , \sa_ctrl_rst_dat[11].f.spare[13] );
tran (\sa_ctrl_rst_dat[11][19] , \sa_ctrl_rst_dat[11].r.part0[19] );
tran (\sa_ctrl_rst_dat[11][19] , \sa_ctrl_rst_dat[11].f.spare[14] );
tran (\sa_ctrl_rst_dat[11][20] , \sa_ctrl_rst_dat[11].r.part0[20] );
tran (\sa_ctrl_rst_dat[11][20] , \sa_ctrl_rst_dat[11].f.spare[15] );
tran (\sa_ctrl_rst_dat[11][21] , \sa_ctrl_rst_dat[11].r.part0[21] );
tran (\sa_ctrl_rst_dat[11][21] , \sa_ctrl_rst_dat[11].f.spare[16] );
tran (\sa_ctrl_rst_dat[11][22] , \sa_ctrl_rst_dat[11].r.part0[22] );
tran (\sa_ctrl_rst_dat[11][22] , \sa_ctrl_rst_dat[11].f.spare[17] );
tran (\sa_ctrl_rst_dat[11][23] , \sa_ctrl_rst_dat[11].r.part0[23] );
tran (\sa_ctrl_rst_dat[11][23] , \sa_ctrl_rst_dat[11].f.spare[18] );
tran (\sa_ctrl_rst_dat[11][24] , \sa_ctrl_rst_dat[11].r.part0[24] );
tran (\sa_ctrl_rst_dat[11][24] , \sa_ctrl_rst_dat[11].f.spare[19] );
tran (\sa_ctrl_rst_dat[11][25] , \sa_ctrl_rst_dat[11].r.part0[25] );
tran (\sa_ctrl_rst_dat[11][25] , \sa_ctrl_rst_dat[11].f.spare[20] );
tran (\sa_ctrl_rst_dat[11][26] , \sa_ctrl_rst_dat[11].r.part0[26] );
tran (\sa_ctrl_rst_dat[11][26] , \sa_ctrl_rst_dat[11].f.spare[21] );
tran (\sa_ctrl_rst_dat[11][27] , \sa_ctrl_rst_dat[11].r.part0[27] );
tran (\sa_ctrl_rst_dat[11][27] , \sa_ctrl_rst_dat[11].f.spare[22] );
tran (\sa_ctrl_rst_dat[11][28] , \sa_ctrl_rst_dat[11].r.part0[28] );
tran (\sa_ctrl_rst_dat[11][28] , \sa_ctrl_rst_dat[11].f.spare[23] );
tran (\sa_ctrl_rst_dat[11][29] , \sa_ctrl_rst_dat[11].r.part0[29] );
tran (\sa_ctrl_rst_dat[11][29] , \sa_ctrl_rst_dat[11].f.spare[24] );
tran (\sa_ctrl_rst_dat[11][30] , \sa_ctrl_rst_dat[11].r.part0[30] );
tran (\sa_ctrl_rst_dat[11][30] , \sa_ctrl_rst_dat[11].f.spare[25] );
tran (\sa_ctrl_rst_dat[11][31] , \sa_ctrl_rst_dat[11].r.part0[31] );
tran (\sa_ctrl_rst_dat[11][31] , \sa_ctrl_rst_dat[11].f.spare[26] );
tran (\sa_ctrl_rst_dat[12][0] , \sa_ctrl_rst_dat[12].r.part0[0] );
tran (\sa_ctrl_rst_dat[12][0] , \sa_ctrl_rst_dat[12].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[12][1] , \sa_ctrl_rst_dat[12].r.part0[1] );
tran (\sa_ctrl_rst_dat[12][1] , \sa_ctrl_rst_dat[12].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[12][2] , \sa_ctrl_rst_dat[12].r.part0[2] );
tran (\sa_ctrl_rst_dat[12][2] , \sa_ctrl_rst_dat[12].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[12][3] , \sa_ctrl_rst_dat[12].r.part0[3] );
tran (\sa_ctrl_rst_dat[12][3] , \sa_ctrl_rst_dat[12].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[12][4] , \sa_ctrl_rst_dat[12].r.part0[4] );
tran (\sa_ctrl_rst_dat[12][4] , \sa_ctrl_rst_dat[12].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[12][5] , \sa_ctrl_rst_dat[12].r.part0[5] );
tran (\sa_ctrl_rst_dat[12][5] , \sa_ctrl_rst_dat[12].f.spare[0] );
tran (\sa_ctrl_rst_dat[12][6] , \sa_ctrl_rst_dat[12].r.part0[6] );
tran (\sa_ctrl_rst_dat[12][6] , \sa_ctrl_rst_dat[12].f.spare[1] );
tran (\sa_ctrl_rst_dat[12][7] , \sa_ctrl_rst_dat[12].r.part0[7] );
tran (\sa_ctrl_rst_dat[12][7] , \sa_ctrl_rst_dat[12].f.spare[2] );
tran (\sa_ctrl_rst_dat[12][8] , \sa_ctrl_rst_dat[12].r.part0[8] );
tran (\sa_ctrl_rst_dat[12][8] , \sa_ctrl_rst_dat[12].f.spare[3] );
tran (\sa_ctrl_rst_dat[12][9] , \sa_ctrl_rst_dat[12].r.part0[9] );
tran (\sa_ctrl_rst_dat[12][9] , \sa_ctrl_rst_dat[12].f.spare[4] );
tran (\sa_ctrl_rst_dat[12][10] , \sa_ctrl_rst_dat[12].r.part0[10] );
tran (\sa_ctrl_rst_dat[12][10] , \sa_ctrl_rst_dat[12].f.spare[5] );
tran (\sa_ctrl_rst_dat[12][11] , \sa_ctrl_rst_dat[12].r.part0[11] );
tran (\sa_ctrl_rst_dat[12][11] , \sa_ctrl_rst_dat[12].f.spare[6] );
tran (\sa_ctrl_rst_dat[12][12] , \sa_ctrl_rst_dat[12].r.part0[12] );
tran (\sa_ctrl_rst_dat[12][12] , \sa_ctrl_rst_dat[12].f.spare[7] );
tran (\sa_ctrl_rst_dat[12][13] , \sa_ctrl_rst_dat[12].r.part0[13] );
tran (\sa_ctrl_rst_dat[12][13] , \sa_ctrl_rst_dat[12].f.spare[8] );
tran (\sa_ctrl_rst_dat[12][14] , \sa_ctrl_rst_dat[12].r.part0[14] );
tran (\sa_ctrl_rst_dat[12][14] , \sa_ctrl_rst_dat[12].f.spare[9] );
tran (\sa_ctrl_rst_dat[12][15] , \sa_ctrl_rst_dat[12].r.part0[15] );
tran (\sa_ctrl_rst_dat[12][15] , \sa_ctrl_rst_dat[12].f.spare[10] );
tran (\sa_ctrl_rst_dat[12][16] , \sa_ctrl_rst_dat[12].r.part0[16] );
tran (\sa_ctrl_rst_dat[12][16] , \sa_ctrl_rst_dat[12].f.spare[11] );
tran (\sa_ctrl_rst_dat[12][17] , \sa_ctrl_rst_dat[12].r.part0[17] );
tran (\sa_ctrl_rst_dat[12][17] , \sa_ctrl_rst_dat[12].f.spare[12] );
tran (\sa_ctrl_rst_dat[12][18] , \sa_ctrl_rst_dat[12].r.part0[18] );
tran (\sa_ctrl_rst_dat[12][18] , \sa_ctrl_rst_dat[12].f.spare[13] );
tran (\sa_ctrl_rst_dat[12][19] , \sa_ctrl_rst_dat[12].r.part0[19] );
tran (\sa_ctrl_rst_dat[12][19] , \sa_ctrl_rst_dat[12].f.spare[14] );
tran (\sa_ctrl_rst_dat[12][20] , \sa_ctrl_rst_dat[12].r.part0[20] );
tran (\sa_ctrl_rst_dat[12][20] , \sa_ctrl_rst_dat[12].f.spare[15] );
tran (\sa_ctrl_rst_dat[12][21] , \sa_ctrl_rst_dat[12].r.part0[21] );
tran (\sa_ctrl_rst_dat[12][21] , \sa_ctrl_rst_dat[12].f.spare[16] );
tran (\sa_ctrl_rst_dat[12][22] , \sa_ctrl_rst_dat[12].r.part0[22] );
tran (\sa_ctrl_rst_dat[12][22] , \sa_ctrl_rst_dat[12].f.spare[17] );
tran (\sa_ctrl_rst_dat[12][23] , \sa_ctrl_rst_dat[12].r.part0[23] );
tran (\sa_ctrl_rst_dat[12][23] , \sa_ctrl_rst_dat[12].f.spare[18] );
tran (\sa_ctrl_rst_dat[12][24] , \sa_ctrl_rst_dat[12].r.part0[24] );
tran (\sa_ctrl_rst_dat[12][24] , \sa_ctrl_rst_dat[12].f.spare[19] );
tran (\sa_ctrl_rst_dat[12][25] , \sa_ctrl_rst_dat[12].r.part0[25] );
tran (\sa_ctrl_rst_dat[12][25] , \sa_ctrl_rst_dat[12].f.spare[20] );
tran (\sa_ctrl_rst_dat[12][26] , \sa_ctrl_rst_dat[12].r.part0[26] );
tran (\sa_ctrl_rst_dat[12][26] , \sa_ctrl_rst_dat[12].f.spare[21] );
tran (\sa_ctrl_rst_dat[12][27] , \sa_ctrl_rst_dat[12].r.part0[27] );
tran (\sa_ctrl_rst_dat[12][27] , \sa_ctrl_rst_dat[12].f.spare[22] );
tran (\sa_ctrl_rst_dat[12][28] , \sa_ctrl_rst_dat[12].r.part0[28] );
tran (\sa_ctrl_rst_dat[12][28] , \sa_ctrl_rst_dat[12].f.spare[23] );
tran (\sa_ctrl_rst_dat[12][29] , \sa_ctrl_rst_dat[12].r.part0[29] );
tran (\sa_ctrl_rst_dat[12][29] , \sa_ctrl_rst_dat[12].f.spare[24] );
tran (\sa_ctrl_rst_dat[12][30] , \sa_ctrl_rst_dat[12].r.part0[30] );
tran (\sa_ctrl_rst_dat[12][30] , \sa_ctrl_rst_dat[12].f.spare[25] );
tran (\sa_ctrl_rst_dat[12][31] , \sa_ctrl_rst_dat[12].r.part0[31] );
tran (\sa_ctrl_rst_dat[12][31] , \sa_ctrl_rst_dat[12].f.spare[26] );
tran (\sa_ctrl_rst_dat[13][0] , \sa_ctrl_rst_dat[13].r.part0[0] );
tran (\sa_ctrl_rst_dat[13][0] , \sa_ctrl_rst_dat[13].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[13][1] , \sa_ctrl_rst_dat[13].r.part0[1] );
tran (\sa_ctrl_rst_dat[13][1] , \sa_ctrl_rst_dat[13].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[13][2] , \sa_ctrl_rst_dat[13].r.part0[2] );
tran (\sa_ctrl_rst_dat[13][2] , \sa_ctrl_rst_dat[13].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[13][3] , \sa_ctrl_rst_dat[13].r.part0[3] );
tran (\sa_ctrl_rst_dat[13][3] , \sa_ctrl_rst_dat[13].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[13][4] , \sa_ctrl_rst_dat[13].r.part0[4] );
tran (\sa_ctrl_rst_dat[13][4] , \sa_ctrl_rst_dat[13].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[13][5] , \sa_ctrl_rst_dat[13].r.part0[5] );
tran (\sa_ctrl_rst_dat[13][5] , \sa_ctrl_rst_dat[13].f.spare[0] );
tran (\sa_ctrl_rst_dat[13][6] , \sa_ctrl_rst_dat[13].r.part0[6] );
tran (\sa_ctrl_rst_dat[13][6] , \sa_ctrl_rst_dat[13].f.spare[1] );
tran (\sa_ctrl_rst_dat[13][7] , \sa_ctrl_rst_dat[13].r.part0[7] );
tran (\sa_ctrl_rst_dat[13][7] , \sa_ctrl_rst_dat[13].f.spare[2] );
tran (\sa_ctrl_rst_dat[13][8] , \sa_ctrl_rst_dat[13].r.part0[8] );
tran (\sa_ctrl_rst_dat[13][8] , \sa_ctrl_rst_dat[13].f.spare[3] );
tran (\sa_ctrl_rst_dat[13][9] , \sa_ctrl_rst_dat[13].r.part0[9] );
tran (\sa_ctrl_rst_dat[13][9] , \sa_ctrl_rst_dat[13].f.spare[4] );
tran (\sa_ctrl_rst_dat[13][10] , \sa_ctrl_rst_dat[13].r.part0[10] );
tran (\sa_ctrl_rst_dat[13][10] , \sa_ctrl_rst_dat[13].f.spare[5] );
tran (\sa_ctrl_rst_dat[13][11] , \sa_ctrl_rst_dat[13].r.part0[11] );
tran (\sa_ctrl_rst_dat[13][11] , \sa_ctrl_rst_dat[13].f.spare[6] );
tran (\sa_ctrl_rst_dat[13][12] , \sa_ctrl_rst_dat[13].r.part0[12] );
tran (\sa_ctrl_rst_dat[13][12] , \sa_ctrl_rst_dat[13].f.spare[7] );
tran (\sa_ctrl_rst_dat[13][13] , \sa_ctrl_rst_dat[13].r.part0[13] );
tran (\sa_ctrl_rst_dat[13][13] , \sa_ctrl_rst_dat[13].f.spare[8] );
tran (\sa_ctrl_rst_dat[13][14] , \sa_ctrl_rst_dat[13].r.part0[14] );
tran (\sa_ctrl_rst_dat[13][14] , \sa_ctrl_rst_dat[13].f.spare[9] );
tran (\sa_ctrl_rst_dat[13][15] , \sa_ctrl_rst_dat[13].r.part0[15] );
tran (\sa_ctrl_rst_dat[13][15] , \sa_ctrl_rst_dat[13].f.spare[10] );
tran (\sa_ctrl_rst_dat[13][16] , \sa_ctrl_rst_dat[13].r.part0[16] );
tran (\sa_ctrl_rst_dat[13][16] , \sa_ctrl_rst_dat[13].f.spare[11] );
tran (\sa_ctrl_rst_dat[13][17] , \sa_ctrl_rst_dat[13].r.part0[17] );
tran (\sa_ctrl_rst_dat[13][17] , \sa_ctrl_rst_dat[13].f.spare[12] );
tran (\sa_ctrl_rst_dat[13][18] , \sa_ctrl_rst_dat[13].r.part0[18] );
tran (\sa_ctrl_rst_dat[13][18] , \sa_ctrl_rst_dat[13].f.spare[13] );
tran (\sa_ctrl_rst_dat[13][19] , \sa_ctrl_rst_dat[13].r.part0[19] );
tran (\sa_ctrl_rst_dat[13][19] , \sa_ctrl_rst_dat[13].f.spare[14] );
tran (\sa_ctrl_rst_dat[13][20] , \sa_ctrl_rst_dat[13].r.part0[20] );
tran (\sa_ctrl_rst_dat[13][20] , \sa_ctrl_rst_dat[13].f.spare[15] );
tran (\sa_ctrl_rst_dat[13][21] , \sa_ctrl_rst_dat[13].r.part0[21] );
tran (\sa_ctrl_rst_dat[13][21] , \sa_ctrl_rst_dat[13].f.spare[16] );
tran (\sa_ctrl_rst_dat[13][22] , \sa_ctrl_rst_dat[13].r.part0[22] );
tran (\sa_ctrl_rst_dat[13][22] , \sa_ctrl_rst_dat[13].f.spare[17] );
tran (\sa_ctrl_rst_dat[13][23] , \sa_ctrl_rst_dat[13].r.part0[23] );
tran (\sa_ctrl_rst_dat[13][23] , \sa_ctrl_rst_dat[13].f.spare[18] );
tran (\sa_ctrl_rst_dat[13][24] , \sa_ctrl_rst_dat[13].r.part0[24] );
tran (\sa_ctrl_rst_dat[13][24] , \sa_ctrl_rst_dat[13].f.spare[19] );
tran (\sa_ctrl_rst_dat[13][25] , \sa_ctrl_rst_dat[13].r.part0[25] );
tran (\sa_ctrl_rst_dat[13][25] , \sa_ctrl_rst_dat[13].f.spare[20] );
tran (\sa_ctrl_rst_dat[13][26] , \sa_ctrl_rst_dat[13].r.part0[26] );
tran (\sa_ctrl_rst_dat[13][26] , \sa_ctrl_rst_dat[13].f.spare[21] );
tran (\sa_ctrl_rst_dat[13][27] , \sa_ctrl_rst_dat[13].r.part0[27] );
tran (\sa_ctrl_rst_dat[13][27] , \sa_ctrl_rst_dat[13].f.spare[22] );
tran (\sa_ctrl_rst_dat[13][28] , \sa_ctrl_rst_dat[13].r.part0[28] );
tran (\sa_ctrl_rst_dat[13][28] , \sa_ctrl_rst_dat[13].f.spare[23] );
tran (\sa_ctrl_rst_dat[13][29] , \sa_ctrl_rst_dat[13].r.part0[29] );
tran (\sa_ctrl_rst_dat[13][29] , \sa_ctrl_rst_dat[13].f.spare[24] );
tran (\sa_ctrl_rst_dat[13][30] , \sa_ctrl_rst_dat[13].r.part0[30] );
tran (\sa_ctrl_rst_dat[13][30] , \sa_ctrl_rst_dat[13].f.spare[25] );
tran (\sa_ctrl_rst_dat[13][31] , \sa_ctrl_rst_dat[13].r.part0[31] );
tran (\sa_ctrl_rst_dat[13][31] , \sa_ctrl_rst_dat[13].f.spare[26] );
tran (\sa_ctrl_rst_dat[14][0] , \sa_ctrl_rst_dat[14].r.part0[0] );
tran (\sa_ctrl_rst_dat[14][0] , \sa_ctrl_rst_dat[14].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[14][1] , \sa_ctrl_rst_dat[14].r.part0[1] );
tran (\sa_ctrl_rst_dat[14][1] , \sa_ctrl_rst_dat[14].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[14][2] , \sa_ctrl_rst_dat[14].r.part0[2] );
tran (\sa_ctrl_rst_dat[14][2] , \sa_ctrl_rst_dat[14].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[14][3] , \sa_ctrl_rst_dat[14].r.part0[3] );
tran (\sa_ctrl_rst_dat[14][3] , \sa_ctrl_rst_dat[14].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[14][4] , \sa_ctrl_rst_dat[14].r.part0[4] );
tran (\sa_ctrl_rst_dat[14][4] , \sa_ctrl_rst_dat[14].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[14][5] , \sa_ctrl_rst_dat[14].r.part0[5] );
tran (\sa_ctrl_rst_dat[14][5] , \sa_ctrl_rst_dat[14].f.spare[0] );
tran (\sa_ctrl_rst_dat[14][6] , \sa_ctrl_rst_dat[14].r.part0[6] );
tran (\sa_ctrl_rst_dat[14][6] , \sa_ctrl_rst_dat[14].f.spare[1] );
tran (\sa_ctrl_rst_dat[14][7] , \sa_ctrl_rst_dat[14].r.part0[7] );
tran (\sa_ctrl_rst_dat[14][7] , \sa_ctrl_rst_dat[14].f.spare[2] );
tran (\sa_ctrl_rst_dat[14][8] , \sa_ctrl_rst_dat[14].r.part0[8] );
tran (\sa_ctrl_rst_dat[14][8] , \sa_ctrl_rst_dat[14].f.spare[3] );
tran (\sa_ctrl_rst_dat[14][9] , \sa_ctrl_rst_dat[14].r.part0[9] );
tran (\sa_ctrl_rst_dat[14][9] , \sa_ctrl_rst_dat[14].f.spare[4] );
tran (\sa_ctrl_rst_dat[14][10] , \sa_ctrl_rst_dat[14].r.part0[10] );
tran (\sa_ctrl_rst_dat[14][10] , \sa_ctrl_rst_dat[14].f.spare[5] );
tran (\sa_ctrl_rst_dat[14][11] , \sa_ctrl_rst_dat[14].r.part0[11] );
tran (\sa_ctrl_rst_dat[14][11] , \sa_ctrl_rst_dat[14].f.spare[6] );
tran (\sa_ctrl_rst_dat[14][12] , \sa_ctrl_rst_dat[14].r.part0[12] );
tran (\sa_ctrl_rst_dat[14][12] , \sa_ctrl_rst_dat[14].f.spare[7] );
tran (\sa_ctrl_rst_dat[14][13] , \sa_ctrl_rst_dat[14].r.part0[13] );
tran (\sa_ctrl_rst_dat[14][13] , \sa_ctrl_rst_dat[14].f.spare[8] );
tran (\sa_ctrl_rst_dat[14][14] , \sa_ctrl_rst_dat[14].r.part0[14] );
tran (\sa_ctrl_rst_dat[14][14] , \sa_ctrl_rst_dat[14].f.spare[9] );
tran (\sa_ctrl_rst_dat[14][15] , \sa_ctrl_rst_dat[14].r.part0[15] );
tran (\sa_ctrl_rst_dat[14][15] , \sa_ctrl_rst_dat[14].f.spare[10] );
tran (\sa_ctrl_rst_dat[14][16] , \sa_ctrl_rst_dat[14].r.part0[16] );
tran (\sa_ctrl_rst_dat[14][16] , \sa_ctrl_rst_dat[14].f.spare[11] );
tran (\sa_ctrl_rst_dat[14][17] , \sa_ctrl_rst_dat[14].r.part0[17] );
tran (\sa_ctrl_rst_dat[14][17] , \sa_ctrl_rst_dat[14].f.spare[12] );
tran (\sa_ctrl_rst_dat[14][18] , \sa_ctrl_rst_dat[14].r.part0[18] );
tran (\sa_ctrl_rst_dat[14][18] , \sa_ctrl_rst_dat[14].f.spare[13] );
tran (\sa_ctrl_rst_dat[14][19] , \sa_ctrl_rst_dat[14].r.part0[19] );
tran (\sa_ctrl_rst_dat[14][19] , \sa_ctrl_rst_dat[14].f.spare[14] );
tran (\sa_ctrl_rst_dat[14][20] , \sa_ctrl_rst_dat[14].r.part0[20] );
tran (\sa_ctrl_rst_dat[14][20] , \sa_ctrl_rst_dat[14].f.spare[15] );
tran (\sa_ctrl_rst_dat[14][21] , \sa_ctrl_rst_dat[14].r.part0[21] );
tran (\sa_ctrl_rst_dat[14][21] , \sa_ctrl_rst_dat[14].f.spare[16] );
tran (\sa_ctrl_rst_dat[14][22] , \sa_ctrl_rst_dat[14].r.part0[22] );
tran (\sa_ctrl_rst_dat[14][22] , \sa_ctrl_rst_dat[14].f.spare[17] );
tran (\sa_ctrl_rst_dat[14][23] , \sa_ctrl_rst_dat[14].r.part0[23] );
tran (\sa_ctrl_rst_dat[14][23] , \sa_ctrl_rst_dat[14].f.spare[18] );
tran (\sa_ctrl_rst_dat[14][24] , \sa_ctrl_rst_dat[14].r.part0[24] );
tran (\sa_ctrl_rst_dat[14][24] , \sa_ctrl_rst_dat[14].f.spare[19] );
tran (\sa_ctrl_rst_dat[14][25] , \sa_ctrl_rst_dat[14].r.part0[25] );
tran (\sa_ctrl_rst_dat[14][25] , \sa_ctrl_rst_dat[14].f.spare[20] );
tran (\sa_ctrl_rst_dat[14][26] , \sa_ctrl_rst_dat[14].r.part0[26] );
tran (\sa_ctrl_rst_dat[14][26] , \sa_ctrl_rst_dat[14].f.spare[21] );
tran (\sa_ctrl_rst_dat[14][27] , \sa_ctrl_rst_dat[14].r.part0[27] );
tran (\sa_ctrl_rst_dat[14][27] , \sa_ctrl_rst_dat[14].f.spare[22] );
tran (\sa_ctrl_rst_dat[14][28] , \sa_ctrl_rst_dat[14].r.part0[28] );
tran (\sa_ctrl_rst_dat[14][28] , \sa_ctrl_rst_dat[14].f.spare[23] );
tran (\sa_ctrl_rst_dat[14][29] , \sa_ctrl_rst_dat[14].r.part0[29] );
tran (\sa_ctrl_rst_dat[14][29] , \sa_ctrl_rst_dat[14].f.spare[24] );
tran (\sa_ctrl_rst_dat[14][30] , \sa_ctrl_rst_dat[14].r.part0[30] );
tran (\sa_ctrl_rst_dat[14][30] , \sa_ctrl_rst_dat[14].f.spare[25] );
tran (\sa_ctrl_rst_dat[14][31] , \sa_ctrl_rst_dat[14].r.part0[31] );
tran (\sa_ctrl_rst_dat[14][31] , \sa_ctrl_rst_dat[14].f.spare[26] );
tran (\sa_ctrl_rst_dat[15][0] , \sa_ctrl_rst_dat[15].r.part0[0] );
tran (\sa_ctrl_rst_dat[15][0] , \sa_ctrl_rst_dat[15].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[15][1] , \sa_ctrl_rst_dat[15].r.part0[1] );
tran (\sa_ctrl_rst_dat[15][1] , \sa_ctrl_rst_dat[15].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[15][2] , \sa_ctrl_rst_dat[15].r.part0[2] );
tran (\sa_ctrl_rst_dat[15][2] , \sa_ctrl_rst_dat[15].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[15][3] , \sa_ctrl_rst_dat[15].r.part0[3] );
tran (\sa_ctrl_rst_dat[15][3] , \sa_ctrl_rst_dat[15].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[15][4] , \sa_ctrl_rst_dat[15].r.part0[4] );
tran (\sa_ctrl_rst_dat[15][4] , \sa_ctrl_rst_dat[15].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[15][5] , \sa_ctrl_rst_dat[15].r.part0[5] );
tran (\sa_ctrl_rst_dat[15][5] , \sa_ctrl_rst_dat[15].f.spare[0] );
tran (\sa_ctrl_rst_dat[15][6] , \sa_ctrl_rst_dat[15].r.part0[6] );
tran (\sa_ctrl_rst_dat[15][6] , \sa_ctrl_rst_dat[15].f.spare[1] );
tran (\sa_ctrl_rst_dat[15][7] , \sa_ctrl_rst_dat[15].r.part0[7] );
tran (\sa_ctrl_rst_dat[15][7] , \sa_ctrl_rst_dat[15].f.spare[2] );
tran (\sa_ctrl_rst_dat[15][8] , \sa_ctrl_rst_dat[15].r.part0[8] );
tran (\sa_ctrl_rst_dat[15][8] , \sa_ctrl_rst_dat[15].f.spare[3] );
tran (\sa_ctrl_rst_dat[15][9] , \sa_ctrl_rst_dat[15].r.part0[9] );
tran (\sa_ctrl_rst_dat[15][9] , \sa_ctrl_rst_dat[15].f.spare[4] );
tran (\sa_ctrl_rst_dat[15][10] , \sa_ctrl_rst_dat[15].r.part0[10] );
tran (\sa_ctrl_rst_dat[15][10] , \sa_ctrl_rst_dat[15].f.spare[5] );
tran (\sa_ctrl_rst_dat[15][11] , \sa_ctrl_rst_dat[15].r.part0[11] );
tran (\sa_ctrl_rst_dat[15][11] , \sa_ctrl_rst_dat[15].f.spare[6] );
tran (\sa_ctrl_rst_dat[15][12] , \sa_ctrl_rst_dat[15].r.part0[12] );
tran (\sa_ctrl_rst_dat[15][12] , \sa_ctrl_rst_dat[15].f.spare[7] );
tran (\sa_ctrl_rst_dat[15][13] , \sa_ctrl_rst_dat[15].r.part0[13] );
tran (\sa_ctrl_rst_dat[15][13] , \sa_ctrl_rst_dat[15].f.spare[8] );
tran (\sa_ctrl_rst_dat[15][14] , \sa_ctrl_rst_dat[15].r.part0[14] );
tran (\sa_ctrl_rst_dat[15][14] , \sa_ctrl_rst_dat[15].f.spare[9] );
tran (\sa_ctrl_rst_dat[15][15] , \sa_ctrl_rst_dat[15].r.part0[15] );
tran (\sa_ctrl_rst_dat[15][15] , \sa_ctrl_rst_dat[15].f.spare[10] );
tran (\sa_ctrl_rst_dat[15][16] , \sa_ctrl_rst_dat[15].r.part0[16] );
tran (\sa_ctrl_rst_dat[15][16] , \sa_ctrl_rst_dat[15].f.spare[11] );
tran (\sa_ctrl_rst_dat[15][17] , \sa_ctrl_rst_dat[15].r.part0[17] );
tran (\sa_ctrl_rst_dat[15][17] , \sa_ctrl_rst_dat[15].f.spare[12] );
tran (\sa_ctrl_rst_dat[15][18] , \sa_ctrl_rst_dat[15].r.part0[18] );
tran (\sa_ctrl_rst_dat[15][18] , \sa_ctrl_rst_dat[15].f.spare[13] );
tran (\sa_ctrl_rst_dat[15][19] , \sa_ctrl_rst_dat[15].r.part0[19] );
tran (\sa_ctrl_rst_dat[15][19] , \sa_ctrl_rst_dat[15].f.spare[14] );
tran (\sa_ctrl_rst_dat[15][20] , \sa_ctrl_rst_dat[15].r.part0[20] );
tran (\sa_ctrl_rst_dat[15][20] , \sa_ctrl_rst_dat[15].f.spare[15] );
tran (\sa_ctrl_rst_dat[15][21] , \sa_ctrl_rst_dat[15].r.part0[21] );
tran (\sa_ctrl_rst_dat[15][21] , \sa_ctrl_rst_dat[15].f.spare[16] );
tran (\sa_ctrl_rst_dat[15][22] , \sa_ctrl_rst_dat[15].r.part0[22] );
tran (\sa_ctrl_rst_dat[15][22] , \sa_ctrl_rst_dat[15].f.spare[17] );
tran (\sa_ctrl_rst_dat[15][23] , \sa_ctrl_rst_dat[15].r.part0[23] );
tran (\sa_ctrl_rst_dat[15][23] , \sa_ctrl_rst_dat[15].f.spare[18] );
tran (\sa_ctrl_rst_dat[15][24] , \sa_ctrl_rst_dat[15].r.part0[24] );
tran (\sa_ctrl_rst_dat[15][24] , \sa_ctrl_rst_dat[15].f.spare[19] );
tran (\sa_ctrl_rst_dat[15][25] , \sa_ctrl_rst_dat[15].r.part0[25] );
tran (\sa_ctrl_rst_dat[15][25] , \sa_ctrl_rst_dat[15].f.spare[20] );
tran (\sa_ctrl_rst_dat[15][26] , \sa_ctrl_rst_dat[15].r.part0[26] );
tran (\sa_ctrl_rst_dat[15][26] , \sa_ctrl_rst_dat[15].f.spare[21] );
tran (\sa_ctrl_rst_dat[15][27] , \sa_ctrl_rst_dat[15].r.part0[27] );
tran (\sa_ctrl_rst_dat[15][27] , \sa_ctrl_rst_dat[15].f.spare[22] );
tran (\sa_ctrl_rst_dat[15][28] , \sa_ctrl_rst_dat[15].r.part0[28] );
tran (\sa_ctrl_rst_dat[15][28] , \sa_ctrl_rst_dat[15].f.spare[23] );
tran (\sa_ctrl_rst_dat[15][29] , \sa_ctrl_rst_dat[15].r.part0[29] );
tran (\sa_ctrl_rst_dat[15][29] , \sa_ctrl_rst_dat[15].f.spare[24] );
tran (\sa_ctrl_rst_dat[15][30] , \sa_ctrl_rst_dat[15].r.part0[30] );
tran (\sa_ctrl_rst_dat[15][30] , \sa_ctrl_rst_dat[15].f.spare[25] );
tran (\sa_ctrl_rst_dat[15][31] , \sa_ctrl_rst_dat[15].r.part0[31] );
tran (\sa_ctrl_rst_dat[15][31] , \sa_ctrl_rst_dat[15].f.spare[26] );
tran (\sa_ctrl_rst_dat[16][0] , \sa_ctrl_rst_dat[16].r.part0[0] );
tran (\sa_ctrl_rst_dat[16][0] , \sa_ctrl_rst_dat[16].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[16][1] , \sa_ctrl_rst_dat[16].r.part0[1] );
tran (\sa_ctrl_rst_dat[16][1] , \sa_ctrl_rst_dat[16].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[16][2] , \sa_ctrl_rst_dat[16].r.part0[2] );
tran (\sa_ctrl_rst_dat[16][2] , \sa_ctrl_rst_dat[16].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[16][3] , \sa_ctrl_rst_dat[16].r.part0[3] );
tran (\sa_ctrl_rst_dat[16][3] , \sa_ctrl_rst_dat[16].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[16][4] , \sa_ctrl_rst_dat[16].r.part0[4] );
tran (\sa_ctrl_rst_dat[16][4] , \sa_ctrl_rst_dat[16].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[16][5] , \sa_ctrl_rst_dat[16].r.part0[5] );
tran (\sa_ctrl_rst_dat[16][5] , \sa_ctrl_rst_dat[16].f.spare[0] );
tran (\sa_ctrl_rst_dat[16][6] , \sa_ctrl_rst_dat[16].r.part0[6] );
tran (\sa_ctrl_rst_dat[16][6] , \sa_ctrl_rst_dat[16].f.spare[1] );
tran (\sa_ctrl_rst_dat[16][7] , \sa_ctrl_rst_dat[16].r.part0[7] );
tran (\sa_ctrl_rst_dat[16][7] , \sa_ctrl_rst_dat[16].f.spare[2] );
tran (\sa_ctrl_rst_dat[16][8] , \sa_ctrl_rst_dat[16].r.part0[8] );
tran (\sa_ctrl_rst_dat[16][8] , \sa_ctrl_rst_dat[16].f.spare[3] );
tran (\sa_ctrl_rst_dat[16][9] , \sa_ctrl_rst_dat[16].r.part0[9] );
tran (\sa_ctrl_rst_dat[16][9] , \sa_ctrl_rst_dat[16].f.spare[4] );
tran (\sa_ctrl_rst_dat[16][10] , \sa_ctrl_rst_dat[16].r.part0[10] );
tran (\sa_ctrl_rst_dat[16][10] , \sa_ctrl_rst_dat[16].f.spare[5] );
tran (\sa_ctrl_rst_dat[16][11] , \sa_ctrl_rst_dat[16].r.part0[11] );
tran (\sa_ctrl_rst_dat[16][11] , \sa_ctrl_rst_dat[16].f.spare[6] );
tran (\sa_ctrl_rst_dat[16][12] , \sa_ctrl_rst_dat[16].r.part0[12] );
tran (\sa_ctrl_rst_dat[16][12] , \sa_ctrl_rst_dat[16].f.spare[7] );
tran (\sa_ctrl_rst_dat[16][13] , \sa_ctrl_rst_dat[16].r.part0[13] );
tran (\sa_ctrl_rst_dat[16][13] , \sa_ctrl_rst_dat[16].f.spare[8] );
tran (\sa_ctrl_rst_dat[16][14] , \sa_ctrl_rst_dat[16].r.part0[14] );
tran (\sa_ctrl_rst_dat[16][14] , \sa_ctrl_rst_dat[16].f.spare[9] );
tran (\sa_ctrl_rst_dat[16][15] , \sa_ctrl_rst_dat[16].r.part0[15] );
tran (\sa_ctrl_rst_dat[16][15] , \sa_ctrl_rst_dat[16].f.spare[10] );
tran (\sa_ctrl_rst_dat[16][16] , \sa_ctrl_rst_dat[16].r.part0[16] );
tran (\sa_ctrl_rst_dat[16][16] , \sa_ctrl_rst_dat[16].f.spare[11] );
tran (\sa_ctrl_rst_dat[16][17] , \sa_ctrl_rst_dat[16].r.part0[17] );
tran (\sa_ctrl_rst_dat[16][17] , \sa_ctrl_rst_dat[16].f.spare[12] );
tran (\sa_ctrl_rst_dat[16][18] , \sa_ctrl_rst_dat[16].r.part0[18] );
tran (\sa_ctrl_rst_dat[16][18] , \sa_ctrl_rst_dat[16].f.spare[13] );
tran (\sa_ctrl_rst_dat[16][19] , \sa_ctrl_rst_dat[16].r.part0[19] );
tran (\sa_ctrl_rst_dat[16][19] , \sa_ctrl_rst_dat[16].f.spare[14] );
tran (\sa_ctrl_rst_dat[16][20] , \sa_ctrl_rst_dat[16].r.part0[20] );
tran (\sa_ctrl_rst_dat[16][20] , \sa_ctrl_rst_dat[16].f.spare[15] );
tran (\sa_ctrl_rst_dat[16][21] , \sa_ctrl_rst_dat[16].r.part0[21] );
tran (\sa_ctrl_rst_dat[16][21] , \sa_ctrl_rst_dat[16].f.spare[16] );
tran (\sa_ctrl_rst_dat[16][22] , \sa_ctrl_rst_dat[16].r.part0[22] );
tran (\sa_ctrl_rst_dat[16][22] , \sa_ctrl_rst_dat[16].f.spare[17] );
tran (\sa_ctrl_rst_dat[16][23] , \sa_ctrl_rst_dat[16].r.part0[23] );
tran (\sa_ctrl_rst_dat[16][23] , \sa_ctrl_rst_dat[16].f.spare[18] );
tran (\sa_ctrl_rst_dat[16][24] , \sa_ctrl_rst_dat[16].r.part0[24] );
tran (\sa_ctrl_rst_dat[16][24] , \sa_ctrl_rst_dat[16].f.spare[19] );
tran (\sa_ctrl_rst_dat[16][25] , \sa_ctrl_rst_dat[16].r.part0[25] );
tran (\sa_ctrl_rst_dat[16][25] , \sa_ctrl_rst_dat[16].f.spare[20] );
tran (\sa_ctrl_rst_dat[16][26] , \sa_ctrl_rst_dat[16].r.part0[26] );
tran (\sa_ctrl_rst_dat[16][26] , \sa_ctrl_rst_dat[16].f.spare[21] );
tran (\sa_ctrl_rst_dat[16][27] , \sa_ctrl_rst_dat[16].r.part0[27] );
tran (\sa_ctrl_rst_dat[16][27] , \sa_ctrl_rst_dat[16].f.spare[22] );
tran (\sa_ctrl_rst_dat[16][28] , \sa_ctrl_rst_dat[16].r.part0[28] );
tran (\sa_ctrl_rst_dat[16][28] , \sa_ctrl_rst_dat[16].f.spare[23] );
tran (\sa_ctrl_rst_dat[16][29] , \sa_ctrl_rst_dat[16].r.part0[29] );
tran (\sa_ctrl_rst_dat[16][29] , \sa_ctrl_rst_dat[16].f.spare[24] );
tran (\sa_ctrl_rst_dat[16][30] , \sa_ctrl_rst_dat[16].r.part0[30] );
tran (\sa_ctrl_rst_dat[16][30] , \sa_ctrl_rst_dat[16].f.spare[25] );
tran (\sa_ctrl_rst_dat[16][31] , \sa_ctrl_rst_dat[16].r.part0[31] );
tran (\sa_ctrl_rst_dat[16][31] , \sa_ctrl_rst_dat[16].f.spare[26] );
tran (\sa_ctrl_rst_dat[17][0] , \sa_ctrl_rst_dat[17].r.part0[0] );
tran (\sa_ctrl_rst_dat[17][0] , \sa_ctrl_rst_dat[17].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[17][1] , \sa_ctrl_rst_dat[17].r.part0[1] );
tran (\sa_ctrl_rst_dat[17][1] , \sa_ctrl_rst_dat[17].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[17][2] , \sa_ctrl_rst_dat[17].r.part0[2] );
tran (\sa_ctrl_rst_dat[17][2] , \sa_ctrl_rst_dat[17].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[17][3] , \sa_ctrl_rst_dat[17].r.part0[3] );
tran (\sa_ctrl_rst_dat[17][3] , \sa_ctrl_rst_dat[17].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[17][4] , \sa_ctrl_rst_dat[17].r.part0[4] );
tran (\sa_ctrl_rst_dat[17][4] , \sa_ctrl_rst_dat[17].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[17][5] , \sa_ctrl_rst_dat[17].r.part0[5] );
tran (\sa_ctrl_rst_dat[17][5] , \sa_ctrl_rst_dat[17].f.spare[0] );
tran (\sa_ctrl_rst_dat[17][6] , \sa_ctrl_rst_dat[17].r.part0[6] );
tran (\sa_ctrl_rst_dat[17][6] , \sa_ctrl_rst_dat[17].f.spare[1] );
tran (\sa_ctrl_rst_dat[17][7] , \sa_ctrl_rst_dat[17].r.part0[7] );
tran (\sa_ctrl_rst_dat[17][7] , \sa_ctrl_rst_dat[17].f.spare[2] );
tran (\sa_ctrl_rst_dat[17][8] , \sa_ctrl_rst_dat[17].r.part0[8] );
tran (\sa_ctrl_rst_dat[17][8] , \sa_ctrl_rst_dat[17].f.spare[3] );
tran (\sa_ctrl_rst_dat[17][9] , \sa_ctrl_rst_dat[17].r.part0[9] );
tran (\sa_ctrl_rst_dat[17][9] , \sa_ctrl_rst_dat[17].f.spare[4] );
tran (\sa_ctrl_rst_dat[17][10] , \sa_ctrl_rst_dat[17].r.part0[10] );
tran (\sa_ctrl_rst_dat[17][10] , \sa_ctrl_rst_dat[17].f.spare[5] );
tran (\sa_ctrl_rst_dat[17][11] , \sa_ctrl_rst_dat[17].r.part0[11] );
tran (\sa_ctrl_rst_dat[17][11] , \sa_ctrl_rst_dat[17].f.spare[6] );
tran (\sa_ctrl_rst_dat[17][12] , \sa_ctrl_rst_dat[17].r.part0[12] );
tran (\sa_ctrl_rst_dat[17][12] , \sa_ctrl_rst_dat[17].f.spare[7] );
tran (\sa_ctrl_rst_dat[17][13] , \sa_ctrl_rst_dat[17].r.part0[13] );
tran (\sa_ctrl_rst_dat[17][13] , \sa_ctrl_rst_dat[17].f.spare[8] );
tran (\sa_ctrl_rst_dat[17][14] , \sa_ctrl_rst_dat[17].r.part0[14] );
tran (\sa_ctrl_rst_dat[17][14] , \sa_ctrl_rst_dat[17].f.spare[9] );
tran (\sa_ctrl_rst_dat[17][15] , \sa_ctrl_rst_dat[17].r.part0[15] );
tran (\sa_ctrl_rst_dat[17][15] , \sa_ctrl_rst_dat[17].f.spare[10] );
tran (\sa_ctrl_rst_dat[17][16] , \sa_ctrl_rst_dat[17].r.part0[16] );
tran (\sa_ctrl_rst_dat[17][16] , \sa_ctrl_rst_dat[17].f.spare[11] );
tran (\sa_ctrl_rst_dat[17][17] , \sa_ctrl_rst_dat[17].r.part0[17] );
tran (\sa_ctrl_rst_dat[17][17] , \sa_ctrl_rst_dat[17].f.spare[12] );
tran (\sa_ctrl_rst_dat[17][18] , \sa_ctrl_rst_dat[17].r.part0[18] );
tran (\sa_ctrl_rst_dat[17][18] , \sa_ctrl_rst_dat[17].f.spare[13] );
tran (\sa_ctrl_rst_dat[17][19] , \sa_ctrl_rst_dat[17].r.part0[19] );
tran (\sa_ctrl_rst_dat[17][19] , \sa_ctrl_rst_dat[17].f.spare[14] );
tran (\sa_ctrl_rst_dat[17][20] , \sa_ctrl_rst_dat[17].r.part0[20] );
tran (\sa_ctrl_rst_dat[17][20] , \sa_ctrl_rst_dat[17].f.spare[15] );
tran (\sa_ctrl_rst_dat[17][21] , \sa_ctrl_rst_dat[17].r.part0[21] );
tran (\sa_ctrl_rst_dat[17][21] , \sa_ctrl_rst_dat[17].f.spare[16] );
tran (\sa_ctrl_rst_dat[17][22] , \sa_ctrl_rst_dat[17].r.part0[22] );
tran (\sa_ctrl_rst_dat[17][22] , \sa_ctrl_rst_dat[17].f.spare[17] );
tran (\sa_ctrl_rst_dat[17][23] , \sa_ctrl_rst_dat[17].r.part0[23] );
tran (\sa_ctrl_rst_dat[17][23] , \sa_ctrl_rst_dat[17].f.spare[18] );
tran (\sa_ctrl_rst_dat[17][24] , \sa_ctrl_rst_dat[17].r.part0[24] );
tran (\sa_ctrl_rst_dat[17][24] , \sa_ctrl_rst_dat[17].f.spare[19] );
tran (\sa_ctrl_rst_dat[17][25] , \sa_ctrl_rst_dat[17].r.part0[25] );
tran (\sa_ctrl_rst_dat[17][25] , \sa_ctrl_rst_dat[17].f.spare[20] );
tran (\sa_ctrl_rst_dat[17][26] , \sa_ctrl_rst_dat[17].r.part0[26] );
tran (\sa_ctrl_rst_dat[17][26] , \sa_ctrl_rst_dat[17].f.spare[21] );
tran (\sa_ctrl_rst_dat[17][27] , \sa_ctrl_rst_dat[17].r.part0[27] );
tran (\sa_ctrl_rst_dat[17][27] , \sa_ctrl_rst_dat[17].f.spare[22] );
tran (\sa_ctrl_rst_dat[17][28] , \sa_ctrl_rst_dat[17].r.part0[28] );
tran (\sa_ctrl_rst_dat[17][28] , \sa_ctrl_rst_dat[17].f.spare[23] );
tran (\sa_ctrl_rst_dat[17][29] , \sa_ctrl_rst_dat[17].r.part0[29] );
tran (\sa_ctrl_rst_dat[17][29] , \sa_ctrl_rst_dat[17].f.spare[24] );
tran (\sa_ctrl_rst_dat[17][30] , \sa_ctrl_rst_dat[17].r.part0[30] );
tran (\sa_ctrl_rst_dat[17][30] , \sa_ctrl_rst_dat[17].f.spare[25] );
tran (\sa_ctrl_rst_dat[17][31] , \sa_ctrl_rst_dat[17].r.part0[31] );
tran (\sa_ctrl_rst_dat[17][31] , \sa_ctrl_rst_dat[17].f.spare[26] );
tran (\sa_ctrl_rst_dat[18][0] , \sa_ctrl_rst_dat[18].r.part0[0] );
tran (\sa_ctrl_rst_dat[18][0] , \sa_ctrl_rst_dat[18].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[18][1] , \sa_ctrl_rst_dat[18].r.part0[1] );
tran (\sa_ctrl_rst_dat[18][1] , \sa_ctrl_rst_dat[18].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[18][2] , \sa_ctrl_rst_dat[18].r.part0[2] );
tran (\sa_ctrl_rst_dat[18][2] , \sa_ctrl_rst_dat[18].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[18][3] , \sa_ctrl_rst_dat[18].r.part0[3] );
tran (\sa_ctrl_rst_dat[18][3] , \sa_ctrl_rst_dat[18].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[18][4] , \sa_ctrl_rst_dat[18].r.part0[4] );
tran (\sa_ctrl_rst_dat[18][4] , \sa_ctrl_rst_dat[18].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[18][5] , \sa_ctrl_rst_dat[18].r.part0[5] );
tran (\sa_ctrl_rst_dat[18][5] , \sa_ctrl_rst_dat[18].f.spare[0] );
tran (\sa_ctrl_rst_dat[18][6] , \sa_ctrl_rst_dat[18].r.part0[6] );
tran (\sa_ctrl_rst_dat[18][6] , \sa_ctrl_rst_dat[18].f.spare[1] );
tran (\sa_ctrl_rst_dat[18][7] , \sa_ctrl_rst_dat[18].r.part0[7] );
tran (\sa_ctrl_rst_dat[18][7] , \sa_ctrl_rst_dat[18].f.spare[2] );
tran (\sa_ctrl_rst_dat[18][8] , \sa_ctrl_rst_dat[18].r.part0[8] );
tran (\sa_ctrl_rst_dat[18][8] , \sa_ctrl_rst_dat[18].f.spare[3] );
tran (\sa_ctrl_rst_dat[18][9] , \sa_ctrl_rst_dat[18].r.part0[9] );
tran (\sa_ctrl_rst_dat[18][9] , \sa_ctrl_rst_dat[18].f.spare[4] );
tran (\sa_ctrl_rst_dat[18][10] , \sa_ctrl_rst_dat[18].r.part0[10] );
tran (\sa_ctrl_rst_dat[18][10] , \sa_ctrl_rst_dat[18].f.spare[5] );
tran (\sa_ctrl_rst_dat[18][11] , \sa_ctrl_rst_dat[18].r.part0[11] );
tran (\sa_ctrl_rst_dat[18][11] , \sa_ctrl_rst_dat[18].f.spare[6] );
tran (\sa_ctrl_rst_dat[18][12] , \sa_ctrl_rst_dat[18].r.part0[12] );
tran (\sa_ctrl_rst_dat[18][12] , \sa_ctrl_rst_dat[18].f.spare[7] );
tran (\sa_ctrl_rst_dat[18][13] , \sa_ctrl_rst_dat[18].r.part0[13] );
tran (\sa_ctrl_rst_dat[18][13] , \sa_ctrl_rst_dat[18].f.spare[8] );
tran (\sa_ctrl_rst_dat[18][14] , \sa_ctrl_rst_dat[18].r.part0[14] );
tran (\sa_ctrl_rst_dat[18][14] , \sa_ctrl_rst_dat[18].f.spare[9] );
tran (\sa_ctrl_rst_dat[18][15] , \sa_ctrl_rst_dat[18].r.part0[15] );
tran (\sa_ctrl_rst_dat[18][15] , \sa_ctrl_rst_dat[18].f.spare[10] );
tran (\sa_ctrl_rst_dat[18][16] , \sa_ctrl_rst_dat[18].r.part0[16] );
tran (\sa_ctrl_rst_dat[18][16] , \sa_ctrl_rst_dat[18].f.spare[11] );
tran (\sa_ctrl_rst_dat[18][17] , \sa_ctrl_rst_dat[18].r.part0[17] );
tran (\sa_ctrl_rst_dat[18][17] , \sa_ctrl_rst_dat[18].f.spare[12] );
tran (\sa_ctrl_rst_dat[18][18] , \sa_ctrl_rst_dat[18].r.part0[18] );
tran (\sa_ctrl_rst_dat[18][18] , \sa_ctrl_rst_dat[18].f.spare[13] );
tran (\sa_ctrl_rst_dat[18][19] , \sa_ctrl_rst_dat[18].r.part0[19] );
tran (\sa_ctrl_rst_dat[18][19] , \sa_ctrl_rst_dat[18].f.spare[14] );
tran (\sa_ctrl_rst_dat[18][20] , \sa_ctrl_rst_dat[18].r.part0[20] );
tran (\sa_ctrl_rst_dat[18][20] , \sa_ctrl_rst_dat[18].f.spare[15] );
tran (\sa_ctrl_rst_dat[18][21] , \sa_ctrl_rst_dat[18].r.part0[21] );
tran (\sa_ctrl_rst_dat[18][21] , \sa_ctrl_rst_dat[18].f.spare[16] );
tran (\sa_ctrl_rst_dat[18][22] , \sa_ctrl_rst_dat[18].r.part0[22] );
tran (\sa_ctrl_rst_dat[18][22] , \sa_ctrl_rst_dat[18].f.spare[17] );
tran (\sa_ctrl_rst_dat[18][23] , \sa_ctrl_rst_dat[18].r.part0[23] );
tran (\sa_ctrl_rst_dat[18][23] , \sa_ctrl_rst_dat[18].f.spare[18] );
tran (\sa_ctrl_rst_dat[18][24] , \sa_ctrl_rst_dat[18].r.part0[24] );
tran (\sa_ctrl_rst_dat[18][24] , \sa_ctrl_rst_dat[18].f.spare[19] );
tran (\sa_ctrl_rst_dat[18][25] , \sa_ctrl_rst_dat[18].r.part0[25] );
tran (\sa_ctrl_rst_dat[18][25] , \sa_ctrl_rst_dat[18].f.spare[20] );
tran (\sa_ctrl_rst_dat[18][26] , \sa_ctrl_rst_dat[18].r.part0[26] );
tran (\sa_ctrl_rst_dat[18][26] , \sa_ctrl_rst_dat[18].f.spare[21] );
tran (\sa_ctrl_rst_dat[18][27] , \sa_ctrl_rst_dat[18].r.part0[27] );
tran (\sa_ctrl_rst_dat[18][27] , \sa_ctrl_rst_dat[18].f.spare[22] );
tran (\sa_ctrl_rst_dat[18][28] , \sa_ctrl_rst_dat[18].r.part0[28] );
tran (\sa_ctrl_rst_dat[18][28] , \sa_ctrl_rst_dat[18].f.spare[23] );
tran (\sa_ctrl_rst_dat[18][29] , \sa_ctrl_rst_dat[18].r.part0[29] );
tran (\sa_ctrl_rst_dat[18][29] , \sa_ctrl_rst_dat[18].f.spare[24] );
tran (\sa_ctrl_rst_dat[18][30] , \sa_ctrl_rst_dat[18].r.part0[30] );
tran (\sa_ctrl_rst_dat[18][30] , \sa_ctrl_rst_dat[18].f.spare[25] );
tran (\sa_ctrl_rst_dat[18][31] , \sa_ctrl_rst_dat[18].r.part0[31] );
tran (\sa_ctrl_rst_dat[18][31] , \sa_ctrl_rst_dat[18].f.spare[26] );
tran (\sa_ctrl_rst_dat[19][0] , \sa_ctrl_rst_dat[19].r.part0[0] );
tran (\sa_ctrl_rst_dat[19][0] , \sa_ctrl_rst_dat[19].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[19][1] , \sa_ctrl_rst_dat[19].r.part0[1] );
tran (\sa_ctrl_rst_dat[19][1] , \sa_ctrl_rst_dat[19].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[19][2] , \sa_ctrl_rst_dat[19].r.part0[2] );
tran (\sa_ctrl_rst_dat[19][2] , \sa_ctrl_rst_dat[19].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[19][3] , \sa_ctrl_rst_dat[19].r.part0[3] );
tran (\sa_ctrl_rst_dat[19][3] , \sa_ctrl_rst_dat[19].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[19][4] , \sa_ctrl_rst_dat[19].r.part0[4] );
tran (\sa_ctrl_rst_dat[19][4] , \sa_ctrl_rst_dat[19].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[19][5] , \sa_ctrl_rst_dat[19].r.part0[5] );
tran (\sa_ctrl_rst_dat[19][5] , \sa_ctrl_rst_dat[19].f.spare[0] );
tran (\sa_ctrl_rst_dat[19][6] , \sa_ctrl_rst_dat[19].r.part0[6] );
tran (\sa_ctrl_rst_dat[19][6] , \sa_ctrl_rst_dat[19].f.spare[1] );
tran (\sa_ctrl_rst_dat[19][7] , \sa_ctrl_rst_dat[19].r.part0[7] );
tran (\sa_ctrl_rst_dat[19][7] , \sa_ctrl_rst_dat[19].f.spare[2] );
tran (\sa_ctrl_rst_dat[19][8] , \sa_ctrl_rst_dat[19].r.part0[8] );
tran (\sa_ctrl_rst_dat[19][8] , \sa_ctrl_rst_dat[19].f.spare[3] );
tran (\sa_ctrl_rst_dat[19][9] , \sa_ctrl_rst_dat[19].r.part0[9] );
tran (\sa_ctrl_rst_dat[19][9] , \sa_ctrl_rst_dat[19].f.spare[4] );
tran (\sa_ctrl_rst_dat[19][10] , \sa_ctrl_rst_dat[19].r.part0[10] );
tran (\sa_ctrl_rst_dat[19][10] , \sa_ctrl_rst_dat[19].f.spare[5] );
tran (\sa_ctrl_rst_dat[19][11] , \sa_ctrl_rst_dat[19].r.part0[11] );
tran (\sa_ctrl_rst_dat[19][11] , \sa_ctrl_rst_dat[19].f.spare[6] );
tran (\sa_ctrl_rst_dat[19][12] , \sa_ctrl_rst_dat[19].r.part0[12] );
tran (\sa_ctrl_rst_dat[19][12] , \sa_ctrl_rst_dat[19].f.spare[7] );
tran (\sa_ctrl_rst_dat[19][13] , \sa_ctrl_rst_dat[19].r.part0[13] );
tran (\sa_ctrl_rst_dat[19][13] , \sa_ctrl_rst_dat[19].f.spare[8] );
tran (\sa_ctrl_rst_dat[19][14] , \sa_ctrl_rst_dat[19].r.part0[14] );
tran (\sa_ctrl_rst_dat[19][14] , \sa_ctrl_rst_dat[19].f.spare[9] );
tran (\sa_ctrl_rst_dat[19][15] , \sa_ctrl_rst_dat[19].r.part0[15] );
tran (\sa_ctrl_rst_dat[19][15] , \sa_ctrl_rst_dat[19].f.spare[10] );
tran (\sa_ctrl_rst_dat[19][16] , \sa_ctrl_rst_dat[19].r.part0[16] );
tran (\sa_ctrl_rst_dat[19][16] , \sa_ctrl_rst_dat[19].f.spare[11] );
tran (\sa_ctrl_rst_dat[19][17] , \sa_ctrl_rst_dat[19].r.part0[17] );
tran (\sa_ctrl_rst_dat[19][17] , \sa_ctrl_rst_dat[19].f.spare[12] );
tran (\sa_ctrl_rst_dat[19][18] , \sa_ctrl_rst_dat[19].r.part0[18] );
tran (\sa_ctrl_rst_dat[19][18] , \sa_ctrl_rst_dat[19].f.spare[13] );
tran (\sa_ctrl_rst_dat[19][19] , \sa_ctrl_rst_dat[19].r.part0[19] );
tran (\sa_ctrl_rst_dat[19][19] , \sa_ctrl_rst_dat[19].f.spare[14] );
tran (\sa_ctrl_rst_dat[19][20] , \sa_ctrl_rst_dat[19].r.part0[20] );
tran (\sa_ctrl_rst_dat[19][20] , \sa_ctrl_rst_dat[19].f.spare[15] );
tran (\sa_ctrl_rst_dat[19][21] , \sa_ctrl_rst_dat[19].r.part0[21] );
tran (\sa_ctrl_rst_dat[19][21] , \sa_ctrl_rst_dat[19].f.spare[16] );
tran (\sa_ctrl_rst_dat[19][22] , \sa_ctrl_rst_dat[19].r.part0[22] );
tran (\sa_ctrl_rst_dat[19][22] , \sa_ctrl_rst_dat[19].f.spare[17] );
tran (\sa_ctrl_rst_dat[19][23] , \sa_ctrl_rst_dat[19].r.part0[23] );
tran (\sa_ctrl_rst_dat[19][23] , \sa_ctrl_rst_dat[19].f.spare[18] );
tran (\sa_ctrl_rst_dat[19][24] , \sa_ctrl_rst_dat[19].r.part0[24] );
tran (\sa_ctrl_rst_dat[19][24] , \sa_ctrl_rst_dat[19].f.spare[19] );
tran (\sa_ctrl_rst_dat[19][25] , \sa_ctrl_rst_dat[19].r.part0[25] );
tran (\sa_ctrl_rst_dat[19][25] , \sa_ctrl_rst_dat[19].f.spare[20] );
tran (\sa_ctrl_rst_dat[19][26] , \sa_ctrl_rst_dat[19].r.part0[26] );
tran (\sa_ctrl_rst_dat[19][26] , \sa_ctrl_rst_dat[19].f.spare[21] );
tran (\sa_ctrl_rst_dat[19][27] , \sa_ctrl_rst_dat[19].r.part0[27] );
tran (\sa_ctrl_rst_dat[19][27] , \sa_ctrl_rst_dat[19].f.spare[22] );
tran (\sa_ctrl_rst_dat[19][28] , \sa_ctrl_rst_dat[19].r.part0[28] );
tran (\sa_ctrl_rst_dat[19][28] , \sa_ctrl_rst_dat[19].f.spare[23] );
tran (\sa_ctrl_rst_dat[19][29] , \sa_ctrl_rst_dat[19].r.part0[29] );
tran (\sa_ctrl_rst_dat[19][29] , \sa_ctrl_rst_dat[19].f.spare[24] );
tran (\sa_ctrl_rst_dat[19][30] , \sa_ctrl_rst_dat[19].r.part0[30] );
tran (\sa_ctrl_rst_dat[19][30] , \sa_ctrl_rst_dat[19].f.spare[25] );
tran (\sa_ctrl_rst_dat[19][31] , \sa_ctrl_rst_dat[19].r.part0[31] );
tran (\sa_ctrl_rst_dat[19][31] , \sa_ctrl_rst_dat[19].f.spare[26] );
tran (\sa_ctrl_rst_dat[20][0] , \sa_ctrl_rst_dat[20].r.part0[0] );
tran (\sa_ctrl_rst_dat[20][0] , \sa_ctrl_rst_dat[20].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[20][1] , \sa_ctrl_rst_dat[20].r.part0[1] );
tran (\sa_ctrl_rst_dat[20][1] , \sa_ctrl_rst_dat[20].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[20][2] , \sa_ctrl_rst_dat[20].r.part0[2] );
tran (\sa_ctrl_rst_dat[20][2] , \sa_ctrl_rst_dat[20].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[20][3] , \sa_ctrl_rst_dat[20].r.part0[3] );
tran (\sa_ctrl_rst_dat[20][3] , \sa_ctrl_rst_dat[20].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[20][4] , \sa_ctrl_rst_dat[20].r.part0[4] );
tran (\sa_ctrl_rst_dat[20][4] , \sa_ctrl_rst_dat[20].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[20][5] , \sa_ctrl_rst_dat[20].r.part0[5] );
tran (\sa_ctrl_rst_dat[20][5] , \sa_ctrl_rst_dat[20].f.spare[0] );
tran (\sa_ctrl_rst_dat[20][6] , \sa_ctrl_rst_dat[20].r.part0[6] );
tran (\sa_ctrl_rst_dat[20][6] , \sa_ctrl_rst_dat[20].f.spare[1] );
tran (\sa_ctrl_rst_dat[20][7] , \sa_ctrl_rst_dat[20].r.part0[7] );
tran (\sa_ctrl_rst_dat[20][7] , \sa_ctrl_rst_dat[20].f.spare[2] );
tran (\sa_ctrl_rst_dat[20][8] , \sa_ctrl_rst_dat[20].r.part0[8] );
tran (\sa_ctrl_rst_dat[20][8] , \sa_ctrl_rst_dat[20].f.spare[3] );
tran (\sa_ctrl_rst_dat[20][9] , \sa_ctrl_rst_dat[20].r.part0[9] );
tran (\sa_ctrl_rst_dat[20][9] , \sa_ctrl_rst_dat[20].f.spare[4] );
tran (\sa_ctrl_rst_dat[20][10] , \sa_ctrl_rst_dat[20].r.part0[10] );
tran (\sa_ctrl_rst_dat[20][10] , \sa_ctrl_rst_dat[20].f.spare[5] );
tran (\sa_ctrl_rst_dat[20][11] , \sa_ctrl_rst_dat[20].r.part0[11] );
tran (\sa_ctrl_rst_dat[20][11] , \sa_ctrl_rst_dat[20].f.spare[6] );
tran (\sa_ctrl_rst_dat[20][12] , \sa_ctrl_rst_dat[20].r.part0[12] );
tran (\sa_ctrl_rst_dat[20][12] , \sa_ctrl_rst_dat[20].f.spare[7] );
tran (\sa_ctrl_rst_dat[20][13] , \sa_ctrl_rst_dat[20].r.part0[13] );
tran (\sa_ctrl_rst_dat[20][13] , \sa_ctrl_rst_dat[20].f.spare[8] );
tran (\sa_ctrl_rst_dat[20][14] , \sa_ctrl_rst_dat[20].r.part0[14] );
tran (\sa_ctrl_rst_dat[20][14] , \sa_ctrl_rst_dat[20].f.spare[9] );
tran (\sa_ctrl_rst_dat[20][15] , \sa_ctrl_rst_dat[20].r.part0[15] );
tran (\sa_ctrl_rst_dat[20][15] , \sa_ctrl_rst_dat[20].f.spare[10] );
tran (\sa_ctrl_rst_dat[20][16] , \sa_ctrl_rst_dat[20].r.part0[16] );
tran (\sa_ctrl_rst_dat[20][16] , \sa_ctrl_rst_dat[20].f.spare[11] );
tran (\sa_ctrl_rst_dat[20][17] , \sa_ctrl_rst_dat[20].r.part0[17] );
tran (\sa_ctrl_rst_dat[20][17] , \sa_ctrl_rst_dat[20].f.spare[12] );
tran (\sa_ctrl_rst_dat[20][18] , \sa_ctrl_rst_dat[20].r.part0[18] );
tran (\sa_ctrl_rst_dat[20][18] , \sa_ctrl_rst_dat[20].f.spare[13] );
tran (\sa_ctrl_rst_dat[20][19] , \sa_ctrl_rst_dat[20].r.part0[19] );
tran (\sa_ctrl_rst_dat[20][19] , \sa_ctrl_rst_dat[20].f.spare[14] );
tran (\sa_ctrl_rst_dat[20][20] , \sa_ctrl_rst_dat[20].r.part0[20] );
tran (\sa_ctrl_rst_dat[20][20] , \sa_ctrl_rst_dat[20].f.spare[15] );
tran (\sa_ctrl_rst_dat[20][21] , \sa_ctrl_rst_dat[20].r.part0[21] );
tran (\sa_ctrl_rst_dat[20][21] , \sa_ctrl_rst_dat[20].f.spare[16] );
tran (\sa_ctrl_rst_dat[20][22] , \sa_ctrl_rst_dat[20].r.part0[22] );
tran (\sa_ctrl_rst_dat[20][22] , \sa_ctrl_rst_dat[20].f.spare[17] );
tran (\sa_ctrl_rst_dat[20][23] , \sa_ctrl_rst_dat[20].r.part0[23] );
tran (\sa_ctrl_rst_dat[20][23] , \sa_ctrl_rst_dat[20].f.spare[18] );
tran (\sa_ctrl_rst_dat[20][24] , \sa_ctrl_rst_dat[20].r.part0[24] );
tran (\sa_ctrl_rst_dat[20][24] , \sa_ctrl_rst_dat[20].f.spare[19] );
tran (\sa_ctrl_rst_dat[20][25] , \sa_ctrl_rst_dat[20].r.part0[25] );
tran (\sa_ctrl_rst_dat[20][25] , \sa_ctrl_rst_dat[20].f.spare[20] );
tran (\sa_ctrl_rst_dat[20][26] , \sa_ctrl_rst_dat[20].r.part0[26] );
tran (\sa_ctrl_rst_dat[20][26] , \sa_ctrl_rst_dat[20].f.spare[21] );
tran (\sa_ctrl_rst_dat[20][27] , \sa_ctrl_rst_dat[20].r.part0[27] );
tran (\sa_ctrl_rst_dat[20][27] , \sa_ctrl_rst_dat[20].f.spare[22] );
tran (\sa_ctrl_rst_dat[20][28] , \sa_ctrl_rst_dat[20].r.part0[28] );
tran (\sa_ctrl_rst_dat[20][28] , \sa_ctrl_rst_dat[20].f.spare[23] );
tran (\sa_ctrl_rst_dat[20][29] , \sa_ctrl_rst_dat[20].r.part0[29] );
tran (\sa_ctrl_rst_dat[20][29] , \sa_ctrl_rst_dat[20].f.spare[24] );
tran (\sa_ctrl_rst_dat[20][30] , \sa_ctrl_rst_dat[20].r.part0[30] );
tran (\sa_ctrl_rst_dat[20][30] , \sa_ctrl_rst_dat[20].f.spare[25] );
tran (\sa_ctrl_rst_dat[20][31] , \sa_ctrl_rst_dat[20].r.part0[31] );
tran (\sa_ctrl_rst_dat[20][31] , \sa_ctrl_rst_dat[20].f.spare[26] );
tran (\sa_ctrl_rst_dat[21][0] , \sa_ctrl_rst_dat[21].r.part0[0] );
tran (\sa_ctrl_rst_dat[21][0] , \sa_ctrl_rst_dat[21].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[21][1] , \sa_ctrl_rst_dat[21].r.part0[1] );
tran (\sa_ctrl_rst_dat[21][1] , \sa_ctrl_rst_dat[21].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[21][2] , \sa_ctrl_rst_dat[21].r.part0[2] );
tran (\sa_ctrl_rst_dat[21][2] , \sa_ctrl_rst_dat[21].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[21][3] , \sa_ctrl_rst_dat[21].r.part0[3] );
tran (\sa_ctrl_rst_dat[21][3] , \sa_ctrl_rst_dat[21].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[21][4] , \sa_ctrl_rst_dat[21].r.part0[4] );
tran (\sa_ctrl_rst_dat[21][4] , \sa_ctrl_rst_dat[21].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[21][5] , \sa_ctrl_rst_dat[21].r.part0[5] );
tran (\sa_ctrl_rst_dat[21][5] , \sa_ctrl_rst_dat[21].f.spare[0] );
tran (\sa_ctrl_rst_dat[21][6] , \sa_ctrl_rst_dat[21].r.part0[6] );
tran (\sa_ctrl_rst_dat[21][6] , \sa_ctrl_rst_dat[21].f.spare[1] );
tran (\sa_ctrl_rst_dat[21][7] , \sa_ctrl_rst_dat[21].r.part0[7] );
tran (\sa_ctrl_rst_dat[21][7] , \sa_ctrl_rst_dat[21].f.spare[2] );
tran (\sa_ctrl_rst_dat[21][8] , \sa_ctrl_rst_dat[21].r.part0[8] );
tran (\sa_ctrl_rst_dat[21][8] , \sa_ctrl_rst_dat[21].f.spare[3] );
tran (\sa_ctrl_rst_dat[21][9] , \sa_ctrl_rst_dat[21].r.part0[9] );
tran (\sa_ctrl_rst_dat[21][9] , \sa_ctrl_rst_dat[21].f.spare[4] );
tran (\sa_ctrl_rst_dat[21][10] , \sa_ctrl_rst_dat[21].r.part0[10] );
tran (\sa_ctrl_rst_dat[21][10] , \sa_ctrl_rst_dat[21].f.spare[5] );
tran (\sa_ctrl_rst_dat[21][11] , \sa_ctrl_rst_dat[21].r.part0[11] );
tran (\sa_ctrl_rst_dat[21][11] , \sa_ctrl_rst_dat[21].f.spare[6] );
tran (\sa_ctrl_rst_dat[21][12] , \sa_ctrl_rst_dat[21].r.part0[12] );
tran (\sa_ctrl_rst_dat[21][12] , \sa_ctrl_rst_dat[21].f.spare[7] );
tran (\sa_ctrl_rst_dat[21][13] , \sa_ctrl_rst_dat[21].r.part0[13] );
tran (\sa_ctrl_rst_dat[21][13] , \sa_ctrl_rst_dat[21].f.spare[8] );
tran (\sa_ctrl_rst_dat[21][14] , \sa_ctrl_rst_dat[21].r.part0[14] );
tran (\sa_ctrl_rst_dat[21][14] , \sa_ctrl_rst_dat[21].f.spare[9] );
tran (\sa_ctrl_rst_dat[21][15] , \sa_ctrl_rst_dat[21].r.part0[15] );
tran (\sa_ctrl_rst_dat[21][15] , \sa_ctrl_rst_dat[21].f.spare[10] );
tran (\sa_ctrl_rst_dat[21][16] , \sa_ctrl_rst_dat[21].r.part0[16] );
tran (\sa_ctrl_rst_dat[21][16] , \sa_ctrl_rst_dat[21].f.spare[11] );
tran (\sa_ctrl_rst_dat[21][17] , \sa_ctrl_rst_dat[21].r.part0[17] );
tran (\sa_ctrl_rst_dat[21][17] , \sa_ctrl_rst_dat[21].f.spare[12] );
tran (\sa_ctrl_rst_dat[21][18] , \sa_ctrl_rst_dat[21].r.part0[18] );
tran (\sa_ctrl_rst_dat[21][18] , \sa_ctrl_rst_dat[21].f.spare[13] );
tran (\sa_ctrl_rst_dat[21][19] , \sa_ctrl_rst_dat[21].r.part0[19] );
tran (\sa_ctrl_rst_dat[21][19] , \sa_ctrl_rst_dat[21].f.spare[14] );
tran (\sa_ctrl_rst_dat[21][20] , \sa_ctrl_rst_dat[21].r.part0[20] );
tran (\sa_ctrl_rst_dat[21][20] , \sa_ctrl_rst_dat[21].f.spare[15] );
tran (\sa_ctrl_rst_dat[21][21] , \sa_ctrl_rst_dat[21].r.part0[21] );
tran (\sa_ctrl_rst_dat[21][21] , \sa_ctrl_rst_dat[21].f.spare[16] );
tran (\sa_ctrl_rst_dat[21][22] , \sa_ctrl_rst_dat[21].r.part0[22] );
tran (\sa_ctrl_rst_dat[21][22] , \sa_ctrl_rst_dat[21].f.spare[17] );
tran (\sa_ctrl_rst_dat[21][23] , \sa_ctrl_rst_dat[21].r.part0[23] );
tran (\sa_ctrl_rst_dat[21][23] , \sa_ctrl_rst_dat[21].f.spare[18] );
tran (\sa_ctrl_rst_dat[21][24] , \sa_ctrl_rst_dat[21].r.part0[24] );
tran (\sa_ctrl_rst_dat[21][24] , \sa_ctrl_rst_dat[21].f.spare[19] );
tran (\sa_ctrl_rst_dat[21][25] , \sa_ctrl_rst_dat[21].r.part0[25] );
tran (\sa_ctrl_rst_dat[21][25] , \sa_ctrl_rst_dat[21].f.spare[20] );
tran (\sa_ctrl_rst_dat[21][26] , \sa_ctrl_rst_dat[21].r.part0[26] );
tran (\sa_ctrl_rst_dat[21][26] , \sa_ctrl_rst_dat[21].f.spare[21] );
tran (\sa_ctrl_rst_dat[21][27] , \sa_ctrl_rst_dat[21].r.part0[27] );
tran (\sa_ctrl_rst_dat[21][27] , \sa_ctrl_rst_dat[21].f.spare[22] );
tran (\sa_ctrl_rst_dat[21][28] , \sa_ctrl_rst_dat[21].r.part0[28] );
tran (\sa_ctrl_rst_dat[21][28] , \sa_ctrl_rst_dat[21].f.spare[23] );
tran (\sa_ctrl_rst_dat[21][29] , \sa_ctrl_rst_dat[21].r.part0[29] );
tran (\sa_ctrl_rst_dat[21][29] , \sa_ctrl_rst_dat[21].f.spare[24] );
tran (\sa_ctrl_rst_dat[21][30] , \sa_ctrl_rst_dat[21].r.part0[30] );
tran (\sa_ctrl_rst_dat[21][30] , \sa_ctrl_rst_dat[21].f.spare[25] );
tran (\sa_ctrl_rst_dat[21][31] , \sa_ctrl_rst_dat[21].r.part0[31] );
tran (\sa_ctrl_rst_dat[21][31] , \sa_ctrl_rst_dat[21].f.spare[26] );
tran (\sa_ctrl_rst_dat[22][0] , \sa_ctrl_rst_dat[22].r.part0[0] );
tran (\sa_ctrl_rst_dat[22][0] , \sa_ctrl_rst_dat[22].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[22][1] , \sa_ctrl_rst_dat[22].r.part0[1] );
tran (\sa_ctrl_rst_dat[22][1] , \sa_ctrl_rst_dat[22].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[22][2] , \sa_ctrl_rst_dat[22].r.part0[2] );
tran (\sa_ctrl_rst_dat[22][2] , \sa_ctrl_rst_dat[22].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[22][3] , \sa_ctrl_rst_dat[22].r.part0[3] );
tran (\sa_ctrl_rst_dat[22][3] , \sa_ctrl_rst_dat[22].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[22][4] , \sa_ctrl_rst_dat[22].r.part0[4] );
tran (\sa_ctrl_rst_dat[22][4] , \sa_ctrl_rst_dat[22].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[22][5] , \sa_ctrl_rst_dat[22].r.part0[5] );
tran (\sa_ctrl_rst_dat[22][5] , \sa_ctrl_rst_dat[22].f.spare[0] );
tran (\sa_ctrl_rst_dat[22][6] , \sa_ctrl_rst_dat[22].r.part0[6] );
tran (\sa_ctrl_rst_dat[22][6] , \sa_ctrl_rst_dat[22].f.spare[1] );
tran (\sa_ctrl_rst_dat[22][7] , \sa_ctrl_rst_dat[22].r.part0[7] );
tran (\sa_ctrl_rst_dat[22][7] , \sa_ctrl_rst_dat[22].f.spare[2] );
tran (\sa_ctrl_rst_dat[22][8] , \sa_ctrl_rst_dat[22].r.part0[8] );
tran (\sa_ctrl_rst_dat[22][8] , \sa_ctrl_rst_dat[22].f.spare[3] );
tran (\sa_ctrl_rst_dat[22][9] , \sa_ctrl_rst_dat[22].r.part0[9] );
tran (\sa_ctrl_rst_dat[22][9] , \sa_ctrl_rst_dat[22].f.spare[4] );
tran (\sa_ctrl_rst_dat[22][10] , \sa_ctrl_rst_dat[22].r.part0[10] );
tran (\sa_ctrl_rst_dat[22][10] , \sa_ctrl_rst_dat[22].f.spare[5] );
tran (\sa_ctrl_rst_dat[22][11] , \sa_ctrl_rst_dat[22].r.part0[11] );
tran (\sa_ctrl_rst_dat[22][11] , \sa_ctrl_rst_dat[22].f.spare[6] );
tran (\sa_ctrl_rst_dat[22][12] , \sa_ctrl_rst_dat[22].r.part0[12] );
tran (\sa_ctrl_rst_dat[22][12] , \sa_ctrl_rst_dat[22].f.spare[7] );
tran (\sa_ctrl_rst_dat[22][13] , \sa_ctrl_rst_dat[22].r.part0[13] );
tran (\sa_ctrl_rst_dat[22][13] , \sa_ctrl_rst_dat[22].f.spare[8] );
tran (\sa_ctrl_rst_dat[22][14] , \sa_ctrl_rst_dat[22].r.part0[14] );
tran (\sa_ctrl_rst_dat[22][14] , \sa_ctrl_rst_dat[22].f.spare[9] );
tran (\sa_ctrl_rst_dat[22][15] , \sa_ctrl_rst_dat[22].r.part0[15] );
tran (\sa_ctrl_rst_dat[22][15] , \sa_ctrl_rst_dat[22].f.spare[10] );
tran (\sa_ctrl_rst_dat[22][16] , \sa_ctrl_rst_dat[22].r.part0[16] );
tran (\sa_ctrl_rst_dat[22][16] , \sa_ctrl_rst_dat[22].f.spare[11] );
tran (\sa_ctrl_rst_dat[22][17] , \sa_ctrl_rst_dat[22].r.part0[17] );
tran (\sa_ctrl_rst_dat[22][17] , \sa_ctrl_rst_dat[22].f.spare[12] );
tran (\sa_ctrl_rst_dat[22][18] , \sa_ctrl_rst_dat[22].r.part0[18] );
tran (\sa_ctrl_rst_dat[22][18] , \sa_ctrl_rst_dat[22].f.spare[13] );
tran (\sa_ctrl_rst_dat[22][19] , \sa_ctrl_rst_dat[22].r.part0[19] );
tran (\sa_ctrl_rst_dat[22][19] , \sa_ctrl_rst_dat[22].f.spare[14] );
tran (\sa_ctrl_rst_dat[22][20] , \sa_ctrl_rst_dat[22].r.part0[20] );
tran (\sa_ctrl_rst_dat[22][20] , \sa_ctrl_rst_dat[22].f.spare[15] );
tran (\sa_ctrl_rst_dat[22][21] , \sa_ctrl_rst_dat[22].r.part0[21] );
tran (\sa_ctrl_rst_dat[22][21] , \sa_ctrl_rst_dat[22].f.spare[16] );
tran (\sa_ctrl_rst_dat[22][22] , \sa_ctrl_rst_dat[22].r.part0[22] );
tran (\sa_ctrl_rst_dat[22][22] , \sa_ctrl_rst_dat[22].f.spare[17] );
tran (\sa_ctrl_rst_dat[22][23] , \sa_ctrl_rst_dat[22].r.part0[23] );
tran (\sa_ctrl_rst_dat[22][23] , \sa_ctrl_rst_dat[22].f.spare[18] );
tran (\sa_ctrl_rst_dat[22][24] , \sa_ctrl_rst_dat[22].r.part0[24] );
tran (\sa_ctrl_rst_dat[22][24] , \sa_ctrl_rst_dat[22].f.spare[19] );
tran (\sa_ctrl_rst_dat[22][25] , \sa_ctrl_rst_dat[22].r.part0[25] );
tran (\sa_ctrl_rst_dat[22][25] , \sa_ctrl_rst_dat[22].f.spare[20] );
tran (\sa_ctrl_rst_dat[22][26] , \sa_ctrl_rst_dat[22].r.part0[26] );
tran (\sa_ctrl_rst_dat[22][26] , \sa_ctrl_rst_dat[22].f.spare[21] );
tran (\sa_ctrl_rst_dat[22][27] , \sa_ctrl_rst_dat[22].r.part0[27] );
tran (\sa_ctrl_rst_dat[22][27] , \sa_ctrl_rst_dat[22].f.spare[22] );
tran (\sa_ctrl_rst_dat[22][28] , \sa_ctrl_rst_dat[22].r.part0[28] );
tran (\sa_ctrl_rst_dat[22][28] , \sa_ctrl_rst_dat[22].f.spare[23] );
tran (\sa_ctrl_rst_dat[22][29] , \sa_ctrl_rst_dat[22].r.part0[29] );
tran (\sa_ctrl_rst_dat[22][29] , \sa_ctrl_rst_dat[22].f.spare[24] );
tran (\sa_ctrl_rst_dat[22][30] , \sa_ctrl_rst_dat[22].r.part0[30] );
tran (\sa_ctrl_rst_dat[22][30] , \sa_ctrl_rst_dat[22].f.spare[25] );
tran (\sa_ctrl_rst_dat[22][31] , \sa_ctrl_rst_dat[22].r.part0[31] );
tran (\sa_ctrl_rst_dat[22][31] , \sa_ctrl_rst_dat[22].f.spare[26] );
tran (\sa_ctrl_rst_dat[23][0] , \sa_ctrl_rst_dat[23].r.part0[0] );
tran (\sa_ctrl_rst_dat[23][0] , \sa_ctrl_rst_dat[23].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[23][1] , \sa_ctrl_rst_dat[23].r.part0[1] );
tran (\sa_ctrl_rst_dat[23][1] , \sa_ctrl_rst_dat[23].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[23][2] , \sa_ctrl_rst_dat[23].r.part0[2] );
tran (\sa_ctrl_rst_dat[23][2] , \sa_ctrl_rst_dat[23].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[23][3] , \sa_ctrl_rst_dat[23].r.part0[3] );
tran (\sa_ctrl_rst_dat[23][3] , \sa_ctrl_rst_dat[23].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[23][4] , \sa_ctrl_rst_dat[23].r.part0[4] );
tran (\sa_ctrl_rst_dat[23][4] , \sa_ctrl_rst_dat[23].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[23][5] , \sa_ctrl_rst_dat[23].r.part0[5] );
tran (\sa_ctrl_rst_dat[23][5] , \sa_ctrl_rst_dat[23].f.spare[0] );
tran (\sa_ctrl_rst_dat[23][6] , \sa_ctrl_rst_dat[23].r.part0[6] );
tran (\sa_ctrl_rst_dat[23][6] , \sa_ctrl_rst_dat[23].f.spare[1] );
tran (\sa_ctrl_rst_dat[23][7] , \sa_ctrl_rst_dat[23].r.part0[7] );
tran (\sa_ctrl_rst_dat[23][7] , \sa_ctrl_rst_dat[23].f.spare[2] );
tran (\sa_ctrl_rst_dat[23][8] , \sa_ctrl_rst_dat[23].r.part0[8] );
tran (\sa_ctrl_rst_dat[23][8] , \sa_ctrl_rst_dat[23].f.spare[3] );
tran (\sa_ctrl_rst_dat[23][9] , \sa_ctrl_rst_dat[23].r.part0[9] );
tran (\sa_ctrl_rst_dat[23][9] , \sa_ctrl_rst_dat[23].f.spare[4] );
tran (\sa_ctrl_rst_dat[23][10] , \sa_ctrl_rst_dat[23].r.part0[10] );
tran (\sa_ctrl_rst_dat[23][10] , \sa_ctrl_rst_dat[23].f.spare[5] );
tran (\sa_ctrl_rst_dat[23][11] , \sa_ctrl_rst_dat[23].r.part0[11] );
tran (\sa_ctrl_rst_dat[23][11] , \sa_ctrl_rst_dat[23].f.spare[6] );
tran (\sa_ctrl_rst_dat[23][12] , \sa_ctrl_rst_dat[23].r.part0[12] );
tran (\sa_ctrl_rst_dat[23][12] , \sa_ctrl_rst_dat[23].f.spare[7] );
tran (\sa_ctrl_rst_dat[23][13] , \sa_ctrl_rst_dat[23].r.part0[13] );
tran (\sa_ctrl_rst_dat[23][13] , \sa_ctrl_rst_dat[23].f.spare[8] );
tran (\sa_ctrl_rst_dat[23][14] , \sa_ctrl_rst_dat[23].r.part0[14] );
tran (\sa_ctrl_rst_dat[23][14] , \sa_ctrl_rst_dat[23].f.spare[9] );
tran (\sa_ctrl_rst_dat[23][15] , \sa_ctrl_rst_dat[23].r.part0[15] );
tran (\sa_ctrl_rst_dat[23][15] , \sa_ctrl_rst_dat[23].f.spare[10] );
tran (\sa_ctrl_rst_dat[23][16] , \sa_ctrl_rst_dat[23].r.part0[16] );
tran (\sa_ctrl_rst_dat[23][16] , \sa_ctrl_rst_dat[23].f.spare[11] );
tran (\sa_ctrl_rst_dat[23][17] , \sa_ctrl_rst_dat[23].r.part0[17] );
tran (\sa_ctrl_rst_dat[23][17] , \sa_ctrl_rst_dat[23].f.spare[12] );
tran (\sa_ctrl_rst_dat[23][18] , \sa_ctrl_rst_dat[23].r.part0[18] );
tran (\sa_ctrl_rst_dat[23][18] , \sa_ctrl_rst_dat[23].f.spare[13] );
tran (\sa_ctrl_rst_dat[23][19] , \sa_ctrl_rst_dat[23].r.part0[19] );
tran (\sa_ctrl_rst_dat[23][19] , \sa_ctrl_rst_dat[23].f.spare[14] );
tran (\sa_ctrl_rst_dat[23][20] , \sa_ctrl_rst_dat[23].r.part0[20] );
tran (\sa_ctrl_rst_dat[23][20] , \sa_ctrl_rst_dat[23].f.spare[15] );
tran (\sa_ctrl_rst_dat[23][21] , \sa_ctrl_rst_dat[23].r.part0[21] );
tran (\sa_ctrl_rst_dat[23][21] , \sa_ctrl_rst_dat[23].f.spare[16] );
tran (\sa_ctrl_rst_dat[23][22] , \sa_ctrl_rst_dat[23].r.part0[22] );
tran (\sa_ctrl_rst_dat[23][22] , \sa_ctrl_rst_dat[23].f.spare[17] );
tran (\sa_ctrl_rst_dat[23][23] , \sa_ctrl_rst_dat[23].r.part0[23] );
tran (\sa_ctrl_rst_dat[23][23] , \sa_ctrl_rst_dat[23].f.spare[18] );
tran (\sa_ctrl_rst_dat[23][24] , \sa_ctrl_rst_dat[23].r.part0[24] );
tran (\sa_ctrl_rst_dat[23][24] , \sa_ctrl_rst_dat[23].f.spare[19] );
tran (\sa_ctrl_rst_dat[23][25] , \sa_ctrl_rst_dat[23].r.part0[25] );
tran (\sa_ctrl_rst_dat[23][25] , \sa_ctrl_rst_dat[23].f.spare[20] );
tran (\sa_ctrl_rst_dat[23][26] , \sa_ctrl_rst_dat[23].r.part0[26] );
tran (\sa_ctrl_rst_dat[23][26] , \sa_ctrl_rst_dat[23].f.spare[21] );
tran (\sa_ctrl_rst_dat[23][27] , \sa_ctrl_rst_dat[23].r.part0[27] );
tran (\sa_ctrl_rst_dat[23][27] , \sa_ctrl_rst_dat[23].f.spare[22] );
tran (\sa_ctrl_rst_dat[23][28] , \sa_ctrl_rst_dat[23].r.part0[28] );
tran (\sa_ctrl_rst_dat[23][28] , \sa_ctrl_rst_dat[23].f.spare[23] );
tran (\sa_ctrl_rst_dat[23][29] , \sa_ctrl_rst_dat[23].r.part0[29] );
tran (\sa_ctrl_rst_dat[23][29] , \sa_ctrl_rst_dat[23].f.spare[24] );
tran (\sa_ctrl_rst_dat[23][30] , \sa_ctrl_rst_dat[23].r.part0[30] );
tran (\sa_ctrl_rst_dat[23][30] , \sa_ctrl_rst_dat[23].f.spare[25] );
tran (\sa_ctrl_rst_dat[23][31] , \sa_ctrl_rst_dat[23].r.part0[31] );
tran (\sa_ctrl_rst_dat[23][31] , \sa_ctrl_rst_dat[23].f.spare[26] );
tran (\sa_ctrl_rst_dat[24][0] , \sa_ctrl_rst_dat[24].r.part0[0] );
tran (\sa_ctrl_rst_dat[24][0] , \sa_ctrl_rst_dat[24].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[24][1] , \sa_ctrl_rst_dat[24].r.part0[1] );
tran (\sa_ctrl_rst_dat[24][1] , \sa_ctrl_rst_dat[24].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[24][2] , \sa_ctrl_rst_dat[24].r.part0[2] );
tran (\sa_ctrl_rst_dat[24][2] , \sa_ctrl_rst_dat[24].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[24][3] , \sa_ctrl_rst_dat[24].r.part0[3] );
tran (\sa_ctrl_rst_dat[24][3] , \sa_ctrl_rst_dat[24].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[24][4] , \sa_ctrl_rst_dat[24].r.part0[4] );
tran (\sa_ctrl_rst_dat[24][4] , \sa_ctrl_rst_dat[24].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[24][5] , \sa_ctrl_rst_dat[24].r.part0[5] );
tran (\sa_ctrl_rst_dat[24][5] , \sa_ctrl_rst_dat[24].f.spare[0] );
tran (\sa_ctrl_rst_dat[24][6] , \sa_ctrl_rst_dat[24].r.part0[6] );
tran (\sa_ctrl_rst_dat[24][6] , \sa_ctrl_rst_dat[24].f.spare[1] );
tran (\sa_ctrl_rst_dat[24][7] , \sa_ctrl_rst_dat[24].r.part0[7] );
tran (\sa_ctrl_rst_dat[24][7] , \sa_ctrl_rst_dat[24].f.spare[2] );
tran (\sa_ctrl_rst_dat[24][8] , \sa_ctrl_rst_dat[24].r.part0[8] );
tran (\sa_ctrl_rst_dat[24][8] , \sa_ctrl_rst_dat[24].f.spare[3] );
tran (\sa_ctrl_rst_dat[24][9] , \sa_ctrl_rst_dat[24].r.part0[9] );
tran (\sa_ctrl_rst_dat[24][9] , \sa_ctrl_rst_dat[24].f.spare[4] );
tran (\sa_ctrl_rst_dat[24][10] , \sa_ctrl_rst_dat[24].r.part0[10] );
tran (\sa_ctrl_rst_dat[24][10] , \sa_ctrl_rst_dat[24].f.spare[5] );
tran (\sa_ctrl_rst_dat[24][11] , \sa_ctrl_rst_dat[24].r.part0[11] );
tran (\sa_ctrl_rst_dat[24][11] , \sa_ctrl_rst_dat[24].f.spare[6] );
tran (\sa_ctrl_rst_dat[24][12] , \sa_ctrl_rst_dat[24].r.part0[12] );
tran (\sa_ctrl_rst_dat[24][12] , \sa_ctrl_rst_dat[24].f.spare[7] );
tran (\sa_ctrl_rst_dat[24][13] , \sa_ctrl_rst_dat[24].r.part0[13] );
tran (\sa_ctrl_rst_dat[24][13] , \sa_ctrl_rst_dat[24].f.spare[8] );
tran (\sa_ctrl_rst_dat[24][14] , \sa_ctrl_rst_dat[24].r.part0[14] );
tran (\sa_ctrl_rst_dat[24][14] , \sa_ctrl_rst_dat[24].f.spare[9] );
tran (\sa_ctrl_rst_dat[24][15] , \sa_ctrl_rst_dat[24].r.part0[15] );
tran (\sa_ctrl_rst_dat[24][15] , \sa_ctrl_rst_dat[24].f.spare[10] );
tran (\sa_ctrl_rst_dat[24][16] , \sa_ctrl_rst_dat[24].r.part0[16] );
tran (\sa_ctrl_rst_dat[24][16] , \sa_ctrl_rst_dat[24].f.spare[11] );
tran (\sa_ctrl_rst_dat[24][17] , \sa_ctrl_rst_dat[24].r.part0[17] );
tran (\sa_ctrl_rst_dat[24][17] , \sa_ctrl_rst_dat[24].f.spare[12] );
tran (\sa_ctrl_rst_dat[24][18] , \sa_ctrl_rst_dat[24].r.part0[18] );
tran (\sa_ctrl_rst_dat[24][18] , \sa_ctrl_rst_dat[24].f.spare[13] );
tran (\sa_ctrl_rst_dat[24][19] , \sa_ctrl_rst_dat[24].r.part0[19] );
tran (\sa_ctrl_rst_dat[24][19] , \sa_ctrl_rst_dat[24].f.spare[14] );
tran (\sa_ctrl_rst_dat[24][20] , \sa_ctrl_rst_dat[24].r.part0[20] );
tran (\sa_ctrl_rst_dat[24][20] , \sa_ctrl_rst_dat[24].f.spare[15] );
tran (\sa_ctrl_rst_dat[24][21] , \sa_ctrl_rst_dat[24].r.part0[21] );
tran (\sa_ctrl_rst_dat[24][21] , \sa_ctrl_rst_dat[24].f.spare[16] );
tran (\sa_ctrl_rst_dat[24][22] , \sa_ctrl_rst_dat[24].r.part0[22] );
tran (\sa_ctrl_rst_dat[24][22] , \sa_ctrl_rst_dat[24].f.spare[17] );
tran (\sa_ctrl_rst_dat[24][23] , \sa_ctrl_rst_dat[24].r.part0[23] );
tran (\sa_ctrl_rst_dat[24][23] , \sa_ctrl_rst_dat[24].f.spare[18] );
tran (\sa_ctrl_rst_dat[24][24] , \sa_ctrl_rst_dat[24].r.part0[24] );
tran (\sa_ctrl_rst_dat[24][24] , \sa_ctrl_rst_dat[24].f.spare[19] );
tran (\sa_ctrl_rst_dat[24][25] , \sa_ctrl_rst_dat[24].r.part0[25] );
tran (\sa_ctrl_rst_dat[24][25] , \sa_ctrl_rst_dat[24].f.spare[20] );
tran (\sa_ctrl_rst_dat[24][26] , \sa_ctrl_rst_dat[24].r.part0[26] );
tran (\sa_ctrl_rst_dat[24][26] , \sa_ctrl_rst_dat[24].f.spare[21] );
tran (\sa_ctrl_rst_dat[24][27] , \sa_ctrl_rst_dat[24].r.part0[27] );
tran (\sa_ctrl_rst_dat[24][27] , \sa_ctrl_rst_dat[24].f.spare[22] );
tran (\sa_ctrl_rst_dat[24][28] , \sa_ctrl_rst_dat[24].r.part0[28] );
tran (\sa_ctrl_rst_dat[24][28] , \sa_ctrl_rst_dat[24].f.spare[23] );
tran (\sa_ctrl_rst_dat[24][29] , \sa_ctrl_rst_dat[24].r.part0[29] );
tran (\sa_ctrl_rst_dat[24][29] , \sa_ctrl_rst_dat[24].f.spare[24] );
tran (\sa_ctrl_rst_dat[24][30] , \sa_ctrl_rst_dat[24].r.part0[30] );
tran (\sa_ctrl_rst_dat[24][30] , \sa_ctrl_rst_dat[24].f.spare[25] );
tran (\sa_ctrl_rst_dat[24][31] , \sa_ctrl_rst_dat[24].r.part0[31] );
tran (\sa_ctrl_rst_dat[24][31] , \sa_ctrl_rst_dat[24].f.spare[26] );
tran (\sa_ctrl_rst_dat[25][0] , \sa_ctrl_rst_dat[25].r.part0[0] );
tran (\sa_ctrl_rst_dat[25][0] , \sa_ctrl_rst_dat[25].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[25][1] , \sa_ctrl_rst_dat[25].r.part0[1] );
tran (\sa_ctrl_rst_dat[25][1] , \sa_ctrl_rst_dat[25].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[25][2] , \sa_ctrl_rst_dat[25].r.part0[2] );
tran (\sa_ctrl_rst_dat[25][2] , \sa_ctrl_rst_dat[25].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[25][3] , \sa_ctrl_rst_dat[25].r.part0[3] );
tran (\sa_ctrl_rst_dat[25][3] , \sa_ctrl_rst_dat[25].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[25][4] , \sa_ctrl_rst_dat[25].r.part0[4] );
tran (\sa_ctrl_rst_dat[25][4] , \sa_ctrl_rst_dat[25].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[25][5] , \sa_ctrl_rst_dat[25].r.part0[5] );
tran (\sa_ctrl_rst_dat[25][5] , \sa_ctrl_rst_dat[25].f.spare[0] );
tran (\sa_ctrl_rst_dat[25][6] , \sa_ctrl_rst_dat[25].r.part0[6] );
tran (\sa_ctrl_rst_dat[25][6] , \sa_ctrl_rst_dat[25].f.spare[1] );
tran (\sa_ctrl_rst_dat[25][7] , \sa_ctrl_rst_dat[25].r.part0[7] );
tran (\sa_ctrl_rst_dat[25][7] , \sa_ctrl_rst_dat[25].f.spare[2] );
tran (\sa_ctrl_rst_dat[25][8] , \sa_ctrl_rst_dat[25].r.part0[8] );
tran (\sa_ctrl_rst_dat[25][8] , \sa_ctrl_rst_dat[25].f.spare[3] );
tran (\sa_ctrl_rst_dat[25][9] , \sa_ctrl_rst_dat[25].r.part0[9] );
tran (\sa_ctrl_rst_dat[25][9] , \sa_ctrl_rst_dat[25].f.spare[4] );
tran (\sa_ctrl_rst_dat[25][10] , \sa_ctrl_rst_dat[25].r.part0[10] );
tran (\sa_ctrl_rst_dat[25][10] , \sa_ctrl_rst_dat[25].f.spare[5] );
tran (\sa_ctrl_rst_dat[25][11] , \sa_ctrl_rst_dat[25].r.part0[11] );
tran (\sa_ctrl_rst_dat[25][11] , \sa_ctrl_rst_dat[25].f.spare[6] );
tran (\sa_ctrl_rst_dat[25][12] , \sa_ctrl_rst_dat[25].r.part0[12] );
tran (\sa_ctrl_rst_dat[25][12] , \sa_ctrl_rst_dat[25].f.spare[7] );
tran (\sa_ctrl_rst_dat[25][13] , \sa_ctrl_rst_dat[25].r.part0[13] );
tran (\sa_ctrl_rst_dat[25][13] , \sa_ctrl_rst_dat[25].f.spare[8] );
tran (\sa_ctrl_rst_dat[25][14] , \sa_ctrl_rst_dat[25].r.part0[14] );
tran (\sa_ctrl_rst_dat[25][14] , \sa_ctrl_rst_dat[25].f.spare[9] );
tran (\sa_ctrl_rst_dat[25][15] , \sa_ctrl_rst_dat[25].r.part0[15] );
tran (\sa_ctrl_rst_dat[25][15] , \sa_ctrl_rst_dat[25].f.spare[10] );
tran (\sa_ctrl_rst_dat[25][16] , \sa_ctrl_rst_dat[25].r.part0[16] );
tran (\sa_ctrl_rst_dat[25][16] , \sa_ctrl_rst_dat[25].f.spare[11] );
tran (\sa_ctrl_rst_dat[25][17] , \sa_ctrl_rst_dat[25].r.part0[17] );
tran (\sa_ctrl_rst_dat[25][17] , \sa_ctrl_rst_dat[25].f.spare[12] );
tran (\sa_ctrl_rst_dat[25][18] , \sa_ctrl_rst_dat[25].r.part0[18] );
tran (\sa_ctrl_rst_dat[25][18] , \sa_ctrl_rst_dat[25].f.spare[13] );
tran (\sa_ctrl_rst_dat[25][19] , \sa_ctrl_rst_dat[25].r.part0[19] );
tran (\sa_ctrl_rst_dat[25][19] , \sa_ctrl_rst_dat[25].f.spare[14] );
tran (\sa_ctrl_rst_dat[25][20] , \sa_ctrl_rst_dat[25].r.part0[20] );
tran (\sa_ctrl_rst_dat[25][20] , \sa_ctrl_rst_dat[25].f.spare[15] );
tran (\sa_ctrl_rst_dat[25][21] , \sa_ctrl_rst_dat[25].r.part0[21] );
tran (\sa_ctrl_rst_dat[25][21] , \sa_ctrl_rst_dat[25].f.spare[16] );
tran (\sa_ctrl_rst_dat[25][22] , \sa_ctrl_rst_dat[25].r.part0[22] );
tran (\sa_ctrl_rst_dat[25][22] , \sa_ctrl_rst_dat[25].f.spare[17] );
tran (\sa_ctrl_rst_dat[25][23] , \sa_ctrl_rst_dat[25].r.part0[23] );
tran (\sa_ctrl_rst_dat[25][23] , \sa_ctrl_rst_dat[25].f.spare[18] );
tran (\sa_ctrl_rst_dat[25][24] , \sa_ctrl_rst_dat[25].r.part0[24] );
tran (\sa_ctrl_rst_dat[25][24] , \sa_ctrl_rst_dat[25].f.spare[19] );
tran (\sa_ctrl_rst_dat[25][25] , \sa_ctrl_rst_dat[25].r.part0[25] );
tran (\sa_ctrl_rst_dat[25][25] , \sa_ctrl_rst_dat[25].f.spare[20] );
tran (\sa_ctrl_rst_dat[25][26] , \sa_ctrl_rst_dat[25].r.part0[26] );
tran (\sa_ctrl_rst_dat[25][26] , \sa_ctrl_rst_dat[25].f.spare[21] );
tran (\sa_ctrl_rst_dat[25][27] , \sa_ctrl_rst_dat[25].r.part0[27] );
tran (\sa_ctrl_rst_dat[25][27] , \sa_ctrl_rst_dat[25].f.spare[22] );
tran (\sa_ctrl_rst_dat[25][28] , \sa_ctrl_rst_dat[25].r.part0[28] );
tran (\sa_ctrl_rst_dat[25][28] , \sa_ctrl_rst_dat[25].f.spare[23] );
tran (\sa_ctrl_rst_dat[25][29] , \sa_ctrl_rst_dat[25].r.part0[29] );
tran (\sa_ctrl_rst_dat[25][29] , \sa_ctrl_rst_dat[25].f.spare[24] );
tran (\sa_ctrl_rst_dat[25][30] , \sa_ctrl_rst_dat[25].r.part0[30] );
tran (\sa_ctrl_rst_dat[25][30] , \sa_ctrl_rst_dat[25].f.spare[25] );
tran (\sa_ctrl_rst_dat[25][31] , \sa_ctrl_rst_dat[25].r.part0[31] );
tran (\sa_ctrl_rst_dat[25][31] , \sa_ctrl_rst_dat[25].f.spare[26] );
tran (\sa_ctrl_rst_dat[26][0] , \sa_ctrl_rst_dat[26].r.part0[0] );
tran (\sa_ctrl_rst_dat[26][0] , \sa_ctrl_rst_dat[26].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[26][1] , \sa_ctrl_rst_dat[26].r.part0[1] );
tran (\sa_ctrl_rst_dat[26][1] , \sa_ctrl_rst_dat[26].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[26][2] , \sa_ctrl_rst_dat[26].r.part0[2] );
tran (\sa_ctrl_rst_dat[26][2] , \sa_ctrl_rst_dat[26].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[26][3] , \sa_ctrl_rst_dat[26].r.part0[3] );
tran (\sa_ctrl_rst_dat[26][3] , \sa_ctrl_rst_dat[26].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[26][4] , \sa_ctrl_rst_dat[26].r.part0[4] );
tran (\sa_ctrl_rst_dat[26][4] , \sa_ctrl_rst_dat[26].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[26][5] , \sa_ctrl_rst_dat[26].r.part0[5] );
tran (\sa_ctrl_rst_dat[26][5] , \sa_ctrl_rst_dat[26].f.spare[0] );
tran (\sa_ctrl_rst_dat[26][6] , \sa_ctrl_rst_dat[26].r.part0[6] );
tran (\sa_ctrl_rst_dat[26][6] , \sa_ctrl_rst_dat[26].f.spare[1] );
tran (\sa_ctrl_rst_dat[26][7] , \sa_ctrl_rst_dat[26].r.part0[7] );
tran (\sa_ctrl_rst_dat[26][7] , \sa_ctrl_rst_dat[26].f.spare[2] );
tran (\sa_ctrl_rst_dat[26][8] , \sa_ctrl_rst_dat[26].r.part0[8] );
tran (\sa_ctrl_rst_dat[26][8] , \sa_ctrl_rst_dat[26].f.spare[3] );
tran (\sa_ctrl_rst_dat[26][9] , \sa_ctrl_rst_dat[26].r.part0[9] );
tran (\sa_ctrl_rst_dat[26][9] , \sa_ctrl_rst_dat[26].f.spare[4] );
tran (\sa_ctrl_rst_dat[26][10] , \sa_ctrl_rst_dat[26].r.part0[10] );
tran (\sa_ctrl_rst_dat[26][10] , \sa_ctrl_rst_dat[26].f.spare[5] );
tran (\sa_ctrl_rst_dat[26][11] , \sa_ctrl_rst_dat[26].r.part0[11] );
tran (\sa_ctrl_rst_dat[26][11] , \sa_ctrl_rst_dat[26].f.spare[6] );
tran (\sa_ctrl_rst_dat[26][12] , \sa_ctrl_rst_dat[26].r.part0[12] );
tran (\sa_ctrl_rst_dat[26][12] , \sa_ctrl_rst_dat[26].f.spare[7] );
tran (\sa_ctrl_rst_dat[26][13] , \sa_ctrl_rst_dat[26].r.part0[13] );
tran (\sa_ctrl_rst_dat[26][13] , \sa_ctrl_rst_dat[26].f.spare[8] );
tran (\sa_ctrl_rst_dat[26][14] , \sa_ctrl_rst_dat[26].r.part0[14] );
tran (\sa_ctrl_rst_dat[26][14] , \sa_ctrl_rst_dat[26].f.spare[9] );
tran (\sa_ctrl_rst_dat[26][15] , \sa_ctrl_rst_dat[26].r.part0[15] );
tran (\sa_ctrl_rst_dat[26][15] , \sa_ctrl_rst_dat[26].f.spare[10] );
tran (\sa_ctrl_rst_dat[26][16] , \sa_ctrl_rst_dat[26].r.part0[16] );
tran (\sa_ctrl_rst_dat[26][16] , \sa_ctrl_rst_dat[26].f.spare[11] );
tran (\sa_ctrl_rst_dat[26][17] , \sa_ctrl_rst_dat[26].r.part0[17] );
tran (\sa_ctrl_rst_dat[26][17] , \sa_ctrl_rst_dat[26].f.spare[12] );
tran (\sa_ctrl_rst_dat[26][18] , \sa_ctrl_rst_dat[26].r.part0[18] );
tran (\sa_ctrl_rst_dat[26][18] , \sa_ctrl_rst_dat[26].f.spare[13] );
tran (\sa_ctrl_rst_dat[26][19] , \sa_ctrl_rst_dat[26].r.part0[19] );
tran (\sa_ctrl_rst_dat[26][19] , \sa_ctrl_rst_dat[26].f.spare[14] );
tran (\sa_ctrl_rst_dat[26][20] , \sa_ctrl_rst_dat[26].r.part0[20] );
tran (\sa_ctrl_rst_dat[26][20] , \sa_ctrl_rst_dat[26].f.spare[15] );
tran (\sa_ctrl_rst_dat[26][21] , \sa_ctrl_rst_dat[26].r.part0[21] );
tran (\sa_ctrl_rst_dat[26][21] , \sa_ctrl_rst_dat[26].f.spare[16] );
tran (\sa_ctrl_rst_dat[26][22] , \sa_ctrl_rst_dat[26].r.part0[22] );
tran (\sa_ctrl_rst_dat[26][22] , \sa_ctrl_rst_dat[26].f.spare[17] );
tran (\sa_ctrl_rst_dat[26][23] , \sa_ctrl_rst_dat[26].r.part0[23] );
tran (\sa_ctrl_rst_dat[26][23] , \sa_ctrl_rst_dat[26].f.spare[18] );
tran (\sa_ctrl_rst_dat[26][24] , \sa_ctrl_rst_dat[26].r.part0[24] );
tran (\sa_ctrl_rst_dat[26][24] , \sa_ctrl_rst_dat[26].f.spare[19] );
tran (\sa_ctrl_rst_dat[26][25] , \sa_ctrl_rst_dat[26].r.part0[25] );
tran (\sa_ctrl_rst_dat[26][25] , \sa_ctrl_rst_dat[26].f.spare[20] );
tran (\sa_ctrl_rst_dat[26][26] , \sa_ctrl_rst_dat[26].r.part0[26] );
tran (\sa_ctrl_rst_dat[26][26] , \sa_ctrl_rst_dat[26].f.spare[21] );
tran (\sa_ctrl_rst_dat[26][27] , \sa_ctrl_rst_dat[26].r.part0[27] );
tran (\sa_ctrl_rst_dat[26][27] , \sa_ctrl_rst_dat[26].f.spare[22] );
tran (\sa_ctrl_rst_dat[26][28] , \sa_ctrl_rst_dat[26].r.part0[28] );
tran (\sa_ctrl_rst_dat[26][28] , \sa_ctrl_rst_dat[26].f.spare[23] );
tran (\sa_ctrl_rst_dat[26][29] , \sa_ctrl_rst_dat[26].r.part0[29] );
tran (\sa_ctrl_rst_dat[26][29] , \sa_ctrl_rst_dat[26].f.spare[24] );
tran (\sa_ctrl_rst_dat[26][30] , \sa_ctrl_rst_dat[26].r.part0[30] );
tran (\sa_ctrl_rst_dat[26][30] , \sa_ctrl_rst_dat[26].f.spare[25] );
tran (\sa_ctrl_rst_dat[26][31] , \sa_ctrl_rst_dat[26].r.part0[31] );
tran (\sa_ctrl_rst_dat[26][31] , \sa_ctrl_rst_dat[26].f.spare[26] );
tran (\sa_ctrl_rst_dat[27][0] , \sa_ctrl_rst_dat[27].r.part0[0] );
tran (\sa_ctrl_rst_dat[27][0] , \sa_ctrl_rst_dat[27].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[27][1] , \sa_ctrl_rst_dat[27].r.part0[1] );
tran (\sa_ctrl_rst_dat[27][1] , \sa_ctrl_rst_dat[27].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[27][2] , \sa_ctrl_rst_dat[27].r.part0[2] );
tran (\sa_ctrl_rst_dat[27][2] , \sa_ctrl_rst_dat[27].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[27][3] , \sa_ctrl_rst_dat[27].r.part0[3] );
tran (\sa_ctrl_rst_dat[27][3] , \sa_ctrl_rst_dat[27].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[27][4] , \sa_ctrl_rst_dat[27].r.part0[4] );
tran (\sa_ctrl_rst_dat[27][4] , \sa_ctrl_rst_dat[27].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[27][5] , \sa_ctrl_rst_dat[27].r.part0[5] );
tran (\sa_ctrl_rst_dat[27][5] , \sa_ctrl_rst_dat[27].f.spare[0] );
tran (\sa_ctrl_rst_dat[27][6] , \sa_ctrl_rst_dat[27].r.part0[6] );
tran (\sa_ctrl_rst_dat[27][6] , \sa_ctrl_rst_dat[27].f.spare[1] );
tran (\sa_ctrl_rst_dat[27][7] , \sa_ctrl_rst_dat[27].r.part0[7] );
tran (\sa_ctrl_rst_dat[27][7] , \sa_ctrl_rst_dat[27].f.spare[2] );
tran (\sa_ctrl_rst_dat[27][8] , \sa_ctrl_rst_dat[27].r.part0[8] );
tran (\sa_ctrl_rst_dat[27][8] , \sa_ctrl_rst_dat[27].f.spare[3] );
tran (\sa_ctrl_rst_dat[27][9] , \sa_ctrl_rst_dat[27].r.part0[9] );
tran (\sa_ctrl_rst_dat[27][9] , \sa_ctrl_rst_dat[27].f.spare[4] );
tran (\sa_ctrl_rst_dat[27][10] , \sa_ctrl_rst_dat[27].r.part0[10] );
tran (\sa_ctrl_rst_dat[27][10] , \sa_ctrl_rst_dat[27].f.spare[5] );
tran (\sa_ctrl_rst_dat[27][11] , \sa_ctrl_rst_dat[27].r.part0[11] );
tran (\sa_ctrl_rst_dat[27][11] , \sa_ctrl_rst_dat[27].f.spare[6] );
tran (\sa_ctrl_rst_dat[27][12] , \sa_ctrl_rst_dat[27].r.part0[12] );
tran (\sa_ctrl_rst_dat[27][12] , \sa_ctrl_rst_dat[27].f.spare[7] );
tran (\sa_ctrl_rst_dat[27][13] , \sa_ctrl_rst_dat[27].r.part0[13] );
tran (\sa_ctrl_rst_dat[27][13] , \sa_ctrl_rst_dat[27].f.spare[8] );
tran (\sa_ctrl_rst_dat[27][14] , \sa_ctrl_rst_dat[27].r.part0[14] );
tran (\sa_ctrl_rst_dat[27][14] , \sa_ctrl_rst_dat[27].f.spare[9] );
tran (\sa_ctrl_rst_dat[27][15] , \sa_ctrl_rst_dat[27].r.part0[15] );
tran (\sa_ctrl_rst_dat[27][15] , \sa_ctrl_rst_dat[27].f.spare[10] );
tran (\sa_ctrl_rst_dat[27][16] , \sa_ctrl_rst_dat[27].r.part0[16] );
tran (\sa_ctrl_rst_dat[27][16] , \sa_ctrl_rst_dat[27].f.spare[11] );
tran (\sa_ctrl_rst_dat[27][17] , \sa_ctrl_rst_dat[27].r.part0[17] );
tran (\sa_ctrl_rst_dat[27][17] , \sa_ctrl_rst_dat[27].f.spare[12] );
tran (\sa_ctrl_rst_dat[27][18] , \sa_ctrl_rst_dat[27].r.part0[18] );
tran (\sa_ctrl_rst_dat[27][18] , \sa_ctrl_rst_dat[27].f.spare[13] );
tran (\sa_ctrl_rst_dat[27][19] , \sa_ctrl_rst_dat[27].r.part0[19] );
tran (\sa_ctrl_rst_dat[27][19] , \sa_ctrl_rst_dat[27].f.spare[14] );
tran (\sa_ctrl_rst_dat[27][20] , \sa_ctrl_rst_dat[27].r.part0[20] );
tran (\sa_ctrl_rst_dat[27][20] , \sa_ctrl_rst_dat[27].f.spare[15] );
tran (\sa_ctrl_rst_dat[27][21] , \sa_ctrl_rst_dat[27].r.part0[21] );
tran (\sa_ctrl_rst_dat[27][21] , \sa_ctrl_rst_dat[27].f.spare[16] );
tran (\sa_ctrl_rst_dat[27][22] , \sa_ctrl_rst_dat[27].r.part0[22] );
tran (\sa_ctrl_rst_dat[27][22] , \sa_ctrl_rst_dat[27].f.spare[17] );
tran (\sa_ctrl_rst_dat[27][23] , \sa_ctrl_rst_dat[27].r.part0[23] );
tran (\sa_ctrl_rst_dat[27][23] , \sa_ctrl_rst_dat[27].f.spare[18] );
tran (\sa_ctrl_rst_dat[27][24] , \sa_ctrl_rst_dat[27].r.part0[24] );
tran (\sa_ctrl_rst_dat[27][24] , \sa_ctrl_rst_dat[27].f.spare[19] );
tran (\sa_ctrl_rst_dat[27][25] , \sa_ctrl_rst_dat[27].r.part0[25] );
tran (\sa_ctrl_rst_dat[27][25] , \sa_ctrl_rst_dat[27].f.spare[20] );
tran (\sa_ctrl_rst_dat[27][26] , \sa_ctrl_rst_dat[27].r.part0[26] );
tran (\sa_ctrl_rst_dat[27][26] , \sa_ctrl_rst_dat[27].f.spare[21] );
tran (\sa_ctrl_rst_dat[27][27] , \sa_ctrl_rst_dat[27].r.part0[27] );
tran (\sa_ctrl_rst_dat[27][27] , \sa_ctrl_rst_dat[27].f.spare[22] );
tran (\sa_ctrl_rst_dat[27][28] , \sa_ctrl_rst_dat[27].r.part0[28] );
tran (\sa_ctrl_rst_dat[27][28] , \sa_ctrl_rst_dat[27].f.spare[23] );
tran (\sa_ctrl_rst_dat[27][29] , \sa_ctrl_rst_dat[27].r.part0[29] );
tran (\sa_ctrl_rst_dat[27][29] , \sa_ctrl_rst_dat[27].f.spare[24] );
tran (\sa_ctrl_rst_dat[27][30] , \sa_ctrl_rst_dat[27].r.part0[30] );
tran (\sa_ctrl_rst_dat[27][30] , \sa_ctrl_rst_dat[27].f.spare[25] );
tran (\sa_ctrl_rst_dat[27][31] , \sa_ctrl_rst_dat[27].r.part0[31] );
tran (\sa_ctrl_rst_dat[27][31] , \sa_ctrl_rst_dat[27].f.spare[26] );
tran (\sa_ctrl_rst_dat[28][0] , \sa_ctrl_rst_dat[28].r.part0[0] );
tran (\sa_ctrl_rst_dat[28][0] , \sa_ctrl_rst_dat[28].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[28][1] , \sa_ctrl_rst_dat[28].r.part0[1] );
tran (\sa_ctrl_rst_dat[28][1] , \sa_ctrl_rst_dat[28].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[28][2] , \sa_ctrl_rst_dat[28].r.part0[2] );
tran (\sa_ctrl_rst_dat[28][2] , \sa_ctrl_rst_dat[28].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[28][3] , \sa_ctrl_rst_dat[28].r.part0[3] );
tran (\sa_ctrl_rst_dat[28][3] , \sa_ctrl_rst_dat[28].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[28][4] , \sa_ctrl_rst_dat[28].r.part0[4] );
tran (\sa_ctrl_rst_dat[28][4] , \sa_ctrl_rst_dat[28].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[28][5] , \sa_ctrl_rst_dat[28].r.part0[5] );
tran (\sa_ctrl_rst_dat[28][5] , \sa_ctrl_rst_dat[28].f.spare[0] );
tran (\sa_ctrl_rst_dat[28][6] , \sa_ctrl_rst_dat[28].r.part0[6] );
tran (\sa_ctrl_rst_dat[28][6] , \sa_ctrl_rst_dat[28].f.spare[1] );
tran (\sa_ctrl_rst_dat[28][7] , \sa_ctrl_rst_dat[28].r.part0[7] );
tran (\sa_ctrl_rst_dat[28][7] , \sa_ctrl_rst_dat[28].f.spare[2] );
tran (\sa_ctrl_rst_dat[28][8] , \sa_ctrl_rst_dat[28].r.part0[8] );
tran (\sa_ctrl_rst_dat[28][8] , \sa_ctrl_rst_dat[28].f.spare[3] );
tran (\sa_ctrl_rst_dat[28][9] , \sa_ctrl_rst_dat[28].r.part0[9] );
tran (\sa_ctrl_rst_dat[28][9] , \sa_ctrl_rst_dat[28].f.spare[4] );
tran (\sa_ctrl_rst_dat[28][10] , \sa_ctrl_rst_dat[28].r.part0[10] );
tran (\sa_ctrl_rst_dat[28][10] , \sa_ctrl_rst_dat[28].f.spare[5] );
tran (\sa_ctrl_rst_dat[28][11] , \sa_ctrl_rst_dat[28].r.part0[11] );
tran (\sa_ctrl_rst_dat[28][11] , \sa_ctrl_rst_dat[28].f.spare[6] );
tran (\sa_ctrl_rst_dat[28][12] , \sa_ctrl_rst_dat[28].r.part0[12] );
tran (\sa_ctrl_rst_dat[28][12] , \sa_ctrl_rst_dat[28].f.spare[7] );
tran (\sa_ctrl_rst_dat[28][13] , \sa_ctrl_rst_dat[28].r.part0[13] );
tran (\sa_ctrl_rst_dat[28][13] , \sa_ctrl_rst_dat[28].f.spare[8] );
tran (\sa_ctrl_rst_dat[28][14] , \sa_ctrl_rst_dat[28].r.part0[14] );
tran (\sa_ctrl_rst_dat[28][14] , \sa_ctrl_rst_dat[28].f.spare[9] );
tran (\sa_ctrl_rst_dat[28][15] , \sa_ctrl_rst_dat[28].r.part0[15] );
tran (\sa_ctrl_rst_dat[28][15] , \sa_ctrl_rst_dat[28].f.spare[10] );
tran (\sa_ctrl_rst_dat[28][16] , \sa_ctrl_rst_dat[28].r.part0[16] );
tran (\sa_ctrl_rst_dat[28][16] , \sa_ctrl_rst_dat[28].f.spare[11] );
tran (\sa_ctrl_rst_dat[28][17] , \sa_ctrl_rst_dat[28].r.part0[17] );
tran (\sa_ctrl_rst_dat[28][17] , \sa_ctrl_rst_dat[28].f.spare[12] );
tran (\sa_ctrl_rst_dat[28][18] , \sa_ctrl_rst_dat[28].r.part0[18] );
tran (\sa_ctrl_rst_dat[28][18] , \sa_ctrl_rst_dat[28].f.spare[13] );
tran (\sa_ctrl_rst_dat[28][19] , \sa_ctrl_rst_dat[28].r.part0[19] );
tran (\sa_ctrl_rst_dat[28][19] , \sa_ctrl_rst_dat[28].f.spare[14] );
tran (\sa_ctrl_rst_dat[28][20] , \sa_ctrl_rst_dat[28].r.part0[20] );
tran (\sa_ctrl_rst_dat[28][20] , \sa_ctrl_rst_dat[28].f.spare[15] );
tran (\sa_ctrl_rst_dat[28][21] , \sa_ctrl_rst_dat[28].r.part0[21] );
tran (\sa_ctrl_rst_dat[28][21] , \sa_ctrl_rst_dat[28].f.spare[16] );
tran (\sa_ctrl_rst_dat[28][22] , \sa_ctrl_rst_dat[28].r.part0[22] );
tran (\sa_ctrl_rst_dat[28][22] , \sa_ctrl_rst_dat[28].f.spare[17] );
tran (\sa_ctrl_rst_dat[28][23] , \sa_ctrl_rst_dat[28].r.part0[23] );
tran (\sa_ctrl_rst_dat[28][23] , \sa_ctrl_rst_dat[28].f.spare[18] );
tran (\sa_ctrl_rst_dat[28][24] , \sa_ctrl_rst_dat[28].r.part0[24] );
tran (\sa_ctrl_rst_dat[28][24] , \sa_ctrl_rst_dat[28].f.spare[19] );
tran (\sa_ctrl_rst_dat[28][25] , \sa_ctrl_rst_dat[28].r.part0[25] );
tran (\sa_ctrl_rst_dat[28][25] , \sa_ctrl_rst_dat[28].f.spare[20] );
tran (\sa_ctrl_rst_dat[28][26] , \sa_ctrl_rst_dat[28].r.part0[26] );
tran (\sa_ctrl_rst_dat[28][26] , \sa_ctrl_rst_dat[28].f.spare[21] );
tran (\sa_ctrl_rst_dat[28][27] , \sa_ctrl_rst_dat[28].r.part0[27] );
tran (\sa_ctrl_rst_dat[28][27] , \sa_ctrl_rst_dat[28].f.spare[22] );
tran (\sa_ctrl_rst_dat[28][28] , \sa_ctrl_rst_dat[28].r.part0[28] );
tran (\sa_ctrl_rst_dat[28][28] , \sa_ctrl_rst_dat[28].f.spare[23] );
tran (\sa_ctrl_rst_dat[28][29] , \sa_ctrl_rst_dat[28].r.part0[29] );
tran (\sa_ctrl_rst_dat[28][29] , \sa_ctrl_rst_dat[28].f.spare[24] );
tran (\sa_ctrl_rst_dat[28][30] , \sa_ctrl_rst_dat[28].r.part0[30] );
tran (\sa_ctrl_rst_dat[28][30] , \sa_ctrl_rst_dat[28].f.spare[25] );
tran (\sa_ctrl_rst_dat[28][31] , \sa_ctrl_rst_dat[28].r.part0[31] );
tran (\sa_ctrl_rst_dat[28][31] , \sa_ctrl_rst_dat[28].f.spare[26] );
tran (\sa_ctrl_rst_dat[29][0] , \sa_ctrl_rst_dat[29].r.part0[0] );
tran (\sa_ctrl_rst_dat[29][0] , \sa_ctrl_rst_dat[29].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[29][1] , \sa_ctrl_rst_dat[29].r.part0[1] );
tran (\sa_ctrl_rst_dat[29][1] , \sa_ctrl_rst_dat[29].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[29][2] , \sa_ctrl_rst_dat[29].r.part0[2] );
tran (\sa_ctrl_rst_dat[29][2] , \sa_ctrl_rst_dat[29].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[29][3] , \sa_ctrl_rst_dat[29].r.part0[3] );
tran (\sa_ctrl_rst_dat[29][3] , \sa_ctrl_rst_dat[29].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[29][4] , \sa_ctrl_rst_dat[29].r.part0[4] );
tran (\sa_ctrl_rst_dat[29][4] , \sa_ctrl_rst_dat[29].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[29][5] , \sa_ctrl_rst_dat[29].r.part0[5] );
tran (\sa_ctrl_rst_dat[29][5] , \sa_ctrl_rst_dat[29].f.spare[0] );
tran (\sa_ctrl_rst_dat[29][6] , \sa_ctrl_rst_dat[29].r.part0[6] );
tran (\sa_ctrl_rst_dat[29][6] , \sa_ctrl_rst_dat[29].f.spare[1] );
tran (\sa_ctrl_rst_dat[29][7] , \sa_ctrl_rst_dat[29].r.part0[7] );
tran (\sa_ctrl_rst_dat[29][7] , \sa_ctrl_rst_dat[29].f.spare[2] );
tran (\sa_ctrl_rst_dat[29][8] , \sa_ctrl_rst_dat[29].r.part0[8] );
tran (\sa_ctrl_rst_dat[29][8] , \sa_ctrl_rst_dat[29].f.spare[3] );
tran (\sa_ctrl_rst_dat[29][9] , \sa_ctrl_rst_dat[29].r.part0[9] );
tran (\sa_ctrl_rst_dat[29][9] , \sa_ctrl_rst_dat[29].f.spare[4] );
tran (\sa_ctrl_rst_dat[29][10] , \sa_ctrl_rst_dat[29].r.part0[10] );
tran (\sa_ctrl_rst_dat[29][10] , \sa_ctrl_rst_dat[29].f.spare[5] );
tran (\sa_ctrl_rst_dat[29][11] , \sa_ctrl_rst_dat[29].r.part0[11] );
tran (\sa_ctrl_rst_dat[29][11] , \sa_ctrl_rst_dat[29].f.spare[6] );
tran (\sa_ctrl_rst_dat[29][12] , \sa_ctrl_rst_dat[29].r.part0[12] );
tran (\sa_ctrl_rst_dat[29][12] , \sa_ctrl_rst_dat[29].f.spare[7] );
tran (\sa_ctrl_rst_dat[29][13] , \sa_ctrl_rst_dat[29].r.part0[13] );
tran (\sa_ctrl_rst_dat[29][13] , \sa_ctrl_rst_dat[29].f.spare[8] );
tran (\sa_ctrl_rst_dat[29][14] , \sa_ctrl_rst_dat[29].r.part0[14] );
tran (\sa_ctrl_rst_dat[29][14] , \sa_ctrl_rst_dat[29].f.spare[9] );
tran (\sa_ctrl_rst_dat[29][15] , \sa_ctrl_rst_dat[29].r.part0[15] );
tran (\sa_ctrl_rst_dat[29][15] , \sa_ctrl_rst_dat[29].f.spare[10] );
tran (\sa_ctrl_rst_dat[29][16] , \sa_ctrl_rst_dat[29].r.part0[16] );
tran (\sa_ctrl_rst_dat[29][16] , \sa_ctrl_rst_dat[29].f.spare[11] );
tran (\sa_ctrl_rst_dat[29][17] , \sa_ctrl_rst_dat[29].r.part0[17] );
tran (\sa_ctrl_rst_dat[29][17] , \sa_ctrl_rst_dat[29].f.spare[12] );
tran (\sa_ctrl_rst_dat[29][18] , \sa_ctrl_rst_dat[29].r.part0[18] );
tran (\sa_ctrl_rst_dat[29][18] , \sa_ctrl_rst_dat[29].f.spare[13] );
tran (\sa_ctrl_rst_dat[29][19] , \sa_ctrl_rst_dat[29].r.part0[19] );
tran (\sa_ctrl_rst_dat[29][19] , \sa_ctrl_rst_dat[29].f.spare[14] );
tran (\sa_ctrl_rst_dat[29][20] , \sa_ctrl_rst_dat[29].r.part0[20] );
tran (\sa_ctrl_rst_dat[29][20] , \sa_ctrl_rst_dat[29].f.spare[15] );
tran (\sa_ctrl_rst_dat[29][21] , \sa_ctrl_rst_dat[29].r.part0[21] );
tran (\sa_ctrl_rst_dat[29][21] , \sa_ctrl_rst_dat[29].f.spare[16] );
tran (\sa_ctrl_rst_dat[29][22] , \sa_ctrl_rst_dat[29].r.part0[22] );
tran (\sa_ctrl_rst_dat[29][22] , \sa_ctrl_rst_dat[29].f.spare[17] );
tran (\sa_ctrl_rst_dat[29][23] , \sa_ctrl_rst_dat[29].r.part0[23] );
tran (\sa_ctrl_rst_dat[29][23] , \sa_ctrl_rst_dat[29].f.spare[18] );
tran (\sa_ctrl_rst_dat[29][24] , \sa_ctrl_rst_dat[29].r.part0[24] );
tran (\sa_ctrl_rst_dat[29][24] , \sa_ctrl_rst_dat[29].f.spare[19] );
tran (\sa_ctrl_rst_dat[29][25] , \sa_ctrl_rst_dat[29].r.part0[25] );
tran (\sa_ctrl_rst_dat[29][25] , \sa_ctrl_rst_dat[29].f.spare[20] );
tran (\sa_ctrl_rst_dat[29][26] , \sa_ctrl_rst_dat[29].r.part0[26] );
tran (\sa_ctrl_rst_dat[29][26] , \sa_ctrl_rst_dat[29].f.spare[21] );
tran (\sa_ctrl_rst_dat[29][27] , \sa_ctrl_rst_dat[29].r.part0[27] );
tran (\sa_ctrl_rst_dat[29][27] , \sa_ctrl_rst_dat[29].f.spare[22] );
tran (\sa_ctrl_rst_dat[29][28] , \sa_ctrl_rst_dat[29].r.part0[28] );
tran (\sa_ctrl_rst_dat[29][28] , \sa_ctrl_rst_dat[29].f.spare[23] );
tran (\sa_ctrl_rst_dat[29][29] , \sa_ctrl_rst_dat[29].r.part0[29] );
tran (\sa_ctrl_rst_dat[29][29] , \sa_ctrl_rst_dat[29].f.spare[24] );
tran (\sa_ctrl_rst_dat[29][30] , \sa_ctrl_rst_dat[29].r.part0[30] );
tran (\sa_ctrl_rst_dat[29][30] , \sa_ctrl_rst_dat[29].f.spare[25] );
tran (\sa_ctrl_rst_dat[29][31] , \sa_ctrl_rst_dat[29].r.part0[31] );
tran (\sa_ctrl_rst_dat[29][31] , \sa_ctrl_rst_dat[29].f.spare[26] );
tran (\sa_ctrl_rst_dat[30][0] , \sa_ctrl_rst_dat[30].r.part0[0] );
tran (\sa_ctrl_rst_dat[30][0] , \sa_ctrl_rst_dat[30].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[30][1] , \sa_ctrl_rst_dat[30].r.part0[1] );
tran (\sa_ctrl_rst_dat[30][1] , \sa_ctrl_rst_dat[30].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[30][2] , \sa_ctrl_rst_dat[30].r.part0[2] );
tran (\sa_ctrl_rst_dat[30][2] , \sa_ctrl_rst_dat[30].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[30][3] , \sa_ctrl_rst_dat[30].r.part0[3] );
tran (\sa_ctrl_rst_dat[30][3] , \sa_ctrl_rst_dat[30].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[30][4] , \sa_ctrl_rst_dat[30].r.part0[4] );
tran (\sa_ctrl_rst_dat[30][4] , \sa_ctrl_rst_dat[30].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[30][5] , \sa_ctrl_rst_dat[30].r.part0[5] );
tran (\sa_ctrl_rst_dat[30][5] , \sa_ctrl_rst_dat[30].f.spare[0] );
tran (\sa_ctrl_rst_dat[30][6] , \sa_ctrl_rst_dat[30].r.part0[6] );
tran (\sa_ctrl_rst_dat[30][6] , \sa_ctrl_rst_dat[30].f.spare[1] );
tran (\sa_ctrl_rst_dat[30][7] , \sa_ctrl_rst_dat[30].r.part0[7] );
tran (\sa_ctrl_rst_dat[30][7] , \sa_ctrl_rst_dat[30].f.spare[2] );
tran (\sa_ctrl_rst_dat[30][8] , \sa_ctrl_rst_dat[30].r.part0[8] );
tran (\sa_ctrl_rst_dat[30][8] , \sa_ctrl_rst_dat[30].f.spare[3] );
tran (\sa_ctrl_rst_dat[30][9] , \sa_ctrl_rst_dat[30].r.part0[9] );
tran (\sa_ctrl_rst_dat[30][9] , \sa_ctrl_rst_dat[30].f.spare[4] );
tran (\sa_ctrl_rst_dat[30][10] , \sa_ctrl_rst_dat[30].r.part0[10] );
tran (\sa_ctrl_rst_dat[30][10] , \sa_ctrl_rst_dat[30].f.spare[5] );
tran (\sa_ctrl_rst_dat[30][11] , \sa_ctrl_rst_dat[30].r.part0[11] );
tran (\sa_ctrl_rst_dat[30][11] , \sa_ctrl_rst_dat[30].f.spare[6] );
tran (\sa_ctrl_rst_dat[30][12] , \sa_ctrl_rst_dat[30].r.part0[12] );
tran (\sa_ctrl_rst_dat[30][12] , \sa_ctrl_rst_dat[30].f.spare[7] );
tran (\sa_ctrl_rst_dat[30][13] , \sa_ctrl_rst_dat[30].r.part0[13] );
tran (\sa_ctrl_rst_dat[30][13] , \sa_ctrl_rst_dat[30].f.spare[8] );
tran (\sa_ctrl_rst_dat[30][14] , \sa_ctrl_rst_dat[30].r.part0[14] );
tran (\sa_ctrl_rst_dat[30][14] , \sa_ctrl_rst_dat[30].f.spare[9] );
tran (\sa_ctrl_rst_dat[30][15] , \sa_ctrl_rst_dat[30].r.part0[15] );
tran (\sa_ctrl_rst_dat[30][15] , \sa_ctrl_rst_dat[30].f.spare[10] );
tran (\sa_ctrl_rst_dat[30][16] , \sa_ctrl_rst_dat[30].r.part0[16] );
tran (\sa_ctrl_rst_dat[30][16] , \sa_ctrl_rst_dat[30].f.spare[11] );
tran (\sa_ctrl_rst_dat[30][17] , \sa_ctrl_rst_dat[30].r.part0[17] );
tran (\sa_ctrl_rst_dat[30][17] , \sa_ctrl_rst_dat[30].f.spare[12] );
tran (\sa_ctrl_rst_dat[30][18] , \sa_ctrl_rst_dat[30].r.part0[18] );
tran (\sa_ctrl_rst_dat[30][18] , \sa_ctrl_rst_dat[30].f.spare[13] );
tran (\sa_ctrl_rst_dat[30][19] , \sa_ctrl_rst_dat[30].r.part0[19] );
tran (\sa_ctrl_rst_dat[30][19] , \sa_ctrl_rst_dat[30].f.spare[14] );
tran (\sa_ctrl_rst_dat[30][20] , \sa_ctrl_rst_dat[30].r.part0[20] );
tran (\sa_ctrl_rst_dat[30][20] , \sa_ctrl_rst_dat[30].f.spare[15] );
tran (\sa_ctrl_rst_dat[30][21] , \sa_ctrl_rst_dat[30].r.part0[21] );
tran (\sa_ctrl_rst_dat[30][21] , \sa_ctrl_rst_dat[30].f.spare[16] );
tran (\sa_ctrl_rst_dat[30][22] , \sa_ctrl_rst_dat[30].r.part0[22] );
tran (\sa_ctrl_rst_dat[30][22] , \sa_ctrl_rst_dat[30].f.spare[17] );
tran (\sa_ctrl_rst_dat[30][23] , \sa_ctrl_rst_dat[30].r.part0[23] );
tran (\sa_ctrl_rst_dat[30][23] , \sa_ctrl_rst_dat[30].f.spare[18] );
tran (\sa_ctrl_rst_dat[30][24] , \sa_ctrl_rst_dat[30].r.part0[24] );
tran (\sa_ctrl_rst_dat[30][24] , \sa_ctrl_rst_dat[30].f.spare[19] );
tran (\sa_ctrl_rst_dat[30][25] , \sa_ctrl_rst_dat[30].r.part0[25] );
tran (\sa_ctrl_rst_dat[30][25] , \sa_ctrl_rst_dat[30].f.spare[20] );
tran (\sa_ctrl_rst_dat[30][26] , \sa_ctrl_rst_dat[30].r.part0[26] );
tran (\sa_ctrl_rst_dat[30][26] , \sa_ctrl_rst_dat[30].f.spare[21] );
tran (\sa_ctrl_rst_dat[30][27] , \sa_ctrl_rst_dat[30].r.part0[27] );
tran (\sa_ctrl_rst_dat[30][27] , \sa_ctrl_rst_dat[30].f.spare[22] );
tran (\sa_ctrl_rst_dat[30][28] , \sa_ctrl_rst_dat[30].r.part0[28] );
tran (\sa_ctrl_rst_dat[30][28] , \sa_ctrl_rst_dat[30].f.spare[23] );
tran (\sa_ctrl_rst_dat[30][29] , \sa_ctrl_rst_dat[30].r.part0[29] );
tran (\sa_ctrl_rst_dat[30][29] , \sa_ctrl_rst_dat[30].f.spare[24] );
tran (\sa_ctrl_rst_dat[30][30] , \sa_ctrl_rst_dat[30].r.part0[30] );
tran (\sa_ctrl_rst_dat[30][30] , \sa_ctrl_rst_dat[30].f.spare[25] );
tran (\sa_ctrl_rst_dat[30][31] , \sa_ctrl_rst_dat[30].r.part0[31] );
tran (\sa_ctrl_rst_dat[30][31] , \sa_ctrl_rst_dat[30].f.spare[26] );
tran (\sa_ctrl_rst_dat[31][0] , \sa_ctrl_rst_dat[31].r.part0[0] );
tran (\sa_ctrl_rst_dat[31][0] , \sa_ctrl_rst_dat[31].f.sa_event_sel[0] );
tran (\sa_ctrl_rst_dat[31][1] , \sa_ctrl_rst_dat[31].r.part0[1] );
tran (\sa_ctrl_rst_dat[31][1] , \sa_ctrl_rst_dat[31].f.sa_event_sel[1] );
tran (\sa_ctrl_rst_dat[31][2] , \sa_ctrl_rst_dat[31].r.part0[2] );
tran (\sa_ctrl_rst_dat[31][2] , \sa_ctrl_rst_dat[31].f.sa_event_sel[2] );
tran (\sa_ctrl_rst_dat[31][3] , \sa_ctrl_rst_dat[31].r.part0[3] );
tran (\sa_ctrl_rst_dat[31][3] , \sa_ctrl_rst_dat[31].f.sa_event_sel[3] );
tran (\sa_ctrl_rst_dat[31][4] , \sa_ctrl_rst_dat[31].r.part0[4] );
tran (\sa_ctrl_rst_dat[31][4] , \sa_ctrl_rst_dat[31].f.sa_event_sel[4] );
tran (\sa_ctrl_rst_dat[31][5] , \sa_ctrl_rst_dat[31].r.part0[5] );
tran (\sa_ctrl_rst_dat[31][5] , \sa_ctrl_rst_dat[31].f.spare[0] );
tran (\sa_ctrl_rst_dat[31][6] , \sa_ctrl_rst_dat[31].r.part0[6] );
tran (\sa_ctrl_rst_dat[31][6] , \sa_ctrl_rst_dat[31].f.spare[1] );
tran (\sa_ctrl_rst_dat[31][7] , \sa_ctrl_rst_dat[31].r.part0[7] );
tran (\sa_ctrl_rst_dat[31][7] , \sa_ctrl_rst_dat[31].f.spare[2] );
tran (\sa_ctrl_rst_dat[31][8] , \sa_ctrl_rst_dat[31].r.part0[8] );
tran (\sa_ctrl_rst_dat[31][8] , \sa_ctrl_rst_dat[31].f.spare[3] );
tran (\sa_ctrl_rst_dat[31][9] , \sa_ctrl_rst_dat[31].r.part0[9] );
tran (\sa_ctrl_rst_dat[31][9] , \sa_ctrl_rst_dat[31].f.spare[4] );
tran (\sa_ctrl_rst_dat[31][10] , \sa_ctrl_rst_dat[31].r.part0[10] );
tran (\sa_ctrl_rst_dat[31][10] , \sa_ctrl_rst_dat[31].f.spare[5] );
tran (\sa_ctrl_rst_dat[31][11] , \sa_ctrl_rst_dat[31].r.part0[11] );
tran (\sa_ctrl_rst_dat[31][11] , \sa_ctrl_rst_dat[31].f.spare[6] );
tran (\sa_ctrl_rst_dat[31][12] , \sa_ctrl_rst_dat[31].r.part0[12] );
tran (\sa_ctrl_rst_dat[31][12] , \sa_ctrl_rst_dat[31].f.spare[7] );
tran (\sa_ctrl_rst_dat[31][13] , \sa_ctrl_rst_dat[31].r.part0[13] );
tran (\sa_ctrl_rst_dat[31][13] , \sa_ctrl_rst_dat[31].f.spare[8] );
tran (\sa_ctrl_rst_dat[31][14] , \sa_ctrl_rst_dat[31].r.part0[14] );
tran (\sa_ctrl_rst_dat[31][14] , \sa_ctrl_rst_dat[31].f.spare[9] );
tran (\sa_ctrl_rst_dat[31][15] , \sa_ctrl_rst_dat[31].r.part0[15] );
tran (\sa_ctrl_rst_dat[31][15] , \sa_ctrl_rst_dat[31].f.spare[10] );
tran (\sa_ctrl_rst_dat[31][16] , \sa_ctrl_rst_dat[31].r.part0[16] );
tran (\sa_ctrl_rst_dat[31][16] , \sa_ctrl_rst_dat[31].f.spare[11] );
tran (\sa_ctrl_rst_dat[31][17] , \sa_ctrl_rst_dat[31].r.part0[17] );
tran (\sa_ctrl_rst_dat[31][17] , \sa_ctrl_rst_dat[31].f.spare[12] );
tran (\sa_ctrl_rst_dat[31][18] , \sa_ctrl_rst_dat[31].r.part0[18] );
tran (\sa_ctrl_rst_dat[31][18] , \sa_ctrl_rst_dat[31].f.spare[13] );
tran (\sa_ctrl_rst_dat[31][19] , \sa_ctrl_rst_dat[31].r.part0[19] );
tran (\sa_ctrl_rst_dat[31][19] , \sa_ctrl_rst_dat[31].f.spare[14] );
tran (\sa_ctrl_rst_dat[31][20] , \sa_ctrl_rst_dat[31].r.part0[20] );
tran (\sa_ctrl_rst_dat[31][20] , \sa_ctrl_rst_dat[31].f.spare[15] );
tran (\sa_ctrl_rst_dat[31][21] , \sa_ctrl_rst_dat[31].r.part0[21] );
tran (\sa_ctrl_rst_dat[31][21] , \sa_ctrl_rst_dat[31].f.spare[16] );
tran (\sa_ctrl_rst_dat[31][22] , \sa_ctrl_rst_dat[31].r.part0[22] );
tran (\sa_ctrl_rst_dat[31][22] , \sa_ctrl_rst_dat[31].f.spare[17] );
tran (\sa_ctrl_rst_dat[31][23] , \sa_ctrl_rst_dat[31].r.part0[23] );
tran (\sa_ctrl_rst_dat[31][23] , \sa_ctrl_rst_dat[31].f.spare[18] );
tran (\sa_ctrl_rst_dat[31][24] , \sa_ctrl_rst_dat[31].r.part0[24] );
tran (\sa_ctrl_rst_dat[31][24] , \sa_ctrl_rst_dat[31].f.spare[19] );
tran (\sa_ctrl_rst_dat[31][25] , \sa_ctrl_rst_dat[31].r.part0[25] );
tran (\sa_ctrl_rst_dat[31][25] , \sa_ctrl_rst_dat[31].f.spare[20] );
tran (\sa_ctrl_rst_dat[31][26] , \sa_ctrl_rst_dat[31].r.part0[26] );
tran (\sa_ctrl_rst_dat[31][26] , \sa_ctrl_rst_dat[31].f.spare[21] );
tran (\sa_ctrl_rst_dat[31][27] , \sa_ctrl_rst_dat[31].r.part0[27] );
tran (\sa_ctrl_rst_dat[31][27] , \sa_ctrl_rst_dat[31].f.spare[22] );
tran (\sa_ctrl_rst_dat[31][28] , \sa_ctrl_rst_dat[31].r.part0[28] );
tran (\sa_ctrl_rst_dat[31][28] , \sa_ctrl_rst_dat[31].f.spare[23] );
tran (\sa_ctrl_rst_dat[31][29] , \sa_ctrl_rst_dat[31].r.part0[29] );
tran (\sa_ctrl_rst_dat[31][29] , \sa_ctrl_rst_dat[31].f.spare[24] );
tran (\sa_ctrl_rst_dat[31][30] , \sa_ctrl_rst_dat[31].r.part0[30] );
tran (\sa_ctrl_rst_dat[31][30] , \sa_ctrl_rst_dat[31].f.spare[25] );
tran (\sa_ctrl_rst_dat[31][31] , \sa_ctrl_rst_dat[31].r.part0[31] );
tran (\sa_ctrl_rst_dat[31][31] , \sa_ctrl_rst_dat[31].f.spare[26] );
Q_BUF U0 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][31] ));
Q_BUF U1 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][30] ));
Q_BUF U2 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][29] ));
Q_BUF U3 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][28] ));
Q_BUF U4 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][27] ));
Q_BUF U5 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][26] ));
Q_BUF U6 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][25] ));
Q_BUF U7 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][24] ));
Q_BUF U8 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][23] ));
Q_BUF U9 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][22] ));
Q_BUF U10 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][21] ));
Q_BUF U11 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][20] ));
Q_BUF U12 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][19] ));
Q_BUF U13 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][18] ));
Q_BUF U14 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][17] ));
Q_BUF U15 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][16] ));
Q_BUF U16 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][15] ));
Q_BUF U17 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][14] ));
Q_BUF U18 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][13] ));
Q_BUF U19 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][12] ));
Q_BUF U20 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][11] ));
Q_BUF U21 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][10] ));
Q_BUF U22 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][9] ));
Q_BUF U23 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][8] ));
Q_BUF U24 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][7] ));
Q_BUF U25 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][6] ));
Q_BUF U26 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][5] ));
Q_BUF U27 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][4] ));
Q_BUF U28 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][3] ));
Q_BUF U29 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][2] ));
Q_BUF U30 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][1] ));
Q_BUF U31 ( .A(n2), .Z(\sa_ctrl_rst_dat[31][0] ));
Q_BUF U32 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][31] ));
Q_BUF U33 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][30] ));
Q_BUF U34 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][29] ));
Q_BUF U35 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][28] ));
Q_BUF U36 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][27] ));
Q_BUF U37 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][26] ));
Q_BUF U38 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][25] ));
Q_BUF U39 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][24] ));
Q_BUF U40 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][23] ));
Q_BUF U41 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][22] ));
Q_BUF U42 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][21] ));
Q_BUF U43 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][20] ));
Q_BUF U44 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][19] ));
Q_BUF U45 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][18] ));
Q_BUF U46 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][17] ));
Q_BUF U47 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][16] ));
Q_BUF U48 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][15] ));
Q_BUF U49 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][14] ));
Q_BUF U50 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][13] ));
Q_BUF U51 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][12] ));
Q_BUF U52 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][11] ));
Q_BUF U53 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][10] ));
Q_BUF U54 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][9] ));
Q_BUF U55 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][8] ));
Q_BUF U56 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][7] ));
Q_BUF U57 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][6] ));
Q_BUF U58 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][5] ));
Q_BUF U59 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][4] ));
Q_BUF U60 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][3] ));
Q_BUF U61 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][2] ));
Q_BUF U62 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][1] ));
Q_BUF U63 ( .A(n2), .Z(\sa_ctrl_rst_dat[30][0] ));
Q_BUF U64 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][31] ));
Q_BUF U65 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][30] ));
Q_BUF U66 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][29] ));
Q_BUF U67 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][28] ));
Q_BUF U68 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][27] ));
Q_BUF U69 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][26] ));
Q_BUF U70 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][25] ));
Q_BUF U71 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][24] ));
Q_BUF U72 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][23] ));
Q_BUF U73 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][22] ));
Q_BUF U74 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][21] ));
Q_BUF U75 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][20] ));
Q_BUF U76 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][19] ));
Q_BUF U77 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][18] ));
Q_BUF U78 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][17] ));
Q_BUF U79 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][16] ));
Q_BUF U80 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][15] ));
Q_BUF U81 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][14] ));
Q_BUF U82 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][13] ));
Q_BUF U83 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][12] ));
Q_BUF U84 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][11] ));
Q_BUF U85 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][10] ));
Q_BUF U86 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][9] ));
Q_BUF U87 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][8] ));
Q_BUF U88 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][7] ));
Q_BUF U89 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][6] ));
Q_BUF U90 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][5] ));
Q_BUF U91 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][4] ));
Q_BUF U92 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][3] ));
Q_BUF U93 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][2] ));
Q_BUF U94 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][1] ));
Q_BUF U95 ( .A(n2), .Z(\sa_ctrl_rst_dat[29][0] ));
Q_BUF U96 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][31] ));
Q_BUF U97 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][30] ));
Q_BUF U98 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][29] ));
Q_BUF U99 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][28] ));
Q_BUF U100 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][27] ));
Q_BUF U101 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][26] ));
Q_BUF U102 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][25] ));
Q_BUF U103 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][24] ));
Q_BUF U104 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][23] ));
Q_BUF U105 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][22] ));
Q_BUF U106 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][21] ));
Q_BUF U107 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][20] ));
Q_BUF U108 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][19] ));
Q_BUF U109 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][18] ));
Q_BUF U110 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][17] ));
Q_BUF U111 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][16] ));
Q_BUF U112 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][15] ));
Q_BUF U113 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][14] ));
Q_BUF U114 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][13] ));
Q_BUF U115 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][12] ));
Q_BUF U116 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][11] ));
Q_BUF U117 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][10] ));
Q_BUF U118 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][9] ));
Q_BUF U119 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][8] ));
Q_BUF U120 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][7] ));
Q_BUF U121 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][6] ));
Q_BUF U122 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][5] ));
Q_BUF U123 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][4] ));
Q_BUF U124 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][3] ));
Q_BUF U125 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][2] ));
Q_BUF U126 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][1] ));
Q_BUF U127 ( .A(n2), .Z(\sa_ctrl_rst_dat[28][0] ));
Q_BUF U128 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][31] ));
Q_BUF U129 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][30] ));
Q_BUF U130 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][29] ));
Q_BUF U131 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][28] ));
Q_BUF U132 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][27] ));
Q_BUF U133 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][26] ));
Q_BUF U134 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][25] ));
Q_BUF U135 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][24] ));
Q_BUF U136 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][23] ));
Q_BUF U137 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][22] ));
Q_BUF U138 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][21] ));
Q_BUF U139 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][20] ));
Q_BUF U140 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][19] ));
Q_BUF U141 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][18] ));
Q_BUF U142 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][17] ));
Q_BUF U143 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][16] ));
Q_BUF U144 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][15] ));
Q_BUF U145 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][14] ));
Q_BUF U146 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][13] ));
Q_BUF U147 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][12] ));
Q_BUF U148 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][11] ));
Q_BUF U149 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][10] ));
Q_BUF U150 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][9] ));
Q_BUF U151 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][8] ));
Q_BUF U152 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][7] ));
Q_BUF U153 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][6] ));
Q_BUF U154 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][5] ));
Q_BUF U155 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][4] ));
Q_BUF U156 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][3] ));
Q_BUF U157 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][2] ));
Q_BUF U158 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][1] ));
Q_BUF U159 ( .A(n2), .Z(\sa_ctrl_rst_dat[27][0] ));
Q_BUF U160 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][31] ));
Q_BUF U161 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][30] ));
Q_BUF U162 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][29] ));
Q_BUF U163 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][28] ));
Q_BUF U164 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][27] ));
Q_BUF U165 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][26] ));
Q_BUF U166 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][25] ));
Q_BUF U167 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][24] ));
Q_BUF U168 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][23] ));
Q_BUF U169 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][22] ));
Q_BUF U170 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][21] ));
Q_BUF U171 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][20] ));
Q_BUF U172 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][19] ));
Q_BUF U173 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][18] ));
Q_BUF U174 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][17] ));
Q_BUF U175 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][16] ));
Q_BUF U176 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][15] ));
Q_BUF U177 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][14] ));
Q_BUF U178 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][13] ));
Q_BUF U179 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][12] ));
Q_BUF U180 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][11] ));
Q_BUF U181 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][10] ));
Q_BUF U182 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][9] ));
Q_BUF U183 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][8] ));
Q_BUF U184 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][7] ));
Q_BUF U185 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][6] ));
Q_BUF U186 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][5] ));
Q_BUF U187 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][4] ));
Q_BUF U188 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][3] ));
Q_BUF U189 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][2] ));
Q_BUF U190 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][1] ));
Q_BUF U191 ( .A(n2), .Z(\sa_ctrl_rst_dat[26][0] ));
Q_BUF U192 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][31] ));
Q_BUF U193 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][30] ));
Q_BUF U194 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][29] ));
Q_BUF U195 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][28] ));
Q_BUF U196 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][27] ));
Q_BUF U197 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][26] ));
Q_BUF U198 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][25] ));
Q_BUF U199 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][24] ));
Q_BUF U200 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][23] ));
Q_BUF U201 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][22] ));
Q_BUF U202 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][21] ));
Q_BUF U203 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][20] ));
Q_BUF U204 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][19] ));
Q_BUF U205 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][18] ));
Q_BUF U206 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][17] ));
Q_BUF U207 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][16] ));
Q_BUF U208 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][15] ));
Q_BUF U209 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][14] ));
Q_BUF U210 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][13] ));
Q_BUF U211 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][12] ));
Q_BUF U212 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][11] ));
Q_BUF U213 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][10] ));
Q_BUF U214 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][9] ));
Q_BUF U215 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][8] ));
Q_BUF U216 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][7] ));
Q_BUF U217 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][6] ));
Q_BUF U218 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][5] ));
Q_BUF U219 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][4] ));
Q_BUF U220 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][3] ));
Q_BUF U221 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][2] ));
Q_BUF U222 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][1] ));
Q_BUF U223 ( .A(n2), .Z(\sa_ctrl_rst_dat[25][0] ));
Q_BUF U224 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][31] ));
Q_BUF U225 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][30] ));
Q_BUF U226 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][29] ));
Q_BUF U227 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][28] ));
Q_BUF U228 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][27] ));
Q_BUF U229 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][26] ));
Q_BUF U230 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][25] ));
Q_BUF U231 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][24] ));
Q_BUF U232 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][23] ));
Q_BUF U233 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][22] ));
Q_BUF U234 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][21] ));
Q_BUF U235 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][20] ));
Q_BUF U236 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][19] ));
Q_BUF U237 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][18] ));
Q_BUF U238 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][17] ));
Q_BUF U239 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][16] ));
Q_BUF U240 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][15] ));
Q_BUF U241 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][14] ));
Q_BUF U242 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][13] ));
Q_BUF U243 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][12] ));
Q_BUF U244 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][11] ));
Q_BUF U245 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][10] ));
Q_BUF U246 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][9] ));
Q_BUF U247 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][8] ));
Q_BUF U248 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][7] ));
Q_BUF U249 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][6] ));
Q_BUF U250 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][5] ));
Q_BUF U251 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][4] ));
Q_BUF U252 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][3] ));
Q_BUF U253 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][2] ));
Q_BUF U254 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][1] ));
Q_BUF U255 ( .A(n2), .Z(\sa_ctrl_rst_dat[24][0] ));
Q_BUF U256 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][31] ));
Q_BUF U257 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][30] ));
Q_BUF U258 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][29] ));
Q_BUF U259 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][28] ));
Q_BUF U260 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][27] ));
Q_BUF U261 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][26] ));
Q_BUF U262 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][25] ));
Q_BUF U263 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][24] ));
Q_BUF U264 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][23] ));
Q_BUF U265 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][22] ));
Q_BUF U266 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][21] ));
Q_BUF U267 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][20] ));
Q_BUF U268 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][19] ));
Q_BUF U269 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][18] ));
Q_BUF U270 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][17] ));
Q_BUF U271 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][16] ));
Q_BUF U272 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][15] ));
Q_BUF U273 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][14] ));
Q_BUF U274 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][13] ));
Q_BUF U275 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][12] ));
Q_BUF U276 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][11] ));
Q_BUF U277 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][10] ));
Q_BUF U278 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][9] ));
Q_BUF U279 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][8] ));
Q_BUF U280 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][7] ));
Q_BUF U281 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][6] ));
Q_BUF U282 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][5] ));
Q_BUF U283 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][4] ));
Q_BUF U284 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][3] ));
Q_BUF U285 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][2] ));
Q_BUF U286 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][1] ));
Q_BUF U287 ( .A(n2), .Z(\sa_ctrl_rst_dat[23][0] ));
Q_BUF U288 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][31] ));
Q_BUF U289 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][30] ));
Q_BUF U290 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][29] ));
Q_BUF U291 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][28] ));
Q_BUF U292 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][27] ));
Q_BUF U293 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][26] ));
Q_BUF U294 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][25] ));
Q_BUF U295 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][24] ));
Q_BUF U296 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][23] ));
Q_BUF U297 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][22] ));
Q_BUF U298 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][21] ));
Q_BUF U299 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][20] ));
Q_BUF U300 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][19] ));
Q_BUF U301 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][18] ));
Q_BUF U302 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][17] ));
Q_BUF U303 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][16] ));
Q_BUF U304 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][15] ));
Q_BUF U305 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][14] ));
Q_BUF U306 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][13] ));
Q_BUF U307 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][12] ));
Q_BUF U308 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][11] ));
Q_BUF U309 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][10] ));
Q_BUF U310 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][9] ));
Q_BUF U311 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][8] ));
Q_BUF U312 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][7] ));
Q_BUF U313 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][6] ));
Q_BUF U314 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][5] ));
Q_BUF U315 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][4] ));
Q_BUF U316 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][3] ));
Q_BUF U317 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][2] ));
Q_BUF U318 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][1] ));
Q_BUF U319 ( .A(n2), .Z(\sa_ctrl_rst_dat[22][0] ));
Q_BUF U320 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][31] ));
Q_BUF U321 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][30] ));
Q_BUF U322 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][29] ));
Q_BUF U323 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][28] ));
Q_BUF U324 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][27] ));
Q_BUF U325 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][26] ));
Q_BUF U326 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][25] ));
Q_BUF U327 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][24] ));
Q_BUF U328 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][23] ));
Q_BUF U329 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][22] ));
Q_BUF U330 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][21] ));
Q_BUF U331 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][20] ));
Q_BUF U332 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][19] ));
Q_BUF U333 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][18] ));
Q_BUF U334 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][17] ));
Q_BUF U335 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][16] ));
Q_BUF U336 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][15] ));
Q_BUF U337 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][14] ));
Q_BUF U338 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][13] ));
Q_BUF U339 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][12] ));
Q_BUF U340 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][11] ));
Q_BUF U341 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][10] ));
Q_BUF U342 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][9] ));
Q_BUF U343 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][8] ));
Q_BUF U344 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][7] ));
Q_BUF U345 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][6] ));
Q_BUF U346 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][5] ));
Q_BUF U347 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][4] ));
Q_BUF U348 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][3] ));
Q_BUF U349 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][2] ));
Q_BUF U350 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][1] ));
Q_BUF U351 ( .A(n2), .Z(\sa_ctrl_rst_dat[21][0] ));
Q_BUF U352 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][31] ));
Q_BUF U353 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][30] ));
Q_BUF U354 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][29] ));
Q_BUF U355 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][28] ));
Q_BUF U356 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][27] ));
Q_BUF U357 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][26] ));
Q_BUF U358 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][25] ));
Q_BUF U359 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][24] ));
Q_BUF U360 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][23] ));
Q_BUF U361 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][22] ));
Q_BUF U362 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][21] ));
Q_BUF U363 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][20] ));
Q_BUF U364 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][19] ));
Q_BUF U365 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][18] ));
Q_BUF U366 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][17] ));
Q_BUF U367 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][16] ));
Q_BUF U368 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][15] ));
Q_BUF U369 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][14] ));
Q_BUF U370 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][13] ));
Q_BUF U371 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][12] ));
Q_BUF U372 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][11] ));
Q_BUF U373 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][10] ));
Q_BUF U374 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][9] ));
Q_BUF U375 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][8] ));
Q_BUF U376 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][7] ));
Q_BUF U377 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][6] ));
Q_BUF U378 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][5] ));
Q_BUF U379 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][4] ));
Q_BUF U380 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][3] ));
Q_BUF U381 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][2] ));
Q_BUF U382 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][1] ));
Q_BUF U383 ( .A(n2), .Z(\sa_ctrl_rst_dat[20][0] ));
Q_BUF U384 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][31] ));
Q_BUF U385 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][30] ));
Q_BUF U386 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][29] ));
Q_BUF U387 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][28] ));
Q_BUF U388 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][27] ));
Q_BUF U389 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][26] ));
Q_BUF U390 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][25] ));
Q_BUF U391 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][24] ));
Q_BUF U392 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][23] ));
Q_BUF U393 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][22] ));
Q_BUF U394 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][21] ));
Q_BUF U395 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][20] ));
Q_BUF U396 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][19] ));
Q_BUF U397 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][18] ));
Q_BUF U398 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][17] ));
Q_BUF U399 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][16] ));
Q_BUF U400 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][15] ));
Q_BUF U401 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][14] ));
Q_BUF U402 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][13] ));
Q_BUF U403 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][12] ));
Q_BUF U404 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][11] ));
Q_BUF U405 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][10] ));
Q_BUF U406 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][9] ));
Q_BUF U407 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][8] ));
Q_BUF U408 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][7] ));
Q_BUF U409 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][6] ));
Q_BUF U410 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][5] ));
Q_BUF U411 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][4] ));
Q_BUF U412 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][3] ));
Q_BUF U413 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][2] ));
Q_BUF U414 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][1] ));
Q_BUF U415 ( .A(n2), .Z(\sa_ctrl_rst_dat[19][0] ));
Q_BUF U416 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][31] ));
Q_BUF U417 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][30] ));
Q_BUF U418 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][29] ));
Q_BUF U419 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][28] ));
Q_BUF U420 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][27] ));
Q_BUF U421 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][26] ));
Q_BUF U422 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][25] ));
Q_BUF U423 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][24] ));
Q_BUF U424 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][23] ));
Q_BUF U425 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][22] ));
Q_BUF U426 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][21] ));
Q_BUF U427 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][20] ));
Q_BUF U428 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][19] ));
Q_BUF U429 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][18] ));
Q_BUF U430 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][17] ));
Q_BUF U431 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][16] ));
Q_BUF U432 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][15] ));
Q_BUF U433 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][14] ));
Q_BUF U434 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][13] ));
Q_BUF U435 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][12] ));
Q_BUF U436 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][11] ));
Q_BUF U437 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][10] ));
Q_BUF U438 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][9] ));
Q_BUF U439 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][8] ));
Q_BUF U440 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][7] ));
Q_BUF U441 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][6] ));
Q_BUF U442 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][5] ));
Q_BUF U443 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][4] ));
Q_BUF U444 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][3] ));
Q_BUF U445 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][2] ));
Q_BUF U446 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][1] ));
Q_BUF U447 ( .A(n2), .Z(\sa_ctrl_rst_dat[18][0] ));
Q_BUF U448 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][31] ));
Q_BUF U449 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][30] ));
Q_BUF U450 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][29] ));
Q_BUF U451 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][28] ));
Q_BUF U452 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][27] ));
Q_BUF U453 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][26] ));
Q_BUF U454 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][25] ));
Q_BUF U455 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][24] ));
Q_BUF U456 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][23] ));
Q_BUF U457 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][22] ));
Q_BUF U458 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][21] ));
Q_BUF U459 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][20] ));
Q_BUF U460 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][19] ));
Q_BUF U461 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][18] ));
Q_BUF U462 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][17] ));
Q_BUF U463 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][16] ));
Q_BUF U464 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][15] ));
Q_BUF U465 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][14] ));
Q_BUF U466 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][13] ));
Q_BUF U467 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][12] ));
Q_BUF U468 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][11] ));
Q_BUF U469 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][10] ));
Q_BUF U470 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][9] ));
Q_BUF U471 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][8] ));
Q_BUF U472 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][7] ));
Q_BUF U473 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][6] ));
Q_BUF U474 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][5] ));
Q_BUF U475 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][4] ));
Q_BUF U476 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][3] ));
Q_BUF U477 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][2] ));
Q_BUF U478 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][1] ));
Q_BUF U479 ( .A(n2), .Z(\sa_ctrl_rst_dat[17][0] ));
Q_BUF U480 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][31] ));
Q_BUF U481 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][30] ));
Q_BUF U482 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][29] ));
Q_BUF U483 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][28] ));
Q_BUF U484 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][27] ));
Q_BUF U485 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][26] ));
Q_BUF U486 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][25] ));
Q_BUF U487 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][24] ));
Q_BUF U488 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][23] ));
Q_BUF U489 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][22] ));
Q_BUF U490 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][21] ));
Q_BUF U491 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][20] ));
Q_BUF U492 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][19] ));
Q_BUF U493 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][18] ));
Q_BUF U494 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][17] ));
Q_BUF U495 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][16] ));
Q_BUF U496 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][15] ));
Q_BUF U497 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][14] ));
Q_BUF U498 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][13] ));
Q_BUF U499 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][12] ));
Q_BUF U500 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][11] ));
Q_BUF U501 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][10] ));
Q_BUF U502 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][9] ));
Q_BUF U503 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][8] ));
Q_BUF U504 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][7] ));
Q_BUF U505 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][6] ));
Q_BUF U506 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][5] ));
Q_BUF U507 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][4] ));
Q_BUF U508 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][3] ));
Q_BUF U509 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][2] ));
Q_BUF U510 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][1] ));
Q_BUF U511 ( .A(n2), .Z(\sa_ctrl_rst_dat[16][0] ));
Q_BUF U512 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][31] ));
Q_BUF U513 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][30] ));
Q_BUF U514 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][29] ));
Q_BUF U515 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][28] ));
Q_BUF U516 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][27] ));
Q_BUF U517 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][26] ));
Q_BUF U518 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][25] ));
Q_BUF U519 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][24] ));
Q_BUF U520 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][23] ));
Q_BUF U521 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][22] ));
Q_BUF U522 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][21] ));
Q_BUF U523 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][20] ));
Q_BUF U524 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][19] ));
Q_BUF U525 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][18] ));
Q_BUF U526 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][17] ));
Q_BUF U527 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][16] ));
Q_BUF U528 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][15] ));
Q_BUF U529 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][14] ));
Q_BUF U530 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][13] ));
Q_BUF U531 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][12] ));
Q_BUF U532 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][11] ));
Q_BUF U533 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][10] ));
Q_BUF U534 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][9] ));
Q_BUF U535 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][8] ));
Q_BUF U536 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][7] ));
Q_BUF U537 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][6] ));
Q_BUF U538 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][5] ));
Q_BUF U539 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][4] ));
Q_BUF U540 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][3] ));
Q_BUF U541 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][2] ));
Q_BUF U542 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][1] ));
Q_BUF U543 ( .A(n2), .Z(\sa_ctrl_rst_dat[15][0] ));
Q_BUF U544 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][31] ));
Q_BUF U545 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][30] ));
Q_BUF U546 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][29] ));
Q_BUF U547 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][28] ));
Q_BUF U548 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][27] ));
Q_BUF U549 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][26] ));
Q_BUF U550 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][25] ));
Q_BUF U551 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][24] ));
Q_BUF U552 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][23] ));
Q_BUF U553 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][22] ));
Q_BUF U554 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][21] ));
Q_BUF U555 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][20] ));
Q_BUF U556 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][19] ));
Q_BUF U557 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][18] ));
Q_BUF U558 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][17] ));
Q_BUF U559 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][16] ));
Q_BUF U560 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][15] ));
Q_BUF U561 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][14] ));
Q_BUF U562 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][13] ));
Q_BUF U563 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][12] ));
Q_BUF U564 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][11] ));
Q_BUF U565 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][10] ));
Q_BUF U566 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][9] ));
Q_BUF U567 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][8] ));
Q_BUF U568 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][7] ));
Q_BUF U569 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][6] ));
Q_BUF U570 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][5] ));
Q_BUF U571 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][4] ));
Q_BUF U572 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][3] ));
Q_BUF U573 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][2] ));
Q_BUF U574 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][1] ));
Q_BUF U575 ( .A(n2), .Z(\sa_ctrl_rst_dat[14][0] ));
Q_BUF U576 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][31] ));
Q_BUF U577 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][30] ));
Q_BUF U578 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][29] ));
Q_BUF U579 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][28] ));
Q_BUF U580 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][27] ));
Q_BUF U581 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][26] ));
Q_BUF U582 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][25] ));
Q_BUF U583 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][24] ));
Q_BUF U584 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][23] ));
Q_BUF U585 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][22] ));
Q_BUF U586 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][21] ));
Q_BUF U587 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][20] ));
Q_BUF U588 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][19] ));
Q_BUF U589 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][18] ));
Q_BUF U590 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][17] ));
Q_BUF U591 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][16] ));
Q_BUF U592 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][15] ));
Q_BUF U593 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][14] ));
Q_BUF U594 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][13] ));
Q_BUF U595 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][12] ));
Q_BUF U596 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][11] ));
Q_BUF U597 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][10] ));
Q_BUF U598 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][9] ));
Q_BUF U599 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][8] ));
Q_BUF U600 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][7] ));
Q_BUF U601 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][6] ));
Q_BUF U602 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][5] ));
Q_BUF U603 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][4] ));
Q_BUF U604 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][3] ));
Q_BUF U605 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][2] ));
Q_BUF U606 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][1] ));
Q_BUF U607 ( .A(n2), .Z(\sa_ctrl_rst_dat[13][0] ));
Q_BUF U608 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][31] ));
Q_BUF U609 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][30] ));
Q_BUF U610 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][29] ));
Q_BUF U611 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][28] ));
Q_BUF U612 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][27] ));
Q_BUF U613 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][26] ));
Q_BUF U614 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][25] ));
Q_BUF U615 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][24] ));
Q_BUF U616 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][23] ));
Q_BUF U617 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][22] ));
Q_BUF U618 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][21] ));
Q_BUF U619 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][20] ));
Q_BUF U620 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][19] ));
Q_BUF U621 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][18] ));
Q_BUF U622 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][17] ));
Q_BUF U623 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][16] ));
Q_BUF U624 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][15] ));
Q_BUF U625 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][14] ));
Q_BUF U626 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][13] ));
Q_BUF U627 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][12] ));
Q_BUF U628 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][11] ));
Q_BUF U629 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][10] ));
Q_BUF U630 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][9] ));
Q_BUF U631 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][8] ));
Q_BUF U632 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][7] ));
Q_BUF U633 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][6] ));
Q_BUF U634 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][5] ));
Q_BUF U635 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][4] ));
Q_BUF U636 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][3] ));
Q_BUF U637 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][2] ));
Q_BUF U638 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][1] ));
Q_BUF U639 ( .A(n2), .Z(\sa_ctrl_rst_dat[12][0] ));
Q_BUF U640 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][31] ));
Q_BUF U641 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][30] ));
Q_BUF U642 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][29] ));
Q_BUF U643 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][28] ));
Q_BUF U644 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][27] ));
Q_BUF U645 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][26] ));
Q_BUF U646 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][25] ));
Q_BUF U647 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][24] ));
Q_BUF U648 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][23] ));
Q_BUF U649 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][22] ));
Q_BUF U650 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][21] ));
Q_BUF U651 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][20] ));
Q_BUF U652 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][19] ));
Q_BUF U653 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][18] ));
Q_BUF U654 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][17] ));
Q_BUF U655 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][16] ));
Q_BUF U656 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][15] ));
Q_BUF U657 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][14] ));
Q_BUF U658 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][13] ));
Q_BUF U659 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][12] ));
Q_BUF U660 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][11] ));
Q_BUF U661 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][10] ));
Q_BUF U662 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][9] ));
Q_BUF U663 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][8] ));
Q_BUF U664 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][7] ));
Q_BUF U665 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][6] ));
Q_BUF U666 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][5] ));
Q_BUF U667 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][4] ));
Q_BUF U668 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][3] ));
Q_BUF U669 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][2] ));
Q_BUF U670 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][1] ));
Q_BUF U671 ( .A(n2), .Z(\sa_ctrl_rst_dat[11][0] ));
Q_BUF U672 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][31] ));
Q_BUF U673 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][30] ));
Q_BUF U674 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][29] ));
Q_BUF U675 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][28] ));
Q_BUF U676 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][27] ));
Q_BUF U677 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][26] ));
Q_BUF U678 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][25] ));
Q_BUF U679 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][24] ));
Q_BUF U680 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][23] ));
Q_BUF U681 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][22] ));
Q_BUF U682 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][21] ));
Q_BUF U683 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][20] ));
Q_BUF U684 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][19] ));
Q_BUF U685 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][18] ));
Q_BUF U686 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][17] ));
Q_BUF U687 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][16] ));
Q_BUF U688 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][15] ));
Q_BUF U689 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][14] ));
Q_BUF U690 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][13] ));
Q_BUF U691 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][12] ));
Q_BUF U692 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][11] ));
Q_BUF U693 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][10] ));
Q_BUF U694 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][9] ));
Q_BUF U695 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][8] ));
Q_BUF U696 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][7] ));
Q_BUF U697 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][6] ));
Q_BUF U698 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][5] ));
Q_BUF U699 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][4] ));
Q_BUF U700 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][3] ));
Q_BUF U701 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][2] ));
Q_BUF U702 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][1] ));
Q_BUF U703 ( .A(n2), .Z(\sa_ctrl_rst_dat[10][0] ));
Q_BUF U704 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][31] ));
Q_BUF U705 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][30] ));
Q_BUF U706 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][29] ));
Q_BUF U707 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][28] ));
Q_BUF U708 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][27] ));
Q_BUF U709 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][26] ));
Q_BUF U710 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][25] ));
Q_BUF U711 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][24] ));
Q_BUF U712 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][23] ));
Q_BUF U713 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][22] ));
Q_BUF U714 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][21] ));
Q_BUF U715 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][20] ));
Q_BUF U716 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][19] ));
Q_BUF U717 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][18] ));
Q_BUF U718 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][17] ));
Q_BUF U719 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][16] ));
Q_BUF U720 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][15] ));
Q_BUF U721 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][14] ));
Q_BUF U722 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][13] ));
Q_BUF U723 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][12] ));
Q_BUF U724 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][11] ));
Q_BUF U725 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][10] ));
Q_BUF U726 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][9] ));
Q_BUF U727 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][8] ));
Q_BUF U728 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][7] ));
Q_BUF U729 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][6] ));
Q_BUF U730 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][5] ));
Q_BUF U731 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][4] ));
Q_BUF U732 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][3] ));
Q_BUF U733 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][2] ));
Q_BUF U734 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][1] ));
Q_BUF U735 ( .A(n2), .Z(\sa_ctrl_rst_dat[9][0] ));
Q_BUF U736 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][31] ));
Q_BUF U737 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][30] ));
Q_BUF U738 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][29] ));
Q_BUF U739 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][28] ));
Q_BUF U740 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][27] ));
Q_BUF U741 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][26] ));
Q_BUF U742 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][25] ));
Q_BUF U743 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][24] ));
Q_BUF U744 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][23] ));
Q_BUF U745 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][22] ));
Q_BUF U746 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][21] ));
Q_BUF U747 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][20] ));
Q_BUF U748 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][19] ));
Q_BUF U749 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][18] ));
Q_BUF U750 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][17] ));
Q_BUF U751 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][16] ));
Q_BUF U752 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][15] ));
Q_BUF U753 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][14] ));
Q_BUF U754 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][13] ));
Q_BUF U755 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][12] ));
Q_BUF U756 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][11] ));
Q_BUF U757 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][10] ));
Q_BUF U758 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][9] ));
Q_BUF U759 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][8] ));
Q_BUF U760 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][7] ));
Q_BUF U761 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][6] ));
Q_BUF U762 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][5] ));
Q_BUF U763 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][4] ));
Q_BUF U764 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][3] ));
Q_BUF U765 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][2] ));
Q_BUF U766 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][1] ));
Q_BUF U767 ( .A(n2), .Z(\sa_ctrl_rst_dat[8][0] ));
Q_BUF U768 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][31] ));
Q_BUF U769 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][30] ));
Q_BUF U770 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][29] ));
Q_BUF U771 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][28] ));
Q_BUF U772 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][27] ));
Q_BUF U773 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][26] ));
Q_BUF U774 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][25] ));
Q_BUF U775 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][24] ));
Q_BUF U776 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][23] ));
Q_BUF U777 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][22] ));
Q_BUF U778 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][21] ));
Q_BUF U779 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][20] ));
Q_BUF U780 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][19] ));
Q_BUF U781 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][18] ));
Q_BUF U782 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][17] ));
Q_BUF U783 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][16] ));
Q_BUF U784 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][15] ));
Q_BUF U785 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][14] ));
Q_BUF U786 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][13] ));
Q_BUF U787 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][12] ));
Q_BUF U788 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][11] ));
Q_BUF U789 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][10] ));
Q_BUF U790 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][9] ));
Q_BUF U791 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][8] ));
Q_BUF U792 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][7] ));
Q_BUF U793 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][6] ));
Q_BUF U794 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][5] ));
Q_BUF U795 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][4] ));
Q_BUF U796 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][3] ));
Q_BUF U797 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][2] ));
Q_BUF U798 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][1] ));
Q_BUF U799 ( .A(n2), .Z(\sa_ctrl_rst_dat[7][0] ));
Q_BUF U800 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][31] ));
Q_BUF U801 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][30] ));
Q_BUF U802 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][29] ));
Q_BUF U803 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][28] ));
Q_BUF U804 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][27] ));
Q_BUF U805 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][26] ));
Q_BUF U806 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][25] ));
Q_BUF U807 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][24] ));
Q_BUF U808 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][23] ));
Q_BUF U809 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][22] ));
Q_BUF U810 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][21] ));
Q_BUF U811 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][20] ));
Q_BUF U812 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][19] ));
Q_BUF U813 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][18] ));
Q_BUF U814 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][17] ));
Q_BUF U815 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][16] ));
Q_BUF U816 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][15] ));
Q_BUF U817 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][14] ));
Q_BUF U818 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][13] ));
Q_BUF U819 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][12] ));
Q_BUF U820 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][11] ));
Q_BUF U821 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][10] ));
Q_BUF U822 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][9] ));
Q_BUF U823 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][8] ));
Q_BUF U824 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][7] ));
Q_BUF U825 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][6] ));
Q_BUF U826 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][5] ));
Q_BUF U827 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][4] ));
Q_BUF U828 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][3] ));
Q_BUF U829 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][2] ));
Q_BUF U830 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][1] ));
Q_BUF U831 ( .A(n2), .Z(\sa_ctrl_rst_dat[6][0] ));
Q_BUF U832 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][31] ));
Q_BUF U833 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][30] ));
Q_BUF U834 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][29] ));
Q_BUF U835 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][28] ));
Q_BUF U836 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][27] ));
Q_BUF U837 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][26] ));
Q_BUF U838 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][25] ));
Q_BUF U839 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][24] ));
Q_BUF U840 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][23] ));
Q_BUF U841 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][22] ));
Q_BUF U842 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][21] ));
Q_BUF U843 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][20] ));
Q_BUF U844 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][19] ));
Q_BUF U845 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][18] ));
Q_BUF U846 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][17] ));
Q_BUF U847 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][16] ));
Q_BUF U848 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][15] ));
Q_BUF U849 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][14] ));
Q_BUF U850 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][13] ));
Q_BUF U851 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][12] ));
Q_BUF U852 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][11] ));
Q_BUF U853 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][10] ));
Q_BUF U854 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][9] ));
Q_BUF U855 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][8] ));
Q_BUF U856 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][7] ));
Q_BUF U857 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][6] ));
Q_BUF U858 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][5] ));
Q_BUF U859 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][4] ));
Q_BUF U860 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][3] ));
Q_BUF U861 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][2] ));
Q_BUF U862 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][1] ));
Q_BUF U863 ( .A(n2), .Z(\sa_ctrl_rst_dat[5][0] ));
Q_BUF U864 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][31] ));
Q_BUF U865 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][30] ));
Q_BUF U866 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][29] ));
Q_BUF U867 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][28] ));
Q_BUF U868 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][27] ));
Q_BUF U869 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][26] ));
Q_BUF U870 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][25] ));
Q_BUF U871 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][24] ));
Q_BUF U872 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][23] ));
Q_BUF U873 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][22] ));
Q_BUF U874 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][21] ));
Q_BUF U875 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][20] ));
Q_BUF U876 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][19] ));
Q_BUF U877 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][18] ));
Q_BUF U878 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][17] ));
Q_BUF U879 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][16] ));
Q_BUF U880 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][15] ));
Q_BUF U881 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][14] ));
Q_BUF U882 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][13] ));
Q_BUF U883 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][12] ));
Q_BUF U884 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][11] ));
Q_BUF U885 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][10] ));
Q_BUF U886 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][9] ));
Q_BUF U887 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][8] ));
Q_BUF U888 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][7] ));
Q_BUF U889 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][6] ));
Q_BUF U890 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][5] ));
Q_BUF U891 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][4] ));
Q_BUF U892 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][3] ));
Q_BUF U893 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][2] ));
Q_BUF U894 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][1] ));
Q_BUF U895 ( .A(n2), .Z(\sa_ctrl_rst_dat[4][0] ));
Q_BUF U896 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][31] ));
Q_BUF U897 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][30] ));
Q_BUF U898 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][29] ));
Q_BUF U899 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][28] ));
Q_BUF U900 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][27] ));
Q_BUF U901 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][26] ));
Q_BUF U902 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][25] ));
Q_BUF U903 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][24] ));
Q_BUF U904 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][23] ));
Q_BUF U905 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][22] ));
Q_BUF U906 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][21] ));
Q_BUF U907 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][20] ));
Q_BUF U908 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][19] ));
Q_BUF U909 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][18] ));
Q_BUF U910 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][17] ));
Q_BUF U911 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][16] ));
Q_BUF U912 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][15] ));
Q_BUF U913 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][14] ));
Q_BUF U914 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][13] ));
Q_BUF U915 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][12] ));
Q_BUF U916 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][11] ));
Q_BUF U917 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][10] ));
Q_BUF U918 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][9] ));
Q_BUF U919 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][8] ));
Q_BUF U920 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][7] ));
Q_BUF U921 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][6] ));
Q_BUF U922 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][5] ));
Q_BUF U923 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][4] ));
Q_BUF U924 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][3] ));
Q_BUF U925 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][2] ));
Q_BUF U926 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][1] ));
Q_BUF U927 ( .A(n2), .Z(\sa_ctrl_rst_dat[3][0] ));
Q_BUF U928 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][31] ));
Q_BUF U929 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][30] ));
Q_BUF U930 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][29] ));
Q_BUF U931 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][28] ));
Q_BUF U932 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][27] ));
Q_BUF U933 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][26] ));
Q_BUF U934 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][25] ));
Q_BUF U935 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][24] ));
Q_BUF U936 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][23] ));
Q_BUF U937 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][22] ));
Q_BUF U938 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][21] ));
Q_BUF U939 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][20] ));
Q_BUF U940 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][19] ));
Q_BUF U941 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][18] ));
Q_BUF U942 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][17] ));
Q_BUF U943 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][16] ));
Q_BUF U944 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][15] ));
Q_BUF U945 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][14] ));
Q_BUF U946 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][13] ));
Q_BUF U947 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][12] ));
Q_BUF U948 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][11] ));
Q_BUF U949 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][10] ));
Q_BUF U950 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][9] ));
Q_BUF U951 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][8] ));
Q_BUF U952 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][7] ));
Q_BUF U953 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][6] ));
Q_BUF U954 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][5] ));
Q_BUF U955 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][4] ));
Q_BUF U956 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][3] ));
Q_BUF U957 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][2] ));
Q_BUF U958 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][1] ));
Q_BUF U959 ( .A(n2), .Z(\sa_ctrl_rst_dat[2][0] ));
Q_BUF U960 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][31] ));
Q_BUF U961 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][30] ));
Q_BUF U962 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][29] ));
Q_BUF U963 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][28] ));
Q_BUF U964 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][27] ));
Q_BUF U965 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][26] ));
Q_BUF U966 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][25] ));
Q_BUF U967 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][24] ));
Q_BUF U968 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][23] ));
Q_BUF U969 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][22] ));
Q_BUF U970 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][21] ));
Q_BUF U971 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][20] ));
Q_BUF U972 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][19] ));
Q_BUF U973 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][18] ));
Q_BUF U974 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][17] ));
Q_BUF U975 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][16] ));
Q_BUF U976 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][15] ));
Q_BUF U977 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][14] ));
Q_BUF U978 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][13] ));
Q_BUF U979 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][12] ));
Q_BUF U980 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][11] ));
Q_BUF U981 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][10] ));
Q_BUF U982 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][9] ));
Q_BUF U983 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][8] ));
Q_BUF U984 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][7] ));
Q_BUF U985 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][6] ));
Q_BUF U986 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][5] ));
Q_BUF U987 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][4] ));
Q_BUF U988 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][3] ));
Q_BUF U989 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][2] ));
Q_BUF U990 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][1] ));
Q_BUF U991 ( .A(n2), .Z(\sa_ctrl_rst_dat[1][0] ));
Q_BUF U992 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][31] ));
Q_BUF U993 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][30] ));
Q_BUF U994 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][29] ));
Q_BUF U995 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][28] ));
Q_BUF U996 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][27] ));
Q_BUF U997 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][26] ));
Q_BUF U998 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][25] ));
Q_BUF U999 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][24] ));
Q_BUF U1000 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][23] ));
Q_BUF U1001 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][22] ));
Q_BUF U1002 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][21] ));
Q_BUF U1003 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][20] ));
Q_BUF U1004 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][19] ));
Q_BUF U1005 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][18] ));
Q_BUF U1006 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][17] ));
Q_BUF U1007 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][16] ));
Q_BUF U1008 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][15] ));
Q_BUF U1009 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][14] ));
Q_BUF U1010 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][13] ));
Q_BUF U1011 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][12] ));
Q_BUF U1012 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][11] ));
Q_BUF U1013 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][10] ));
Q_BUF U1014 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][9] ));
Q_BUF U1015 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][8] ));
Q_BUF U1016 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][7] ));
Q_BUF U1017 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][6] ));
Q_BUF U1018 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][5] ));
Q_BUF U1019 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][4] ));
Q_BUF U1020 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][3] ));
Q_BUF U1021 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][2] ));
Q_BUF U1022 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][1] ));
Q_BUF U1023 ( .A(n2), .Z(\sa_ctrl_rst_dat[0][0] ));
Q_BUF U1024 ( .A(n2), .Z(_zy_simnet_cio_681[37]));
Q_BUF U1025 ( .A(n2), .Z(_zy_simnet_cio_681[36]));
Q_BUF U1026 ( .A(n2), .Z(_zy_simnet_cio_681[35]));
Q_BUF U1027 ( .A(n2), .Z(_zy_simnet_cio_681[34]));
Q_BUF U1028 ( .A(n2), .Z(_zy_simnet_cio_681[33]));
Q_BUF U1029 ( .A(n2), .Z(_zy_simnet_cio_681[32]));
Q_BUF U1030 ( .A(n2), .Z(_zy_simnet_cio_681[31]));
Q_BUF U1031 ( .A(n2), .Z(_zy_simnet_cio_681[30]));
Q_BUF U1032 ( .A(n2), .Z(_zy_simnet_cio_681[29]));
Q_BUF U1033 ( .A(n2), .Z(_zy_simnet_cio_681[28]));
Q_BUF U1034 ( .A(n2), .Z(_zy_simnet_cio_681[27]));
Q_BUF U1035 ( .A(n2), .Z(_zy_simnet_cio_681[26]));
Q_BUF U1036 ( .A(n2), .Z(_zy_simnet_cio_681[25]));
Q_BUF U1037 ( .A(n2), .Z(_zy_simnet_cio_681[24]));
Q_BUF U1038 ( .A(n2), .Z(_zy_simnet_cio_681[23]));
Q_BUF U1039 ( .A(n2), .Z(_zy_simnet_cio_681[22]));
Q_BUF U1040 ( .A(n2), .Z(_zy_simnet_cio_681[21]));
Q_BUF U1041 ( .A(n2), .Z(_zy_simnet_cio_681[20]));
Q_BUF U1042 ( .A(n2), .Z(_zy_simnet_cio_681[19]));
Q_BUF U1043 ( .A(n2), .Z(_zy_simnet_cio_681[18]));
Q_BUF U1044 ( .A(n2), .Z(_zy_simnet_cio_681[17]));
Q_BUF U1045 ( .A(n2), .Z(_zy_simnet_cio_681[16]));
Q_BUF U1046 ( .A(n2), .Z(_zy_simnet_cio_681[15]));
Q_BUF U1047 ( .A(n2), .Z(_zy_simnet_cio_681[14]));
Q_BUF U1048 ( .A(n2), .Z(_zy_simnet_cio_681[13]));
Q_BUF U1049 ( .A(n2), .Z(_zy_simnet_cio_681[12]));
Q_BUF U1050 ( .A(n2), .Z(_zy_simnet_cio_681[11]));
Q_BUF U1051 ( .A(n2), .Z(_zy_simnet_cio_681[10]));
Q_BUF U1052 ( .A(n2), .Z(_zy_simnet_cio_681[9]));
Q_BUF U1053 ( .A(n2), .Z(_zy_simnet_cio_681[8]));
Q_BUF U1054 ( .A(n2), .Z(_zy_simnet_cio_681[7]));
Q_BUF U1055 ( .A(n2), .Z(_zy_simnet_cio_681[6]));
Q_BUF U1056 ( .A(n2), .Z(_zy_simnet_cio_681[5]));
Q_BUF U1057 ( .A(n2), .Z(_zy_simnet_cio_681[4]));
Q_BUF U1058 ( .A(n2), .Z(_zy_simnet_cio_681[3]));
Q_BUF U1059 ( .A(n2), .Z(_zy_simnet_cio_681[2]));
Q_BUF U1060 ( .A(n2), .Z(_zy_simnet_cio_681[1]));
Q_BUF U1061 ( .A(n2), .Z(_zy_simnet_cio_681[0]));
Q_BUF U1062 ( .A(n2), .Z(_zy_simnet_cio_680[37]));
Q_BUF U1063 ( .A(n2), .Z(_zy_simnet_cio_680[36]));
Q_BUF U1064 ( .A(n2), .Z(_zy_simnet_cio_680[35]));
Q_BUF U1065 ( .A(n2), .Z(_zy_simnet_cio_680[34]));
Q_BUF U1066 ( .A(n2), .Z(_zy_simnet_cio_680[33]));
Q_BUF U1067 ( .A(n2), .Z(_zy_simnet_cio_680[32]));
Q_BUF U1068 ( .A(n2), .Z(_zy_simnet_cio_680[31]));
Q_BUF U1069 ( .A(n2), .Z(_zy_simnet_cio_680[30]));
Q_BUF U1070 ( .A(n2), .Z(_zy_simnet_cio_680[29]));
Q_BUF U1071 ( .A(n2), .Z(_zy_simnet_cio_680[28]));
Q_BUF U1072 ( .A(n2), .Z(_zy_simnet_cio_680[27]));
Q_BUF U1073 ( .A(n2), .Z(_zy_simnet_cio_680[26]));
Q_BUF U1074 ( .A(n2), .Z(_zy_simnet_cio_680[25]));
Q_BUF U1075 ( .A(n2), .Z(_zy_simnet_cio_680[24]));
Q_BUF U1076 ( .A(n2), .Z(_zy_simnet_cio_680[23]));
Q_BUF U1077 ( .A(n2), .Z(_zy_simnet_cio_680[22]));
Q_BUF U1078 ( .A(n2), .Z(_zy_simnet_cio_680[21]));
Q_BUF U1079 ( .A(n2), .Z(_zy_simnet_cio_680[20]));
Q_BUF U1080 ( .A(n2), .Z(_zy_simnet_cio_680[19]));
Q_BUF U1081 ( .A(n2), .Z(_zy_simnet_cio_680[18]));
Q_BUF U1082 ( .A(n2), .Z(_zy_simnet_cio_680[17]));
Q_BUF U1083 ( .A(n2), .Z(_zy_simnet_cio_680[16]));
Q_BUF U1084 ( .A(n2), .Z(_zy_simnet_cio_680[15]));
Q_BUF U1085 ( .A(n2), .Z(_zy_simnet_cio_680[14]));
Q_BUF U1086 ( .A(n2), .Z(_zy_simnet_cio_680[13]));
Q_BUF U1087 ( .A(n2), .Z(_zy_simnet_cio_680[12]));
Q_BUF U1088 ( .A(n2), .Z(_zy_simnet_cio_680[11]));
Q_BUF U1089 ( .A(n2), .Z(_zy_simnet_cio_680[10]));
Q_BUF U1090 ( .A(n2), .Z(_zy_simnet_cio_680[9]));
Q_BUF U1091 ( .A(n2), .Z(_zy_simnet_cio_680[8]));
Q_BUF U1092 ( .A(n2), .Z(_zy_simnet_cio_680[7]));
Q_BUF U1093 ( .A(n2), .Z(_zy_simnet_cio_680[6]));
Q_BUF U1094 ( .A(n2), .Z(_zy_simnet_cio_680[5]));
Q_BUF U1095 ( .A(n2), .Z(_zy_simnet_cio_680[4]));
Q_BUF U1096 ( .A(n2), .Z(_zy_simnet_cio_680[3]));
Q_BUF U1097 ( .A(n2), .Z(_zy_simnet_cio_680[2]));
Q_BUF U1098 ( .A(n2), .Z(_zy_simnet_cio_680[1]));
Q_BUF U1099 ( .A(n2), .Z(_zy_simnet_cio_680[0]));
Q_BUF U1100 ( .A(n2), .Z(_zy_simnet_cio_679));
Q_BUF U1101 ( .A(n2), .Z(_zy_simnet_cio_674));
Q_BUF U1102 ( .A(n2), .Z(_zy_simnet_cio_661[63]));
Q_BUF U1103 ( .A(n2), .Z(_zy_simnet_cio_661[62]));
Q_BUF U1104 ( .A(n2), .Z(_zy_simnet_cio_661[61]));
Q_BUF U1105 ( .A(n2), .Z(_zy_simnet_cio_661[60]));
Q_BUF U1106 ( .A(n2), .Z(_zy_simnet_cio_661[59]));
Q_BUF U1107 ( .A(n2), .Z(_zy_simnet_cio_661[58]));
Q_BUF U1108 ( .A(n2), .Z(_zy_simnet_cio_661[57]));
Q_BUF U1109 ( .A(n2), .Z(_zy_simnet_cio_661[56]));
Q_BUF U1110 ( .A(n2), .Z(_zy_simnet_cio_661[55]));
Q_BUF U1111 ( .A(n2), .Z(_zy_simnet_cio_661[54]));
Q_BUF U1112 ( .A(n2), .Z(_zy_simnet_cio_661[53]));
Q_BUF U1113 ( .A(n2), .Z(_zy_simnet_cio_661[52]));
Q_BUF U1114 ( .A(n2), .Z(_zy_simnet_cio_661[51]));
Q_BUF U1115 ( .A(n2), .Z(_zy_simnet_cio_661[50]));
Q_BUF U1116 ( .A(n2), .Z(_zy_simnet_cio_661[49]));
Q_BUF U1117 ( .A(n2), .Z(_zy_simnet_cio_661[48]));
Q_BUF U1118 ( .A(n2), .Z(_zy_simnet_cio_661[47]));
Q_BUF U1119 ( .A(n2), .Z(_zy_simnet_cio_661[46]));
Q_BUF U1120 ( .A(n2), .Z(_zy_simnet_cio_661[45]));
Q_BUF U1121 ( .A(n2), .Z(_zy_simnet_cio_661[44]));
Q_BUF U1122 ( .A(n2), .Z(_zy_simnet_cio_661[43]));
Q_BUF U1123 ( .A(n2), .Z(_zy_simnet_cio_661[42]));
Q_BUF U1124 ( .A(n2), .Z(_zy_simnet_cio_661[41]));
Q_BUF U1125 ( .A(n2), .Z(_zy_simnet_cio_661[40]));
Q_BUF U1126 ( .A(n2), .Z(_zy_simnet_cio_661[39]));
Q_BUF U1127 ( .A(n2), .Z(_zy_simnet_cio_661[38]));
Q_BUF U1128 ( .A(n2), .Z(_zy_simnet_cio_661[37]));
Q_BUF U1129 ( .A(n2), .Z(_zy_simnet_cio_661[36]));
Q_BUF U1130 ( .A(n2), .Z(_zy_simnet_cio_661[35]));
Q_BUF U1131 ( .A(n2), .Z(_zy_simnet_cio_661[34]));
Q_BUF U1132 ( .A(n2), .Z(_zy_simnet_cio_661[33]));
Q_BUF U1133 ( .A(n2), .Z(_zy_simnet_cio_661[32]));
Q_BUF U1134 ( .A(n2), .Z(_zy_simnet_cio_661[31]));
Q_BUF U1135 ( .A(n2), .Z(_zy_simnet_cio_661[30]));
Q_BUF U1136 ( .A(n2), .Z(_zy_simnet_cio_661[29]));
Q_BUF U1137 ( .A(n2), .Z(_zy_simnet_cio_661[28]));
Q_BUF U1138 ( .A(n2), .Z(_zy_simnet_cio_661[27]));
Q_BUF U1139 ( .A(n2), .Z(_zy_simnet_cio_661[26]));
Q_BUF U1140 ( .A(n2), .Z(_zy_simnet_cio_661[25]));
Q_BUF U1141 ( .A(n2), .Z(_zy_simnet_cio_661[24]));
Q_BUF U1142 ( .A(n2), .Z(_zy_simnet_cio_661[23]));
Q_BUF U1143 ( .A(n2), .Z(_zy_simnet_cio_661[22]));
Q_BUF U1144 ( .A(n2), .Z(_zy_simnet_cio_661[21]));
Q_BUF U1145 ( .A(n2), .Z(_zy_simnet_cio_661[20]));
Q_BUF U1146 ( .A(n2), .Z(_zy_simnet_cio_661[19]));
Q_BUF U1147 ( .A(n2), .Z(_zy_simnet_cio_661[18]));
Q_BUF U1148 ( .A(n2), .Z(_zy_simnet_cio_661[17]));
Q_BUF U1149 ( .A(n2), .Z(_zy_simnet_cio_661[16]));
Q_BUF U1150 ( .A(n2), .Z(_zy_simnet_cio_661[15]));
Q_BUF U1151 ( .A(n2), .Z(_zy_simnet_cio_661[14]));
Q_BUF U1152 ( .A(n2), .Z(_zy_simnet_cio_661[13]));
Q_BUF U1153 ( .A(n2), .Z(_zy_simnet_cio_661[12]));
Q_BUF U1154 ( .A(n2), .Z(_zy_simnet_cio_661[11]));
Q_BUF U1155 ( .A(n2), .Z(_zy_simnet_cio_661[10]));
Q_BUF U1156 ( .A(n2), .Z(_zy_simnet_cio_661[9]));
Q_BUF U1157 ( .A(n2), .Z(_zy_simnet_cio_661[8]));
Q_BUF U1158 ( .A(n2), .Z(_zy_simnet_cio_661[7]));
Q_BUF U1159 ( .A(n2), .Z(_zy_simnet_cio_661[6]));
Q_BUF U1160 ( .A(n2), .Z(_zy_simnet_cio_661[5]));
Q_BUF U1161 ( .A(n2), .Z(_zy_simnet_cio_661[4]));
Q_BUF U1162 ( .A(n2), .Z(_zy_simnet_cio_661[3]));
Q_BUF U1163 ( .A(n2), .Z(_zy_simnet_cio_661[2]));
Q_BUF U1164 ( .A(n2), .Z(_zy_simnet_cio_661[1]));
Q_BUF U1165 ( .A(n2), .Z(_zy_simnet_cio_661[0]));
Q_BUF U1166 ( .A(n2), .Z(_zy_simnet_cio_660[63]));
Q_BUF U1167 ( .A(n2), .Z(_zy_simnet_cio_660[62]));
Q_BUF U1168 ( .A(n2), .Z(_zy_simnet_cio_660[61]));
Q_BUF U1169 ( .A(n2), .Z(_zy_simnet_cio_660[60]));
Q_BUF U1170 ( .A(n2), .Z(_zy_simnet_cio_660[59]));
Q_BUF U1171 ( .A(n2), .Z(_zy_simnet_cio_660[58]));
Q_BUF U1172 ( .A(n2), .Z(_zy_simnet_cio_660[57]));
Q_BUF U1173 ( .A(n2), .Z(_zy_simnet_cio_660[56]));
Q_BUF U1174 ( .A(n2), .Z(_zy_simnet_cio_660[55]));
Q_BUF U1175 ( .A(n2), .Z(_zy_simnet_cio_660[54]));
Q_BUF U1176 ( .A(n2), .Z(_zy_simnet_cio_660[53]));
Q_BUF U1177 ( .A(n2), .Z(_zy_simnet_cio_660[52]));
Q_BUF U1178 ( .A(n2), .Z(_zy_simnet_cio_660[51]));
Q_BUF U1179 ( .A(n2), .Z(_zy_simnet_cio_660[50]));
Q_BUF U1180 ( .A(n2), .Z(_zy_simnet_cio_660[49]));
Q_BUF U1181 ( .A(n2), .Z(_zy_simnet_cio_660[48]));
Q_BUF U1182 ( .A(n2), .Z(_zy_simnet_cio_660[47]));
Q_BUF U1183 ( .A(n2), .Z(_zy_simnet_cio_660[46]));
Q_BUF U1184 ( .A(n2), .Z(_zy_simnet_cio_660[45]));
Q_BUF U1185 ( .A(n2), .Z(_zy_simnet_cio_660[44]));
Q_BUF U1186 ( .A(n2), .Z(_zy_simnet_cio_660[43]));
Q_BUF U1187 ( .A(n2), .Z(_zy_simnet_cio_660[42]));
Q_BUF U1188 ( .A(n2), .Z(_zy_simnet_cio_660[41]));
Q_BUF U1189 ( .A(n2), .Z(_zy_simnet_cio_660[40]));
Q_BUF U1190 ( .A(n2), .Z(_zy_simnet_cio_660[39]));
Q_BUF U1191 ( .A(n2), .Z(_zy_simnet_cio_660[38]));
Q_BUF U1192 ( .A(n2), .Z(_zy_simnet_cio_660[37]));
Q_BUF U1193 ( .A(n2), .Z(_zy_simnet_cio_660[36]));
Q_BUF U1194 ( .A(n2), .Z(_zy_simnet_cio_660[35]));
Q_BUF U1195 ( .A(n2), .Z(_zy_simnet_cio_660[34]));
Q_BUF U1196 ( .A(n2), .Z(_zy_simnet_cio_660[33]));
Q_BUF U1197 ( .A(n2), .Z(_zy_simnet_cio_660[32]));
Q_BUF U1198 ( .A(n2), .Z(_zy_simnet_cio_660[31]));
Q_BUF U1199 ( .A(n2), .Z(_zy_simnet_cio_660[30]));
Q_BUF U1200 ( .A(n2), .Z(_zy_simnet_cio_660[29]));
Q_BUF U1201 ( .A(n2), .Z(_zy_simnet_cio_660[28]));
Q_BUF U1202 ( .A(n2), .Z(_zy_simnet_cio_660[27]));
Q_BUF U1203 ( .A(n2), .Z(_zy_simnet_cio_660[26]));
Q_BUF U1204 ( .A(n2), .Z(_zy_simnet_cio_660[25]));
Q_BUF U1205 ( .A(n2), .Z(_zy_simnet_cio_660[24]));
Q_BUF U1206 ( .A(n2), .Z(_zy_simnet_cio_660[23]));
Q_BUF U1207 ( .A(n2), .Z(_zy_simnet_cio_660[22]));
Q_BUF U1208 ( .A(n2), .Z(_zy_simnet_cio_660[21]));
Q_BUF U1209 ( .A(n2), .Z(_zy_simnet_cio_660[20]));
Q_BUF U1210 ( .A(n2), .Z(_zy_simnet_cio_660[19]));
Q_BUF U1211 ( .A(n2), .Z(_zy_simnet_cio_660[18]));
Q_BUF U1212 ( .A(n2), .Z(_zy_simnet_cio_660[17]));
Q_BUF U1213 ( .A(n2), .Z(_zy_simnet_cio_660[16]));
Q_BUF U1214 ( .A(n2), .Z(_zy_simnet_cio_660[15]));
Q_BUF U1215 ( .A(n2), .Z(_zy_simnet_cio_660[14]));
Q_BUF U1216 ( .A(n2), .Z(_zy_simnet_cio_660[13]));
Q_BUF U1217 ( .A(n2), .Z(_zy_simnet_cio_660[12]));
Q_BUF U1218 ( .A(n2), .Z(_zy_simnet_cio_660[11]));
Q_BUF U1219 ( .A(n2), .Z(_zy_simnet_cio_660[10]));
Q_BUF U1220 ( .A(n2), .Z(_zy_simnet_cio_660[9]));
Q_BUF U1221 ( .A(n2), .Z(_zy_simnet_cio_660[8]));
Q_BUF U1222 ( .A(n2), .Z(_zy_simnet_cio_660[7]));
Q_BUF U1223 ( .A(n2), .Z(_zy_simnet_cio_660[6]));
Q_BUF U1224 ( .A(n2), .Z(_zy_simnet_cio_660[5]));
Q_BUF U1225 ( .A(n2), .Z(_zy_simnet_cio_660[4]));
Q_BUF U1226 ( .A(n2), .Z(_zy_simnet_cio_660[3]));
Q_BUF U1227 ( .A(n2), .Z(_zy_simnet_cio_660[2]));
Q_BUF U1228 ( .A(n2), .Z(_zy_simnet_cio_660[1]));
Q_BUF U1229 ( .A(n2), .Z(_zy_simnet_cio_660[0]));
Q_BUF U1230 ( .A(n2), .Z(_zy_simnet_cio_659));
Q_BUF U1231 ( .A(n2), .Z(_zy_simnet_cio_654));
Q_BUF U1232 ( .A(n2), .Z(_zy_simnet_cio_573));
Q_BUF U1233 ( .A(n2), .Z(_zy_simnet_cio_549));
Q_BUF U1234 ( .A(n2), .Z(_zy_simnet_cio_525));
Q_BUF U1235 ( .A(n2), .Z(_zy_simnet_cio_501));
Q_BUF U1236 ( .A(n2), .Z(_zy_simnet_cio_477));
Q_BUF U1237 ( .A(n2), .Z(_zy_simnet_cio_453));
Q_BUF U1238 ( .A(n2), .Z(_zy_simnet_cio_429));
Q_BUF U1239 ( .A(n2), .Z(_zy_simnet_cio_405));
Q_BUF U1240 ( .A(n2), .Z(_zy_simnet_cio_315[15]));
Q_BUF U1241 ( .A(n2), .Z(_zy_simnet_cio_315[14]));
Q_BUF U1242 ( .A(n2), .Z(_zy_simnet_cio_315[13]));
Q_BUF U1243 ( .A(n2), .Z(_zy_simnet_cio_315[12]));
Q_BUF U1244 ( .A(n2), .Z(_zy_simnet_cio_315[11]));
Q_BUF U1245 ( .A(n2), .Z(_zy_simnet_cio_315[10]));
Q_BUF U1246 ( .A(n2), .Z(_zy_simnet_cio_315[9]));
Q_BUF U1247 ( .A(n2), .Z(_zy_simnet_cio_315[8]));
Q_BUF U1248 ( .A(n2), .Z(_zy_simnet_cio_315[7]));
Q_BUF U1249 ( .A(n2), .Z(_zy_simnet_cio_315[6]));
Q_BUF U1250 ( .A(n2), .Z(_zy_simnet_cio_315[5]));
Q_BUF U1251 ( .A(n2), .Z(_zy_simnet_cio_315[4]));
Q_BUF U1252 ( .A(n2), .Z(_zy_simnet_cio_315[3]));
Q_BUF U1253 ( .A(n2), .Z(_zy_simnet_cio_315[2]));
Q_BUF U1254 ( .A(n2), .Z(_zy_simnet_cio_315[1]));
Q_BUF U1255 ( .A(n2), .Z(_zy_simnet_cio_315[0]));
Q_BUF U1256 ( .A(n2), .Z(_zy_simnet_cio_282[1]));
Q_BUF U1257 ( .A(n2), .Z(_zy_simnet_cio_282[0]));
Q_BUF U1258 ( .A(n2), .Z(_zy_simnet_cio_275[1]));
Q_BUF U1259 ( .A(n2), .Z(_zy_simnet_cio_275[0]));
Q_BUF U1260 ( .A(n2), .Z(_zy_simnet_cio_268[1]));
Q_BUF U1261 ( .A(n2), .Z(_zy_simnet_cio_268[0]));
Q_BUF U1262 ( .A(n2), .Z(_zy_simnet_cio_261[1]));
Q_BUF U1263 ( .A(n2), .Z(_zy_simnet_cio_261[0]));
Q_BUF U1264 ( .A(n2), .Z(_zy_simnet_cio_254[1]));
Q_BUF U1265 ( .A(n2), .Z(_zy_simnet_cio_254[0]));
Q_BUF U1266 ( .A(n2), .Z(_zy_simnet_cio_247[1]));
Q_BUF U1267 ( .A(n2), .Z(_zy_simnet_cio_247[0]));
Q_BUF U1268 ( .A(n2), .Z(_zy_simnet_cio_240[1]));
Q_BUF U1269 ( .A(n2), .Z(_zy_simnet_cio_240[0]));
Q_BUF U1270 ( .A(n2), .Z(_zy_simnet_cio_233[1]));
Q_BUF U1271 ( .A(n2), .Z(_zy_simnet_cio_233[0]));
Q_BUF U1272 ( .A(n2), .Z(_zy_simnet_cio_24));
Q_BUF U1273 ( .A(n2), .Z(blkid_revid_config[8]));
Q_BUF U1274 ( .A(n2), .Z(blkid_revid_config[9]));
Q_BUF U1275 ( .A(n2), .Z(blkid_revid_config[10]));
Q_BUF U1276 ( .A(n2), .Z(blkid_revid_config[11]));
Q_BUF U1277 ( .A(n2), .Z(blkid_revid_config[12]));
Q_BUF U1278 ( .A(n2), .Z(blkid_revid_config[13]));
Q_BUF U1279 ( .A(n2), .Z(blkid_revid_config[14]));
Q_BUF U1280 ( .A(n2), .Z(blkid_revid_config[15]));
Q_BUF U1281 ( .A(n2), .Z(blkid_revid_config[16]));
Q_BUF U1282 ( .A(n2), .Z(blkid_revid_config[17]));
Q_BUF U1283 ( .A(n2), .Z(blkid_revid_config[18]));
Q_BUF U1284 ( .A(n2), .Z(blkid_revid_config[19]));
Q_BUF U1285 ( .A(n2), .Z(blkid_revid_config[20]));
Q_BUF U1286 ( .A(n2), .Z(blkid_revid_config[21]));
Q_BUF U1287 ( .A(n2), .Z(blkid_revid_config[22]));
Q_BUF U1288 ( .A(n2), .Z(blkid_revid_config[23]));
Q_BUF U1289 ( .A(n1), .Z(blkid_revid_config[24]));
Q_BUF U1290 ( .A(n1), .Z(blkid_revid_config[25]));
Q_BUF U1291 ( .A(n1), .Z(blkid_revid_config[26]));
Q_BUF U1292 ( .A(n1), .Z(blkid_revid_config[27]));
Q_BUF U1293 ( .A(n2), .Z(blkid_revid_config[28]));
Q_BUF U1294 ( .A(n2), .Z(blkid_revid_config[29]));
Q_BUF U1295 ( .A(n1), .Z(blkid_revid_config[30]));
Q_BUF U1296 ( .A(n1), .Z(blkid_revid_config[31]));
Q_BUF U1297 ( .A(n2), .Z(cddip3_im_din[0]));
Q_BUF U1298 ( .A(n2), .Z(cddip3_im_din[1]));
Q_BUF U1299 ( .A(n2), .Z(cddip3_im_din[2]));
Q_BUF U1300 ( .A(n2), .Z(cddip3_im_din[3]));
Q_BUF U1301 ( .A(n2), .Z(cddip3_im_din[4]));
Q_BUF U1302 ( .A(n2), .Z(cddip3_im_din[5]));
Q_BUF U1303 ( .A(n2), .Z(cddip3_im_din[15]));
Q_BUF U1304 ( .A(n2), .Z(cddip3_im_din[16]));
Q_BUF U1305 ( .A(n2), .Z(cddip3_im_din[17]));
Q_BUF U1306 ( .A(n2), .Z(cddip3_im_din[18]));
Q_BUF U1307 ( .A(n2), .Z(cddip3_im_din[19]));
Q_BUF U1308 ( .A(n2), .Z(cddip3_im_din[20]));
Q_BUF U1309 ( .A(n2), .Z(cddip3_im_din[21]));
Q_BUF U1310 ( .A(n2), .Z(cddip3_im_din[22]));
Q_BUF U1311 ( .A(n2), .Z(cceip3_im_din[0]));
Q_BUF U1312 ( .A(n2), .Z(cceip3_im_din[1]));
Q_BUF U1313 ( .A(n2), .Z(cceip3_im_din[2]));
Q_BUF U1314 ( .A(n2), .Z(cceip3_im_din[3]));
Q_BUF U1315 ( .A(n2), .Z(cceip3_im_din[4]));
Q_BUF U1316 ( .A(n2), .Z(cceip3_im_din[5]));
Q_BUF U1317 ( .A(n2), .Z(cceip3_im_din[15]));
Q_BUF U1318 ( .A(n2), .Z(cceip3_im_din[16]));
Q_BUF U1319 ( .A(n2), .Z(cceip3_im_din[17]));
Q_BUF U1320 ( .A(n2), .Z(cceip3_im_din[18]));
Q_BUF U1321 ( .A(n2), .Z(cceip3_im_din[19]));
Q_BUF U1322 ( .A(n2), .Z(cceip3_im_din[20]));
Q_BUF U1323 ( .A(n2), .Z(cceip3_im_din[21]));
Q_BUF U1324 ( .A(n2), .Z(cceip3_im_din[22]));
Q_BUF U1325 ( .A(n2), .Z(cddip2_im_din[0]));
Q_BUF U1326 ( .A(n2), .Z(cddip2_im_din[1]));
Q_BUF U1327 ( .A(n2), .Z(cddip2_im_din[2]));
Q_BUF U1328 ( .A(n2), .Z(cddip2_im_din[3]));
Q_BUF U1329 ( .A(n2), .Z(cddip2_im_din[4]));
Q_BUF U1330 ( .A(n2), .Z(cddip2_im_din[5]));
Q_BUF U1331 ( .A(n2), .Z(cddip2_im_din[15]));
Q_BUF U1332 ( .A(n2), .Z(cddip2_im_din[16]));
Q_BUF U1333 ( .A(n2), .Z(cddip2_im_din[17]));
Q_BUF U1334 ( .A(n2), .Z(cddip2_im_din[18]));
Q_BUF U1335 ( .A(n2), .Z(cddip2_im_din[19]));
Q_BUF U1336 ( .A(n2), .Z(cddip2_im_din[20]));
Q_BUF U1337 ( .A(n2), .Z(cddip2_im_din[21]));
Q_BUF U1338 ( .A(n2), .Z(cddip2_im_din[22]));
Q_BUF U1339 ( .A(n2), .Z(cceip2_im_din[0]));
Q_BUF U1340 ( .A(n2), .Z(cceip2_im_din[1]));
Q_BUF U1341 ( .A(n2), .Z(cceip2_im_din[2]));
Q_BUF U1342 ( .A(n2), .Z(cceip2_im_din[3]));
Q_BUF U1343 ( .A(n2), .Z(cceip2_im_din[4]));
Q_BUF U1344 ( .A(n2), .Z(cceip2_im_din[5]));
Q_BUF U1345 ( .A(n2), .Z(cceip2_im_din[15]));
Q_BUF U1346 ( .A(n2), .Z(cceip2_im_din[16]));
Q_BUF U1347 ( .A(n2), .Z(cceip2_im_din[17]));
Q_BUF U1348 ( .A(n2), .Z(cceip2_im_din[18]));
Q_BUF U1349 ( .A(n2), .Z(cceip2_im_din[19]));
Q_BUF U1350 ( .A(n2), .Z(cceip2_im_din[20]));
Q_BUF U1351 ( .A(n2), .Z(cceip2_im_din[21]));
Q_BUF U1352 ( .A(n2), .Z(cceip2_im_din[22]));
Q_BUF U1353 ( .A(n2), .Z(cddip1_im_din[0]));
Q_BUF U1354 ( .A(n2), .Z(cddip1_im_din[1]));
Q_BUF U1355 ( .A(n2), .Z(cddip1_im_din[2]));
Q_BUF U1356 ( .A(n2), .Z(cddip1_im_din[3]));
Q_BUF U1357 ( .A(n2), .Z(cddip1_im_din[4]));
Q_BUF U1358 ( .A(n2), .Z(cddip1_im_din[5]));
Q_BUF U1359 ( .A(n2), .Z(cddip1_im_din[15]));
Q_BUF U1360 ( .A(n2), .Z(cddip1_im_din[16]));
Q_BUF U1361 ( .A(n2), .Z(cddip1_im_din[17]));
Q_BUF U1362 ( .A(n2), .Z(cddip1_im_din[18]));
Q_BUF U1363 ( .A(n2), .Z(cddip1_im_din[19]));
Q_BUF U1364 ( .A(n2), .Z(cddip1_im_din[20]));
Q_BUF U1365 ( .A(n2), .Z(cddip1_im_din[21]));
Q_BUF U1366 ( .A(n2), .Z(cddip1_im_din[22]));
Q_BUF U1367 ( .A(n2), .Z(cceip1_im_din[0]));
Q_BUF U1368 ( .A(n2), .Z(cceip1_im_din[1]));
Q_BUF U1369 ( .A(n2), .Z(cceip1_im_din[2]));
Q_BUF U1370 ( .A(n2), .Z(cceip1_im_din[3]));
Q_BUF U1371 ( .A(n2), .Z(cceip1_im_din[4]));
Q_BUF U1372 ( .A(n2), .Z(cceip1_im_din[5]));
Q_BUF U1373 ( .A(n2), .Z(cceip1_im_din[15]));
Q_BUF U1374 ( .A(n2), .Z(cceip1_im_din[16]));
Q_BUF U1375 ( .A(n2), .Z(cceip1_im_din[17]));
Q_BUF U1376 ( .A(n2), .Z(cceip1_im_din[18]));
Q_BUF U1377 ( .A(n2), .Z(cceip1_im_din[19]));
Q_BUF U1378 ( .A(n2), .Z(cceip1_im_din[20]));
Q_BUF U1379 ( .A(n2), .Z(cceip1_im_din[21]));
Q_BUF U1380 ( .A(n2), .Z(cceip1_im_din[22]));
Q_BUF U1381 ( .A(n2), .Z(cddip0_im_din[0]));
Q_BUF U1382 ( .A(n2), .Z(cddip0_im_din[1]));
Q_BUF U1383 ( .A(n2), .Z(cddip0_im_din[2]));
Q_BUF U1384 ( .A(n2), .Z(cddip0_im_din[3]));
Q_BUF U1385 ( .A(n2), .Z(cddip0_im_din[4]));
Q_BUF U1386 ( .A(n2), .Z(cddip0_im_din[5]));
Q_BUF U1387 ( .A(n2), .Z(cddip0_im_din[15]));
Q_BUF U1388 ( .A(n2), .Z(cddip0_im_din[16]));
Q_BUF U1389 ( .A(n2), .Z(cddip0_im_din[17]));
Q_BUF U1390 ( .A(n2), .Z(cddip0_im_din[18]));
Q_BUF U1391 ( .A(n2), .Z(cddip0_im_din[19]));
Q_BUF U1392 ( .A(n2), .Z(cddip0_im_din[20]));
Q_BUF U1393 ( .A(n2), .Z(cddip0_im_din[21]));
Q_BUF U1394 ( .A(n2), .Z(cddip0_im_din[22]));
Q_BUF U1395 ( .A(n2), .Z(cceip0_im_din[0]));
Q_BUF U1396 ( .A(n2), .Z(cceip0_im_din[1]));
Q_BUF U1397 ( .A(n2), .Z(cceip0_im_din[2]));
Q_BUF U1398 ( .A(n2), .Z(cceip0_im_din[3]));
Q_BUF U1399 ( .A(n2), .Z(cceip0_im_din[4]));
Q_BUF U1400 ( .A(n2), .Z(cceip0_im_din[5]));
Q_BUF U1401 ( .A(n2), .Z(cceip0_im_din[15]));
Q_BUF U1402 ( .A(n2), .Z(cceip0_im_din[16]));
Q_BUF U1403 ( .A(n2), .Z(cceip0_im_din[17]));
Q_BUF U1404 ( .A(n2), .Z(cceip0_im_din[18]));
Q_BUF U1405 ( .A(n2), .Z(cceip0_im_din[19]));
Q_BUF U1406 ( .A(n2), .Z(cceip0_im_din[20]));
Q_BUF U1407 ( .A(n2), .Z(cceip0_im_din[21]));
Q_BUF U1408 ( .A(n2), .Z(cceip0_im_din[22]));
Q_ASSIGN U1409 ( .B(im_available_kme_cceip0[0]), .A(im_available[0]));
Q_ASSIGN U1410 ( .B(im_available_kme_cceip0[1]), .A(im_available[1]));
Q_ASSIGN U1411 ( .B(im_available_kme_cceip1[0]), .A(im_available[2]));
Q_ASSIGN U1412 ( .B(im_available_kme_cceip1[1]), .A(im_available[3]));
Q_ASSIGN U1413 ( .B(im_available_kme_cceip2[0]), .A(im_available[4]));
Q_ASSIGN U1414 ( .B(im_available_kme_cceip2[1]), .A(im_available[5]));
Q_ASSIGN U1415 ( .B(im_available_kme_cceip3[0]), .A(im_available[6]));
Q_ASSIGN U1416 ( .B(im_available_kme_cceip3[1]), .A(im_available[7]));
Q_ASSIGN U1417 ( .B(im_available_kme_cddip0[0]), .A(im_available[8]));
Q_ASSIGN U1418 ( .B(im_available_kme_cddip0[1]), .A(im_available[9]));
Q_ASSIGN U1419 ( .B(im_available_kme_cddip1[0]), .A(im_available[10]));
Q_ASSIGN U1420 ( .B(im_available_kme_cddip1[1]), .A(im_available[11]));
Q_ASSIGN U1421 ( .B(im_available_kme_cddip2[0]), .A(im_available[12]));
Q_ASSIGN U1422 ( .B(im_available_kme_cddip2[1]), .A(im_available[13]));
Q_ASSIGN U1423 ( .B(im_available_kme_cddip3[0]), .A(im_available[14]));
Q_ASSIGN U1424 ( .B(im_available_kme_cddip3[1]), .A(im_available[15]));
Q_ASSIGN U1425 ( .B(revid_wire[0]), .A(blkid_revid_config[0]));
Q_ASSIGN U1426 ( .B(revid_wire[1]), .A(blkid_revid_config[1]));
Q_ASSIGN U1427 ( .B(revid_wire[2]), .A(blkid_revid_config[2]));
Q_ASSIGN U1428 ( .B(revid_wire[3]), .A(blkid_revid_config[3]));
Q_ASSIGN U1429 ( .B(revid_wire[4]), .A(blkid_revid_config[4]));
Q_ASSIGN U1430 ( .B(revid_wire[5]), .A(blkid_revid_config[5]));
Q_ASSIGN U1431 ( .B(revid_wire[6]), .A(blkid_revid_config[6]));
Q_ASSIGN U1432 ( .B(revid_wire[7]), .A(blkid_revid_config[7]));
Q_ASSIGN U1433 ( .B(kme_cddip3_ob_out_pre[64]), .A(cddip3_im_din[6]));
Q_ASSIGN U1434 ( .B(kme_cddip3_ob_out_pre[66]), .A(cddip3_im_din[8]));
Q_ASSIGN U1435 ( .B(kme_cddip3_ob_out_pre[67]), .A(cddip3_im_din[9]));
Q_ASSIGN U1436 ( .B(kme_cddip3_ob_out_pre[68]), .A(cddip3_im_din[10]));
Q_ASSIGN U1437 ( .B(kme_cddip3_ob_out_pre[69]), .A(cddip3_im_din[11]));
Q_ASSIGN U1438 ( .B(kme_cddip3_ob_out_pre[70]), .A(cddip3_im_din[12]));
Q_ASSIGN U1439 ( .B(kme_cddip3_ob_out_pre[71]), .A(cddip3_im_din[13]));
Q_ASSIGN U1440 ( .B(kme_cddip3_ob_out_pre[80]), .A(cddip3_im_din[14]));
Q_ASSIGN U1441 ( .B(kme_cddip3_ob_out_pre[72]), .A(cddip3_im_din[23]));
Q_ASSIGN U1442 ( .B(kme_cddip3_ob_out_pre[73]), .A(cddip3_im_din[24]));
Q_ASSIGN U1443 ( .B(kme_cddip3_ob_out_pre[74]), .A(cddip3_im_din[25]));
Q_ASSIGN U1444 ( .B(kme_cddip3_ob_out_pre[75]), .A(cddip3_im_din[26]));
Q_ASSIGN U1445 ( .B(kme_cddip3_ob_out_pre[76]), .A(cddip3_im_din[27]));
Q_ASSIGN U1446 ( .B(kme_cddip3_ob_out_pre[77]), .A(cddip3_im_din[28]));
Q_ASSIGN U1447 ( .B(kme_cddip3_ob_out_pre[78]), .A(cddip3_im_din[29]));
Q_ASSIGN U1448 ( .B(kme_cddip3_ob_out_pre[79]), .A(cddip3_im_din[30]));
Q_ASSIGN U1449 ( .B(kme_cddip3_ob_out_pre[65]), .A(cddip3_im_din[31]));
Q_ASSIGN U1450 ( .B(kme_cddip3_ob_out_pre[65]), .A(cddip3_im_din[7]));
Q_ASSIGN U1451 ( .B(kme_cddip3_ob_out_pre[0]), .A(cddip3_im_din[32]));
Q_ASSIGN U1452 ( .B(kme_cddip3_ob_out_pre[1]), .A(cddip3_im_din[33]));
Q_ASSIGN U1453 ( .B(kme_cddip3_ob_out_pre[2]), .A(cddip3_im_din[34]));
Q_ASSIGN U1454 ( .B(kme_cddip3_ob_out_pre[3]), .A(cddip3_im_din[35]));
Q_ASSIGN U1455 ( .B(kme_cddip3_ob_out_pre[4]), .A(cddip3_im_din[36]));
Q_ASSIGN U1456 ( .B(kme_cddip3_ob_out_pre[5]), .A(cddip3_im_din[37]));
Q_ASSIGN U1457 ( .B(kme_cddip3_ob_out_pre[6]), .A(cddip3_im_din[38]));
Q_ASSIGN U1458 ( .B(kme_cddip3_ob_out_pre[7]), .A(cddip3_im_din[39]));
Q_ASSIGN U1459 ( .B(kme_cddip3_ob_out_pre[8]), .A(cddip3_im_din[40]));
Q_ASSIGN U1460 ( .B(kme_cddip3_ob_out_pre[9]), .A(cddip3_im_din[41]));
Q_ASSIGN U1461 ( .B(kme_cddip3_ob_out_pre[10]), .A(cddip3_im_din[42]));
Q_ASSIGN U1462 ( .B(kme_cddip3_ob_out_pre[11]), .A(cddip3_im_din[43]));
Q_ASSIGN U1463 ( .B(kme_cddip3_ob_out_pre[12]), .A(cddip3_im_din[44]));
Q_ASSIGN U1464 ( .B(kme_cddip3_ob_out_pre[13]), .A(cddip3_im_din[45]));
Q_ASSIGN U1465 ( .B(kme_cddip3_ob_out_pre[14]), .A(cddip3_im_din[46]));
Q_ASSIGN U1466 ( .B(kme_cddip3_ob_out_pre[15]), .A(cddip3_im_din[47]));
Q_ASSIGN U1467 ( .B(kme_cddip3_ob_out_pre[16]), .A(cddip3_im_din[48]));
Q_ASSIGN U1468 ( .B(kme_cddip3_ob_out_pre[17]), .A(cddip3_im_din[49]));
Q_ASSIGN U1469 ( .B(kme_cddip3_ob_out_pre[18]), .A(cddip3_im_din[50]));
Q_ASSIGN U1470 ( .B(kme_cddip3_ob_out_pre[19]), .A(cddip3_im_din[51]));
Q_ASSIGN U1471 ( .B(kme_cddip3_ob_out_pre[20]), .A(cddip3_im_din[52]));
Q_ASSIGN U1472 ( .B(kme_cddip3_ob_out_pre[21]), .A(cddip3_im_din[53]));
Q_ASSIGN U1473 ( .B(kme_cddip3_ob_out_pre[22]), .A(cddip3_im_din[54]));
Q_ASSIGN U1474 ( .B(kme_cddip3_ob_out_pre[23]), .A(cddip3_im_din[55]));
Q_ASSIGN U1475 ( .B(kme_cddip3_ob_out_pre[24]), .A(cddip3_im_din[56]));
Q_ASSIGN U1476 ( .B(kme_cddip3_ob_out_pre[25]), .A(cddip3_im_din[57]));
Q_ASSIGN U1477 ( .B(kme_cddip3_ob_out_pre[26]), .A(cddip3_im_din[58]));
Q_ASSIGN U1478 ( .B(kme_cddip3_ob_out_pre[27]), .A(cddip3_im_din[59]));
Q_ASSIGN U1479 ( .B(kme_cddip3_ob_out_pre[28]), .A(cddip3_im_din[60]));
Q_ASSIGN U1480 ( .B(kme_cddip3_ob_out_pre[29]), .A(cddip3_im_din[61]));
Q_ASSIGN U1481 ( .B(kme_cddip3_ob_out_pre[30]), .A(cddip3_im_din[62]));
Q_ASSIGN U1482 ( .B(kme_cddip3_ob_out_pre[31]), .A(cddip3_im_din[63]));
Q_ASSIGN U1483 ( .B(kme_cddip3_ob_out_pre[32]), .A(cddip3_im_din[64]));
Q_ASSIGN U1484 ( .B(kme_cddip3_ob_out_pre[33]), .A(cddip3_im_din[65]));
Q_ASSIGN U1485 ( .B(kme_cddip3_ob_out_pre[34]), .A(cddip3_im_din[66]));
Q_ASSIGN U1486 ( .B(kme_cddip3_ob_out_pre[35]), .A(cddip3_im_din[67]));
Q_ASSIGN U1487 ( .B(kme_cddip3_ob_out_pre[36]), .A(cddip3_im_din[68]));
Q_ASSIGN U1488 ( .B(kme_cddip3_ob_out_pre[37]), .A(cddip3_im_din[69]));
Q_ASSIGN U1489 ( .B(kme_cddip3_ob_out_pre[38]), .A(cddip3_im_din[70]));
Q_ASSIGN U1490 ( .B(kme_cddip3_ob_out_pre[39]), .A(cddip3_im_din[71]));
Q_ASSIGN U1491 ( .B(kme_cddip3_ob_out_pre[40]), .A(cddip3_im_din[72]));
Q_ASSIGN U1492 ( .B(kme_cddip3_ob_out_pre[41]), .A(cddip3_im_din[73]));
Q_ASSIGN U1493 ( .B(kme_cddip3_ob_out_pre[42]), .A(cddip3_im_din[74]));
Q_ASSIGN U1494 ( .B(kme_cddip3_ob_out_pre[43]), .A(cddip3_im_din[75]));
Q_ASSIGN U1495 ( .B(kme_cddip3_ob_out_pre[44]), .A(cddip3_im_din[76]));
Q_ASSIGN U1496 ( .B(kme_cddip3_ob_out_pre[45]), .A(cddip3_im_din[77]));
Q_ASSIGN U1497 ( .B(kme_cddip3_ob_out_pre[46]), .A(cddip3_im_din[78]));
Q_ASSIGN U1498 ( .B(kme_cddip3_ob_out_pre[47]), .A(cddip3_im_din[79]));
Q_ASSIGN U1499 ( .B(kme_cddip3_ob_out_pre[48]), .A(cddip3_im_din[80]));
Q_ASSIGN U1500 ( .B(kme_cddip3_ob_out_pre[49]), .A(cddip3_im_din[81]));
Q_ASSIGN U1501 ( .B(kme_cddip3_ob_out_pre[50]), .A(cddip3_im_din[82]));
Q_ASSIGN U1502 ( .B(kme_cddip3_ob_out_pre[51]), .A(cddip3_im_din[83]));
Q_ASSIGN U1503 ( .B(kme_cddip3_ob_out_pre[52]), .A(cddip3_im_din[84]));
Q_ASSIGN U1504 ( .B(kme_cddip3_ob_out_pre[53]), .A(cddip3_im_din[85]));
Q_ASSIGN U1505 ( .B(kme_cddip3_ob_out_pre[54]), .A(cddip3_im_din[86]));
Q_ASSIGN U1506 ( .B(kme_cddip3_ob_out_pre[55]), .A(cddip3_im_din[87]));
Q_ASSIGN U1507 ( .B(kme_cddip3_ob_out_pre[56]), .A(cddip3_im_din[88]));
Q_ASSIGN U1508 ( .B(kme_cddip3_ob_out_pre[57]), .A(cddip3_im_din[89]));
Q_ASSIGN U1509 ( .B(kme_cddip3_ob_out_pre[58]), .A(cddip3_im_din[90]));
Q_ASSIGN U1510 ( .B(kme_cddip3_ob_out_pre[59]), .A(cddip3_im_din[91]));
Q_ASSIGN U1511 ( .B(kme_cddip3_ob_out_pre[60]), .A(cddip3_im_din[92]));
Q_ASSIGN U1512 ( .B(kme_cddip3_ob_out_pre[61]), .A(cddip3_im_din[93]));
Q_ASSIGN U1513 ( .B(kme_cddip3_ob_out_pre[62]), .A(cddip3_im_din[94]));
Q_ASSIGN U1514 ( .B(kme_cddip3_ob_out_pre[63]), .A(cddip3_im_din[95]));
Q_ASSIGN U1515 ( .B(kme_cceip3_ob_out_pre[64]), .A(cceip3_im_din[6]));
Q_ASSIGN U1516 ( .B(kme_cceip3_ob_out_pre[66]), .A(cceip3_im_din[8]));
Q_ASSIGN U1517 ( .B(kme_cceip3_ob_out_pre[67]), .A(cceip3_im_din[9]));
Q_ASSIGN U1518 ( .B(kme_cceip3_ob_out_pre[68]), .A(cceip3_im_din[10]));
Q_ASSIGN U1519 ( .B(kme_cceip3_ob_out_pre[69]), .A(cceip3_im_din[11]));
Q_ASSIGN U1520 ( .B(kme_cceip3_ob_out_pre[70]), .A(cceip3_im_din[12]));
Q_ASSIGN U1521 ( .B(kme_cceip3_ob_out_pre[71]), .A(cceip3_im_din[13]));
Q_ASSIGN U1522 ( .B(kme_cceip3_ob_out_pre[80]), .A(cceip3_im_din[14]));
Q_ASSIGN U1523 ( .B(kme_cceip3_ob_out_pre[72]), .A(cceip3_im_din[23]));
Q_ASSIGN U1524 ( .B(kme_cceip3_ob_out_pre[73]), .A(cceip3_im_din[24]));
Q_ASSIGN U1525 ( .B(kme_cceip3_ob_out_pre[74]), .A(cceip3_im_din[25]));
Q_ASSIGN U1526 ( .B(kme_cceip3_ob_out_pre[75]), .A(cceip3_im_din[26]));
Q_ASSIGN U1527 ( .B(kme_cceip3_ob_out_pre[76]), .A(cceip3_im_din[27]));
Q_ASSIGN U1528 ( .B(kme_cceip3_ob_out_pre[77]), .A(cceip3_im_din[28]));
Q_ASSIGN U1529 ( .B(kme_cceip3_ob_out_pre[78]), .A(cceip3_im_din[29]));
Q_ASSIGN U1530 ( .B(kme_cceip3_ob_out_pre[79]), .A(cceip3_im_din[30]));
Q_ASSIGN U1531 ( .B(kme_cceip3_ob_out_pre[65]), .A(cceip3_im_din[31]));
Q_ASSIGN U1532 ( .B(kme_cceip3_ob_out_pre[65]), .A(cceip3_im_din[7]));
Q_ASSIGN U1533 ( .B(kme_cceip3_ob_out_pre[0]), .A(cceip3_im_din[32]));
Q_ASSIGN U1534 ( .B(kme_cceip3_ob_out_pre[1]), .A(cceip3_im_din[33]));
Q_ASSIGN U1535 ( .B(kme_cceip3_ob_out_pre[2]), .A(cceip3_im_din[34]));
Q_ASSIGN U1536 ( .B(kme_cceip3_ob_out_pre[3]), .A(cceip3_im_din[35]));
Q_ASSIGN U1537 ( .B(kme_cceip3_ob_out_pre[4]), .A(cceip3_im_din[36]));
Q_ASSIGN U1538 ( .B(kme_cceip3_ob_out_pre[5]), .A(cceip3_im_din[37]));
Q_ASSIGN U1539 ( .B(kme_cceip3_ob_out_pre[6]), .A(cceip3_im_din[38]));
Q_ASSIGN U1540 ( .B(kme_cceip3_ob_out_pre[7]), .A(cceip3_im_din[39]));
Q_ASSIGN U1541 ( .B(kme_cceip3_ob_out_pre[8]), .A(cceip3_im_din[40]));
Q_ASSIGN U1542 ( .B(kme_cceip3_ob_out_pre[9]), .A(cceip3_im_din[41]));
Q_ASSIGN U1543 ( .B(kme_cceip3_ob_out_pre[10]), .A(cceip3_im_din[42]));
Q_ASSIGN U1544 ( .B(kme_cceip3_ob_out_pre[11]), .A(cceip3_im_din[43]));
Q_ASSIGN U1545 ( .B(kme_cceip3_ob_out_pre[12]), .A(cceip3_im_din[44]));
Q_ASSIGN U1546 ( .B(kme_cceip3_ob_out_pre[13]), .A(cceip3_im_din[45]));
Q_ASSIGN U1547 ( .B(kme_cceip3_ob_out_pre[14]), .A(cceip3_im_din[46]));
Q_ASSIGN U1548 ( .B(kme_cceip3_ob_out_pre[15]), .A(cceip3_im_din[47]));
Q_ASSIGN U1549 ( .B(kme_cceip3_ob_out_pre[16]), .A(cceip3_im_din[48]));
Q_ASSIGN U1550 ( .B(kme_cceip3_ob_out_pre[17]), .A(cceip3_im_din[49]));
Q_ASSIGN U1551 ( .B(kme_cceip3_ob_out_pre[18]), .A(cceip3_im_din[50]));
Q_ASSIGN U1552 ( .B(kme_cceip3_ob_out_pre[19]), .A(cceip3_im_din[51]));
Q_ASSIGN U1553 ( .B(kme_cceip3_ob_out_pre[20]), .A(cceip3_im_din[52]));
Q_ASSIGN U1554 ( .B(kme_cceip3_ob_out_pre[21]), .A(cceip3_im_din[53]));
Q_ASSIGN U1555 ( .B(kme_cceip3_ob_out_pre[22]), .A(cceip3_im_din[54]));
Q_ASSIGN U1556 ( .B(kme_cceip3_ob_out_pre[23]), .A(cceip3_im_din[55]));
Q_ASSIGN U1557 ( .B(kme_cceip3_ob_out_pre[24]), .A(cceip3_im_din[56]));
Q_ASSIGN U1558 ( .B(kme_cceip3_ob_out_pre[25]), .A(cceip3_im_din[57]));
Q_ASSIGN U1559 ( .B(kme_cceip3_ob_out_pre[26]), .A(cceip3_im_din[58]));
Q_ASSIGN U1560 ( .B(kme_cceip3_ob_out_pre[27]), .A(cceip3_im_din[59]));
Q_ASSIGN U1561 ( .B(kme_cceip3_ob_out_pre[28]), .A(cceip3_im_din[60]));
Q_ASSIGN U1562 ( .B(kme_cceip3_ob_out_pre[29]), .A(cceip3_im_din[61]));
Q_ASSIGN U1563 ( .B(kme_cceip3_ob_out_pre[30]), .A(cceip3_im_din[62]));
Q_ASSIGN U1564 ( .B(kme_cceip3_ob_out_pre[31]), .A(cceip3_im_din[63]));
Q_ASSIGN U1565 ( .B(kme_cceip3_ob_out_pre[32]), .A(cceip3_im_din[64]));
Q_ASSIGN U1566 ( .B(kme_cceip3_ob_out_pre[33]), .A(cceip3_im_din[65]));
Q_ASSIGN U1567 ( .B(kme_cceip3_ob_out_pre[34]), .A(cceip3_im_din[66]));
Q_ASSIGN U1568 ( .B(kme_cceip3_ob_out_pre[35]), .A(cceip3_im_din[67]));
Q_ASSIGN U1569 ( .B(kme_cceip3_ob_out_pre[36]), .A(cceip3_im_din[68]));
Q_ASSIGN U1570 ( .B(kme_cceip3_ob_out_pre[37]), .A(cceip3_im_din[69]));
Q_ASSIGN U1571 ( .B(kme_cceip3_ob_out_pre[38]), .A(cceip3_im_din[70]));
Q_ASSIGN U1572 ( .B(kme_cceip3_ob_out_pre[39]), .A(cceip3_im_din[71]));
Q_ASSIGN U1573 ( .B(kme_cceip3_ob_out_pre[40]), .A(cceip3_im_din[72]));
Q_ASSIGN U1574 ( .B(kme_cceip3_ob_out_pre[41]), .A(cceip3_im_din[73]));
Q_ASSIGN U1575 ( .B(kme_cceip3_ob_out_pre[42]), .A(cceip3_im_din[74]));
Q_ASSIGN U1576 ( .B(kme_cceip3_ob_out_pre[43]), .A(cceip3_im_din[75]));
Q_ASSIGN U1577 ( .B(kme_cceip3_ob_out_pre[44]), .A(cceip3_im_din[76]));
Q_ASSIGN U1578 ( .B(kme_cceip3_ob_out_pre[45]), .A(cceip3_im_din[77]));
Q_ASSIGN U1579 ( .B(kme_cceip3_ob_out_pre[46]), .A(cceip3_im_din[78]));
Q_ASSIGN U1580 ( .B(kme_cceip3_ob_out_pre[47]), .A(cceip3_im_din[79]));
Q_ASSIGN U1581 ( .B(kme_cceip3_ob_out_pre[48]), .A(cceip3_im_din[80]));
Q_ASSIGN U1582 ( .B(kme_cceip3_ob_out_pre[49]), .A(cceip3_im_din[81]));
Q_ASSIGN U1583 ( .B(kme_cceip3_ob_out_pre[50]), .A(cceip3_im_din[82]));
Q_ASSIGN U1584 ( .B(kme_cceip3_ob_out_pre[51]), .A(cceip3_im_din[83]));
Q_ASSIGN U1585 ( .B(kme_cceip3_ob_out_pre[52]), .A(cceip3_im_din[84]));
Q_ASSIGN U1586 ( .B(kme_cceip3_ob_out_pre[53]), .A(cceip3_im_din[85]));
Q_ASSIGN U1587 ( .B(kme_cceip3_ob_out_pre[54]), .A(cceip3_im_din[86]));
Q_ASSIGN U1588 ( .B(kme_cceip3_ob_out_pre[55]), .A(cceip3_im_din[87]));
Q_ASSIGN U1589 ( .B(kme_cceip3_ob_out_pre[56]), .A(cceip3_im_din[88]));
Q_ASSIGN U1590 ( .B(kme_cceip3_ob_out_pre[57]), .A(cceip3_im_din[89]));
Q_ASSIGN U1591 ( .B(kme_cceip3_ob_out_pre[58]), .A(cceip3_im_din[90]));
Q_ASSIGN U1592 ( .B(kme_cceip3_ob_out_pre[59]), .A(cceip3_im_din[91]));
Q_ASSIGN U1593 ( .B(kme_cceip3_ob_out_pre[60]), .A(cceip3_im_din[92]));
Q_ASSIGN U1594 ( .B(kme_cceip3_ob_out_pre[61]), .A(cceip3_im_din[93]));
Q_ASSIGN U1595 ( .B(kme_cceip3_ob_out_pre[62]), .A(cceip3_im_din[94]));
Q_ASSIGN U1596 ( .B(kme_cceip3_ob_out_pre[63]), .A(cceip3_im_din[95]));
Q_ASSIGN U1597 ( .B(kme_cddip2_ob_out_pre[64]), .A(cddip2_im_din[6]));
Q_ASSIGN U1598 ( .B(kme_cddip2_ob_out_pre[66]), .A(cddip2_im_din[8]));
Q_ASSIGN U1599 ( .B(kme_cddip2_ob_out_pre[67]), .A(cddip2_im_din[9]));
Q_ASSIGN U1600 ( .B(kme_cddip2_ob_out_pre[68]), .A(cddip2_im_din[10]));
Q_ASSIGN U1601 ( .B(kme_cddip2_ob_out_pre[69]), .A(cddip2_im_din[11]));
Q_ASSIGN U1602 ( .B(kme_cddip2_ob_out_pre[70]), .A(cddip2_im_din[12]));
Q_ASSIGN U1603 ( .B(kme_cddip2_ob_out_pre[71]), .A(cddip2_im_din[13]));
Q_ASSIGN U1604 ( .B(kme_cddip2_ob_out_pre[80]), .A(cddip2_im_din[14]));
Q_ASSIGN U1605 ( .B(kme_cddip2_ob_out_pre[72]), .A(cddip2_im_din[23]));
Q_ASSIGN U1606 ( .B(kme_cddip2_ob_out_pre[73]), .A(cddip2_im_din[24]));
Q_ASSIGN U1607 ( .B(kme_cddip2_ob_out_pre[74]), .A(cddip2_im_din[25]));
Q_ASSIGN U1608 ( .B(kme_cddip2_ob_out_pre[75]), .A(cddip2_im_din[26]));
Q_ASSIGN U1609 ( .B(kme_cddip2_ob_out_pre[76]), .A(cddip2_im_din[27]));
Q_ASSIGN U1610 ( .B(kme_cddip2_ob_out_pre[77]), .A(cddip2_im_din[28]));
Q_ASSIGN U1611 ( .B(kme_cddip2_ob_out_pre[78]), .A(cddip2_im_din[29]));
Q_ASSIGN U1612 ( .B(kme_cddip2_ob_out_pre[79]), .A(cddip2_im_din[30]));
Q_ASSIGN U1613 ( .B(kme_cddip2_ob_out_pre[65]), .A(cddip2_im_din[31]));
Q_ASSIGN U1614 ( .B(kme_cddip2_ob_out_pre[65]), .A(cddip2_im_din[7]));
Q_ASSIGN U1615 ( .B(kme_cddip2_ob_out_pre[0]), .A(cddip2_im_din[32]));
Q_ASSIGN U1616 ( .B(kme_cddip2_ob_out_pre[1]), .A(cddip2_im_din[33]));
Q_ASSIGN U1617 ( .B(kme_cddip2_ob_out_pre[2]), .A(cddip2_im_din[34]));
Q_ASSIGN U1618 ( .B(kme_cddip2_ob_out_pre[3]), .A(cddip2_im_din[35]));
Q_ASSIGN U1619 ( .B(kme_cddip2_ob_out_pre[4]), .A(cddip2_im_din[36]));
Q_ASSIGN U1620 ( .B(kme_cddip2_ob_out_pre[5]), .A(cddip2_im_din[37]));
Q_ASSIGN U1621 ( .B(kme_cddip2_ob_out_pre[6]), .A(cddip2_im_din[38]));
Q_ASSIGN U1622 ( .B(kme_cddip2_ob_out_pre[7]), .A(cddip2_im_din[39]));
Q_ASSIGN U1623 ( .B(kme_cddip2_ob_out_pre[8]), .A(cddip2_im_din[40]));
Q_ASSIGN U1624 ( .B(kme_cddip2_ob_out_pre[9]), .A(cddip2_im_din[41]));
Q_ASSIGN U1625 ( .B(kme_cddip2_ob_out_pre[10]), .A(cddip2_im_din[42]));
Q_ASSIGN U1626 ( .B(kme_cddip2_ob_out_pre[11]), .A(cddip2_im_din[43]));
Q_ASSIGN U1627 ( .B(kme_cddip2_ob_out_pre[12]), .A(cddip2_im_din[44]));
Q_ASSIGN U1628 ( .B(kme_cddip2_ob_out_pre[13]), .A(cddip2_im_din[45]));
Q_ASSIGN U1629 ( .B(kme_cddip2_ob_out_pre[14]), .A(cddip2_im_din[46]));
Q_ASSIGN U1630 ( .B(kme_cddip2_ob_out_pre[15]), .A(cddip2_im_din[47]));
Q_ASSIGN U1631 ( .B(kme_cddip2_ob_out_pre[16]), .A(cddip2_im_din[48]));
Q_ASSIGN U1632 ( .B(kme_cddip2_ob_out_pre[17]), .A(cddip2_im_din[49]));
Q_ASSIGN U1633 ( .B(kme_cddip2_ob_out_pre[18]), .A(cddip2_im_din[50]));
Q_ASSIGN U1634 ( .B(kme_cddip2_ob_out_pre[19]), .A(cddip2_im_din[51]));
Q_ASSIGN U1635 ( .B(kme_cddip2_ob_out_pre[20]), .A(cddip2_im_din[52]));
Q_ASSIGN U1636 ( .B(kme_cddip2_ob_out_pre[21]), .A(cddip2_im_din[53]));
Q_ASSIGN U1637 ( .B(kme_cddip2_ob_out_pre[22]), .A(cddip2_im_din[54]));
Q_ASSIGN U1638 ( .B(kme_cddip2_ob_out_pre[23]), .A(cddip2_im_din[55]));
Q_ASSIGN U1639 ( .B(kme_cddip2_ob_out_pre[24]), .A(cddip2_im_din[56]));
Q_ASSIGN U1640 ( .B(kme_cddip2_ob_out_pre[25]), .A(cddip2_im_din[57]));
Q_ASSIGN U1641 ( .B(kme_cddip2_ob_out_pre[26]), .A(cddip2_im_din[58]));
Q_ASSIGN U1642 ( .B(kme_cddip2_ob_out_pre[27]), .A(cddip2_im_din[59]));
Q_ASSIGN U1643 ( .B(kme_cddip2_ob_out_pre[28]), .A(cddip2_im_din[60]));
Q_ASSIGN U1644 ( .B(kme_cddip2_ob_out_pre[29]), .A(cddip2_im_din[61]));
Q_ASSIGN U1645 ( .B(kme_cddip2_ob_out_pre[30]), .A(cddip2_im_din[62]));
Q_ASSIGN U1646 ( .B(kme_cddip2_ob_out_pre[31]), .A(cddip2_im_din[63]));
Q_ASSIGN U1647 ( .B(kme_cddip2_ob_out_pre[32]), .A(cddip2_im_din[64]));
Q_ASSIGN U1648 ( .B(kme_cddip2_ob_out_pre[33]), .A(cddip2_im_din[65]));
Q_ASSIGN U1649 ( .B(kme_cddip2_ob_out_pre[34]), .A(cddip2_im_din[66]));
Q_ASSIGN U1650 ( .B(kme_cddip2_ob_out_pre[35]), .A(cddip2_im_din[67]));
Q_ASSIGN U1651 ( .B(kme_cddip2_ob_out_pre[36]), .A(cddip2_im_din[68]));
Q_ASSIGN U1652 ( .B(kme_cddip2_ob_out_pre[37]), .A(cddip2_im_din[69]));
Q_ASSIGN U1653 ( .B(kme_cddip2_ob_out_pre[38]), .A(cddip2_im_din[70]));
Q_ASSIGN U1654 ( .B(kme_cddip2_ob_out_pre[39]), .A(cddip2_im_din[71]));
Q_ASSIGN U1655 ( .B(kme_cddip2_ob_out_pre[40]), .A(cddip2_im_din[72]));
Q_ASSIGN U1656 ( .B(kme_cddip2_ob_out_pre[41]), .A(cddip2_im_din[73]));
Q_ASSIGN U1657 ( .B(kme_cddip2_ob_out_pre[42]), .A(cddip2_im_din[74]));
Q_ASSIGN U1658 ( .B(kme_cddip2_ob_out_pre[43]), .A(cddip2_im_din[75]));
Q_ASSIGN U1659 ( .B(kme_cddip2_ob_out_pre[44]), .A(cddip2_im_din[76]));
Q_ASSIGN U1660 ( .B(kme_cddip2_ob_out_pre[45]), .A(cddip2_im_din[77]));
Q_ASSIGN U1661 ( .B(kme_cddip2_ob_out_pre[46]), .A(cddip2_im_din[78]));
Q_ASSIGN U1662 ( .B(kme_cddip2_ob_out_pre[47]), .A(cddip2_im_din[79]));
Q_ASSIGN U1663 ( .B(kme_cddip2_ob_out_pre[48]), .A(cddip2_im_din[80]));
Q_ASSIGN U1664 ( .B(kme_cddip2_ob_out_pre[49]), .A(cddip2_im_din[81]));
Q_ASSIGN U1665 ( .B(kme_cddip2_ob_out_pre[50]), .A(cddip2_im_din[82]));
Q_ASSIGN U1666 ( .B(kme_cddip2_ob_out_pre[51]), .A(cddip2_im_din[83]));
Q_ASSIGN U1667 ( .B(kme_cddip2_ob_out_pre[52]), .A(cddip2_im_din[84]));
Q_ASSIGN U1668 ( .B(kme_cddip2_ob_out_pre[53]), .A(cddip2_im_din[85]));
Q_ASSIGN U1669 ( .B(kme_cddip2_ob_out_pre[54]), .A(cddip2_im_din[86]));
Q_ASSIGN U1670 ( .B(kme_cddip2_ob_out_pre[55]), .A(cddip2_im_din[87]));
Q_ASSIGN U1671 ( .B(kme_cddip2_ob_out_pre[56]), .A(cddip2_im_din[88]));
Q_ASSIGN U1672 ( .B(kme_cddip2_ob_out_pre[57]), .A(cddip2_im_din[89]));
Q_ASSIGN U1673 ( .B(kme_cddip2_ob_out_pre[58]), .A(cddip2_im_din[90]));
Q_ASSIGN U1674 ( .B(kme_cddip2_ob_out_pre[59]), .A(cddip2_im_din[91]));
Q_ASSIGN U1675 ( .B(kme_cddip2_ob_out_pre[60]), .A(cddip2_im_din[92]));
Q_ASSIGN U1676 ( .B(kme_cddip2_ob_out_pre[61]), .A(cddip2_im_din[93]));
Q_ASSIGN U1677 ( .B(kme_cddip2_ob_out_pre[62]), .A(cddip2_im_din[94]));
Q_ASSIGN U1678 ( .B(kme_cddip2_ob_out_pre[63]), .A(cddip2_im_din[95]));
Q_ASSIGN U1679 ( .B(kme_cceip2_ob_out_pre[64]), .A(cceip2_im_din[6]));
Q_ASSIGN U1680 ( .B(kme_cceip2_ob_out_pre[66]), .A(cceip2_im_din[8]));
Q_ASSIGN U1681 ( .B(kme_cceip2_ob_out_pre[67]), .A(cceip2_im_din[9]));
Q_ASSIGN U1682 ( .B(kme_cceip2_ob_out_pre[68]), .A(cceip2_im_din[10]));
Q_ASSIGN U1683 ( .B(kme_cceip2_ob_out_pre[69]), .A(cceip2_im_din[11]));
Q_ASSIGN U1684 ( .B(kme_cceip2_ob_out_pre[70]), .A(cceip2_im_din[12]));
Q_ASSIGN U1685 ( .B(kme_cceip2_ob_out_pre[71]), .A(cceip2_im_din[13]));
Q_ASSIGN U1686 ( .B(kme_cceip2_ob_out_pre[80]), .A(cceip2_im_din[14]));
Q_ASSIGN U1687 ( .B(kme_cceip2_ob_out_pre[72]), .A(cceip2_im_din[23]));
Q_ASSIGN U1688 ( .B(kme_cceip2_ob_out_pre[73]), .A(cceip2_im_din[24]));
Q_ASSIGN U1689 ( .B(kme_cceip2_ob_out_pre[74]), .A(cceip2_im_din[25]));
Q_ASSIGN U1690 ( .B(kme_cceip2_ob_out_pre[75]), .A(cceip2_im_din[26]));
Q_ASSIGN U1691 ( .B(kme_cceip2_ob_out_pre[76]), .A(cceip2_im_din[27]));
Q_ASSIGN U1692 ( .B(kme_cceip2_ob_out_pre[77]), .A(cceip2_im_din[28]));
Q_ASSIGN U1693 ( .B(kme_cceip2_ob_out_pre[78]), .A(cceip2_im_din[29]));
Q_ASSIGN U1694 ( .B(kme_cceip2_ob_out_pre[79]), .A(cceip2_im_din[30]));
Q_ASSIGN U1695 ( .B(kme_cceip2_ob_out_pre[65]), .A(cceip2_im_din[31]));
Q_ASSIGN U1696 ( .B(kme_cceip2_ob_out_pre[65]), .A(cceip2_im_din[7]));
Q_ASSIGN U1697 ( .B(kme_cceip2_ob_out_pre[0]), .A(cceip2_im_din[32]));
Q_ASSIGN U1698 ( .B(kme_cceip2_ob_out_pre[1]), .A(cceip2_im_din[33]));
Q_ASSIGN U1699 ( .B(kme_cceip2_ob_out_pre[2]), .A(cceip2_im_din[34]));
Q_ASSIGN U1700 ( .B(kme_cceip2_ob_out_pre[3]), .A(cceip2_im_din[35]));
Q_ASSIGN U1701 ( .B(kme_cceip2_ob_out_pre[4]), .A(cceip2_im_din[36]));
Q_ASSIGN U1702 ( .B(kme_cceip2_ob_out_pre[5]), .A(cceip2_im_din[37]));
Q_ASSIGN U1703 ( .B(kme_cceip2_ob_out_pre[6]), .A(cceip2_im_din[38]));
Q_ASSIGN U1704 ( .B(kme_cceip2_ob_out_pre[7]), .A(cceip2_im_din[39]));
Q_ASSIGN U1705 ( .B(kme_cceip2_ob_out_pre[8]), .A(cceip2_im_din[40]));
Q_ASSIGN U1706 ( .B(kme_cceip2_ob_out_pre[9]), .A(cceip2_im_din[41]));
Q_ASSIGN U1707 ( .B(kme_cceip2_ob_out_pre[10]), .A(cceip2_im_din[42]));
Q_ASSIGN U1708 ( .B(kme_cceip2_ob_out_pre[11]), .A(cceip2_im_din[43]));
Q_ASSIGN U1709 ( .B(kme_cceip2_ob_out_pre[12]), .A(cceip2_im_din[44]));
Q_ASSIGN U1710 ( .B(kme_cceip2_ob_out_pre[13]), .A(cceip2_im_din[45]));
Q_ASSIGN U1711 ( .B(kme_cceip2_ob_out_pre[14]), .A(cceip2_im_din[46]));
Q_ASSIGN U1712 ( .B(kme_cceip2_ob_out_pre[15]), .A(cceip2_im_din[47]));
Q_ASSIGN U1713 ( .B(kme_cceip2_ob_out_pre[16]), .A(cceip2_im_din[48]));
Q_ASSIGN U1714 ( .B(kme_cceip2_ob_out_pre[17]), .A(cceip2_im_din[49]));
Q_ASSIGN U1715 ( .B(kme_cceip2_ob_out_pre[18]), .A(cceip2_im_din[50]));
Q_ASSIGN U1716 ( .B(kme_cceip2_ob_out_pre[19]), .A(cceip2_im_din[51]));
Q_ASSIGN U1717 ( .B(kme_cceip2_ob_out_pre[20]), .A(cceip2_im_din[52]));
Q_ASSIGN U1718 ( .B(kme_cceip2_ob_out_pre[21]), .A(cceip2_im_din[53]));
Q_ASSIGN U1719 ( .B(kme_cceip2_ob_out_pre[22]), .A(cceip2_im_din[54]));
Q_ASSIGN U1720 ( .B(kme_cceip2_ob_out_pre[23]), .A(cceip2_im_din[55]));
Q_ASSIGN U1721 ( .B(kme_cceip2_ob_out_pre[24]), .A(cceip2_im_din[56]));
Q_ASSIGN U1722 ( .B(kme_cceip2_ob_out_pre[25]), .A(cceip2_im_din[57]));
Q_ASSIGN U1723 ( .B(kme_cceip2_ob_out_pre[26]), .A(cceip2_im_din[58]));
Q_ASSIGN U1724 ( .B(kme_cceip2_ob_out_pre[27]), .A(cceip2_im_din[59]));
Q_ASSIGN U1725 ( .B(kme_cceip2_ob_out_pre[28]), .A(cceip2_im_din[60]));
Q_ASSIGN U1726 ( .B(kme_cceip2_ob_out_pre[29]), .A(cceip2_im_din[61]));
Q_ASSIGN U1727 ( .B(kme_cceip2_ob_out_pre[30]), .A(cceip2_im_din[62]));
Q_ASSIGN U1728 ( .B(kme_cceip2_ob_out_pre[31]), .A(cceip2_im_din[63]));
Q_ASSIGN U1729 ( .B(kme_cceip2_ob_out_pre[32]), .A(cceip2_im_din[64]));
Q_ASSIGN U1730 ( .B(kme_cceip2_ob_out_pre[33]), .A(cceip2_im_din[65]));
Q_ASSIGN U1731 ( .B(kme_cceip2_ob_out_pre[34]), .A(cceip2_im_din[66]));
Q_ASSIGN U1732 ( .B(kme_cceip2_ob_out_pre[35]), .A(cceip2_im_din[67]));
Q_ASSIGN U1733 ( .B(kme_cceip2_ob_out_pre[36]), .A(cceip2_im_din[68]));
Q_ASSIGN U1734 ( .B(kme_cceip2_ob_out_pre[37]), .A(cceip2_im_din[69]));
Q_ASSIGN U1735 ( .B(kme_cceip2_ob_out_pre[38]), .A(cceip2_im_din[70]));
Q_ASSIGN U1736 ( .B(kme_cceip2_ob_out_pre[39]), .A(cceip2_im_din[71]));
Q_ASSIGN U1737 ( .B(kme_cceip2_ob_out_pre[40]), .A(cceip2_im_din[72]));
Q_ASSIGN U1738 ( .B(kme_cceip2_ob_out_pre[41]), .A(cceip2_im_din[73]));
Q_ASSIGN U1739 ( .B(kme_cceip2_ob_out_pre[42]), .A(cceip2_im_din[74]));
Q_ASSIGN U1740 ( .B(kme_cceip2_ob_out_pre[43]), .A(cceip2_im_din[75]));
Q_ASSIGN U1741 ( .B(kme_cceip2_ob_out_pre[44]), .A(cceip2_im_din[76]));
Q_ASSIGN U1742 ( .B(kme_cceip2_ob_out_pre[45]), .A(cceip2_im_din[77]));
Q_ASSIGN U1743 ( .B(kme_cceip2_ob_out_pre[46]), .A(cceip2_im_din[78]));
Q_ASSIGN U1744 ( .B(kme_cceip2_ob_out_pre[47]), .A(cceip2_im_din[79]));
Q_ASSIGN U1745 ( .B(kme_cceip2_ob_out_pre[48]), .A(cceip2_im_din[80]));
Q_ASSIGN U1746 ( .B(kme_cceip2_ob_out_pre[49]), .A(cceip2_im_din[81]));
Q_ASSIGN U1747 ( .B(kme_cceip2_ob_out_pre[50]), .A(cceip2_im_din[82]));
Q_ASSIGN U1748 ( .B(kme_cceip2_ob_out_pre[51]), .A(cceip2_im_din[83]));
Q_ASSIGN U1749 ( .B(kme_cceip2_ob_out_pre[52]), .A(cceip2_im_din[84]));
Q_ASSIGN U1750 ( .B(kme_cceip2_ob_out_pre[53]), .A(cceip2_im_din[85]));
Q_ASSIGN U1751 ( .B(kme_cceip2_ob_out_pre[54]), .A(cceip2_im_din[86]));
Q_ASSIGN U1752 ( .B(kme_cceip2_ob_out_pre[55]), .A(cceip2_im_din[87]));
Q_ASSIGN U1753 ( .B(kme_cceip2_ob_out_pre[56]), .A(cceip2_im_din[88]));
Q_ASSIGN U1754 ( .B(kme_cceip2_ob_out_pre[57]), .A(cceip2_im_din[89]));
Q_ASSIGN U1755 ( .B(kme_cceip2_ob_out_pre[58]), .A(cceip2_im_din[90]));
Q_ASSIGN U1756 ( .B(kme_cceip2_ob_out_pre[59]), .A(cceip2_im_din[91]));
Q_ASSIGN U1757 ( .B(kme_cceip2_ob_out_pre[60]), .A(cceip2_im_din[92]));
Q_ASSIGN U1758 ( .B(kme_cceip2_ob_out_pre[61]), .A(cceip2_im_din[93]));
Q_ASSIGN U1759 ( .B(kme_cceip2_ob_out_pre[62]), .A(cceip2_im_din[94]));
Q_ASSIGN U1760 ( .B(kme_cceip2_ob_out_pre[63]), .A(cceip2_im_din[95]));
Q_ASSIGN U1761 ( .B(kme_cddip1_ob_out_pre[64]), .A(cddip1_im_din[6]));
Q_ASSIGN U1762 ( .B(kme_cddip1_ob_out_pre[66]), .A(cddip1_im_din[8]));
Q_ASSIGN U1763 ( .B(kme_cddip1_ob_out_pre[67]), .A(cddip1_im_din[9]));
Q_ASSIGN U1764 ( .B(kme_cddip1_ob_out_pre[68]), .A(cddip1_im_din[10]));
Q_ASSIGN U1765 ( .B(kme_cddip1_ob_out_pre[69]), .A(cddip1_im_din[11]));
Q_ASSIGN U1766 ( .B(kme_cddip1_ob_out_pre[70]), .A(cddip1_im_din[12]));
Q_ASSIGN U1767 ( .B(kme_cddip1_ob_out_pre[71]), .A(cddip1_im_din[13]));
Q_ASSIGN U1768 ( .B(kme_cddip1_ob_out_pre[80]), .A(cddip1_im_din[14]));
Q_ASSIGN U1769 ( .B(kme_cddip1_ob_out_pre[72]), .A(cddip1_im_din[23]));
Q_ASSIGN U1770 ( .B(kme_cddip1_ob_out_pre[73]), .A(cddip1_im_din[24]));
Q_ASSIGN U1771 ( .B(kme_cddip1_ob_out_pre[74]), .A(cddip1_im_din[25]));
Q_ASSIGN U1772 ( .B(kme_cddip1_ob_out_pre[75]), .A(cddip1_im_din[26]));
Q_ASSIGN U1773 ( .B(kme_cddip1_ob_out_pre[76]), .A(cddip1_im_din[27]));
Q_ASSIGN U1774 ( .B(kme_cddip1_ob_out_pre[77]), .A(cddip1_im_din[28]));
Q_ASSIGN U1775 ( .B(kme_cddip1_ob_out_pre[78]), .A(cddip1_im_din[29]));
Q_ASSIGN U1776 ( .B(kme_cddip1_ob_out_pre[79]), .A(cddip1_im_din[30]));
Q_ASSIGN U1777 ( .B(kme_cddip1_ob_out_pre[65]), .A(cddip1_im_din[31]));
Q_ASSIGN U1778 ( .B(kme_cddip1_ob_out_pre[65]), .A(cddip1_im_din[7]));
Q_ASSIGN U1779 ( .B(kme_cddip1_ob_out_pre[0]), .A(cddip1_im_din[32]));
Q_ASSIGN U1780 ( .B(kme_cddip1_ob_out_pre[1]), .A(cddip1_im_din[33]));
Q_ASSIGN U1781 ( .B(kme_cddip1_ob_out_pre[2]), .A(cddip1_im_din[34]));
Q_ASSIGN U1782 ( .B(kme_cddip1_ob_out_pre[3]), .A(cddip1_im_din[35]));
Q_ASSIGN U1783 ( .B(kme_cddip1_ob_out_pre[4]), .A(cddip1_im_din[36]));
Q_ASSIGN U1784 ( .B(kme_cddip1_ob_out_pre[5]), .A(cddip1_im_din[37]));
Q_ASSIGN U1785 ( .B(kme_cddip1_ob_out_pre[6]), .A(cddip1_im_din[38]));
Q_ASSIGN U1786 ( .B(kme_cddip1_ob_out_pre[7]), .A(cddip1_im_din[39]));
Q_ASSIGN U1787 ( .B(kme_cddip1_ob_out_pre[8]), .A(cddip1_im_din[40]));
Q_ASSIGN U1788 ( .B(kme_cddip1_ob_out_pre[9]), .A(cddip1_im_din[41]));
Q_ASSIGN U1789 ( .B(kme_cddip1_ob_out_pre[10]), .A(cddip1_im_din[42]));
Q_ASSIGN U1790 ( .B(kme_cddip1_ob_out_pre[11]), .A(cddip1_im_din[43]));
Q_ASSIGN U1791 ( .B(kme_cddip1_ob_out_pre[12]), .A(cddip1_im_din[44]));
Q_ASSIGN U1792 ( .B(kme_cddip1_ob_out_pre[13]), .A(cddip1_im_din[45]));
Q_ASSIGN U1793 ( .B(kme_cddip1_ob_out_pre[14]), .A(cddip1_im_din[46]));
Q_ASSIGN U1794 ( .B(kme_cddip1_ob_out_pre[15]), .A(cddip1_im_din[47]));
Q_ASSIGN U1795 ( .B(kme_cddip1_ob_out_pre[16]), .A(cddip1_im_din[48]));
Q_ASSIGN U1796 ( .B(kme_cddip1_ob_out_pre[17]), .A(cddip1_im_din[49]));
Q_ASSIGN U1797 ( .B(kme_cddip1_ob_out_pre[18]), .A(cddip1_im_din[50]));
Q_ASSIGN U1798 ( .B(kme_cddip1_ob_out_pre[19]), .A(cddip1_im_din[51]));
Q_ASSIGN U1799 ( .B(kme_cddip1_ob_out_pre[20]), .A(cddip1_im_din[52]));
Q_ASSIGN U1800 ( .B(kme_cddip1_ob_out_pre[21]), .A(cddip1_im_din[53]));
Q_ASSIGN U1801 ( .B(kme_cddip1_ob_out_pre[22]), .A(cddip1_im_din[54]));
Q_ASSIGN U1802 ( .B(kme_cddip1_ob_out_pre[23]), .A(cddip1_im_din[55]));
Q_ASSIGN U1803 ( .B(kme_cddip1_ob_out_pre[24]), .A(cddip1_im_din[56]));
Q_ASSIGN U1804 ( .B(kme_cddip1_ob_out_pre[25]), .A(cddip1_im_din[57]));
Q_ASSIGN U1805 ( .B(kme_cddip1_ob_out_pre[26]), .A(cddip1_im_din[58]));
Q_ASSIGN U1806 ( .B(kme_cddip1_ob_out_pre[27]), .A(cddip1_im_din[59]));
Q_ASSIGN U1807 ( .B(kme_cddip1_ob_out_pre[28]), .A(cddip1_im_din[60]));
Q_ASSIGN U1808 ( .B(kme_cddip1_ob_out_pre[29]), .A(cddip1_im_din[61]));
Q_ASSIGN U1809 ( .B(kme_cddip1_ob_out_pre[30]), .A(cddip1_im_din[62]));
Q_ASSIGN U1810 ( .B(kme_cddip1_ob_out_pre[31]), .A(cddip1_im_din[63]));
Q_ASSIGN U1811 ( .B(kme_cddip1_ob_out_pre[32]), .A(cddip1_im_din[64]));
Q_ASSIGN U1812 ( .B(kme_cddip1_ob_out_pre[33]), .A(cddip1_im_din[65]));
Q_ASSIGN U1813 ( .B(kme_cddip1_ob_out_pre[34]), .A(cddip1_im_din[66]));
Q_ASSIGN U1814 ( .B(kme_cddip1_ob_out_pre[35]), .A(cddip1_im_din[67]));
Q_ASSIGN U1815 ( .B(kme_cddip1_ob_out_pre[36]), .A(cddip1_im_din[68]));
Q_ASSIGN U1816 ( .B(kme_cddip1_ob_out_pre[37]), .A(cddip1_im_din[69]));
Q_ASSIGN U1817 ( .B(kme_cddip1_ob_out_pre[38]), .A(cddip1_im_din[70]));
Q_ASSIGN U1818 ( .B(kme_cddip1_ob_out_pre[39]), .A(cddip1_im_din[71]));
Q_ASSIGN U1819 ( .B(kme_cddip1_ob_out_pre[40]), .A(cddip1_im_din[72]));
Q_ASSIGN U1820 ( .B(kme_cddip1_ob_out_pre[41]), .A(cddip1_im_din[73]));
Q_ASSIGN U1821 ( .B(kme_cddip1_ob_out_pre[42]), .A(cddip1_im_din[74]));
Q_ASSIGN U1822 ( .B(kme_cddip1_ob_out_pre[43]), .A(cddip1_im_din[75]));
Q_ASSIGN U1823 ( .B(kme_cddip1_ob_out_pre[44]), .A(cddip1_im_din[76]));
Q_ASSIGN U1824 ( .B(kme_cddip1_ob_out_pre[45]), .A(cddip1_im_din[77]));
Q_ASSIGN U1825 ( .B(kme_cddip1_ob_out_pre[46]), .A(cddip1_im_din[78]));
Q_ASSIGN U1826 ( .B(kme_cddip1_ob_out_pre[47]), .A(cddip1_im_din[79]));
Q_ASSIGN U1827 ( .B(kme_cddip1_ob_out_pre[48]), .A(cddip1_im_din[80]));
Q_ASSIGN U1828 ( .B(kme_cddip1_ob_out_pre[49]), .A(cddip1_im_din[81]));
Q_ASSIGN U1829 ( .B(kme_cddip1_ob_out_pre[50]), .A(cddip1_im_din[82]));
Q_ASSIGN U1830 ( .B(kme_cddip1_ob_out_pre[51]), .A(cddip1_im_din[83]));
Q_ASSIGN U1831 ( .B(kme_cddip1_ob_out_pre[52]), .A(cddip1_im_din[84]));
Q_ASSIGN U1832 ( .B(kme_cddip1_ob_out_pre[53]), .A(cddip1_im_din[85]));
Q_ASSIGN U1833 ( .B(kme_cddip1_ob_out_pre[54]), .A(cddip1_im_din[86]));
Q_ASSIGN U1834 ( .B(kme_cddip1_ob_out_pre[55]), .A(cddip1_im_din[87]));
Q_ASSIGN U1835 ( .B(kme_cddip1_ob_out_pre[56]), .A(cddip1_im_din[88]));
Q_ASSIGN U1836 ( .B(kme_cddip1_ob_out_pre[57]), .A(cddip1_im_din[89]));
Q_ASSIGN U1837 ( .B(kme_cddip1_ob_out_pre[58]), .A(cddip1_im_din[90]));
Q_ASSIGN U1838 ( .B(kme_cddip1_ob_out_pre[59]), .A(cddip1_im_din[91]));
Q_ASSIGN U1839 ( .B(kme_cddip1_ob_out_pre[60]), .A(cddip1_im_din[92]));
Q_ASSIGN U1840 ( .B(kme_cddip1_ob_out_pre[61]), .A(cddip1_im_din[93]));
Q_ASSIGN U1841 ( .B(kme_cddip1_ob_out_pre[62]), .A(cddip1_im_din[94]));
Q_ASSIGN U1842 ( .B(kme_cddip1_ob_out_pre[63]), .A(cddip1_im_din[95]));
Q_ASSIGN U1843 ( .B(kme_cceip1_ob_out_pre[64]), .A(cceip1_im_din[6]));
Q_ASSIGN U1844 ( .B(kme_cceip1_ob_out_pre[66]), .A(cceip1_im_din[8]));
Q_ASSIGN U1845 ( .B(kme_cceip1_ob_out_pre[67]), .A(cceip1_im_din[9]));
Q_ASSIGN U1846 ( .B(kme_cceip1_ob_out_pre[68]), .A(cceip1_im_din[10]));
Q_ASSIGN U1847 ( .B(kme_cceip1_ob_out_pre[69]), .A(cceip1_im_din[11]));
Q_ASSIGN U1848 ( .B(kme_cceip1_ob_out_pre[70]), .A(cceip1_im_din[12]));
Q_ASSIGN U1849 ( .B(kme_cceip1_ob_out_pre[71]), .A(cceip1_im_din[13]));
Q_ASSIGN U1850 ( .B(kme_cceip1_ob_out_pre[80]), .A(cceip1_im_din[14]));
Q_ASSIGN U1851 ( .B(kme_cceip1_ob_out_pre[72]), .A(cceip1_im_din[23]));
Q_ASSIGN U1852 ( .B(kme_cceip1_ob_out_pre[73]), .A(cceip1_im_din[24]));
Q_ASSIGN U1853 ( .B(kme_cceip1_ob_out_pre[74]), .A(cceip1_im_din[25]));
Q_ASSIGN U1854 ( .B(kme_cceip1_ob_out_pre[75]), .A(cceip1_im_din[26]));
Q_ASSIGN U1855 ( .B(kme_cceip1_ob_out_pre[76]), .A(cceip1_im_din[27]));
Q_ASSIGN U1856 ( .B(kme_cceip1_ob_out_pre[77]), .A(cceip1_im_din[28]));
Q_ASSIGN U1857 ( .B(kme_cceip1_ob_out_pre[78]), .A(cceip1_im_din[29]));
Q_ASSIGN U1858 ( .B(kme_cceip1_ob_out_pre[79]), .A(cceip1_im_din[30]));
Q_ASSIGN U1859 ( .B(kme_cceip1_ob_out_pre[65]), .A(cceip1_im_din[31]));
Q_ASSIGN U1860 ( .B(kme_cceip1_ob_out_pre[65]), .A(cceip1_im_din[7]));
Q_ASSIGN U1861 ( .B(kme_cceip1_ob_out_pre[0]), .A(cceip1_im_din[32]));
Q_ASSIGN U1862 ( .B(kme_cceip1_ob_out_pre[1]), .A(cceip1_im_din[33]));
Q_ASSIGN U1863 ( .B(kme_cceip1_ob_out_pre[2]), .A(cceip1_im_din[34]));
Q_ASSIGN U1864 ( .B(kme_cceip1_ob_out_pre[3]), .A(cceip1_im_din[35]));
Q_ASSIGN U1865 ( .B(kme_cceip1_ob_out_pre[4]), .A(cceip1_im_din[36]));
Q_ASSIGN U1866 ( .B(kme_cceip1_ob_out_pre[5]), .A(cceip1_im_din[37]));
Q_ASSIGN U1867 ( .B(kme_cceip1_ob_out_pre[6]), .A(cceip1_im_din[38]));
Q_ASSIGN U1868 ( .B(kme_cceip1_ob_out_pre[7]), .A(cceip1_im_din[39]));
Q_ASSIGN U1869 ( .B(kme_cceip1_ob_out_pre[8]), .A(cceip1_im_din[40]));
Q_ASSIGN U1870 ( .B(kme_cceip1_ob_out_pre[9]), .A(cceip1_im_din[41]));
Q_ASSIGN U1871 ( .B(kme_cceip1_ob_out_pre[10]), .A(cceip1_im_din[42]));
Q_ASSIGN U1872 ( .B(kme_cceip1_ob_out_pre[11]), .A(cceip1_im_din[43]));
Q_ASSIGN U1873 ( .B(kme_cceip1_ob_out_pre[12]), .A(cceip1_im_din[44]));
Q_ASSIGN U1874 ( .B(kme_cceip1_ob_out_pre[13]), .A(cceip1_im_din[45]));
Q_ASSIGN U1875 ( .B(kme_cceip1_ob_out_pre[14]), .A(cceip1_im_din[46]));
Q_ASSIGN U1876 ( .B(kme_cceip1_ob_out_pre[15]), .A(cceip1_im_din[47]));
Q_ASSIGN U1877 ( .B(kme_cceip1_ob_out_pre[16]), .A(cceip1_im_din[48]));
Q_ASSIGN U1878 ( .B(kme_cceip1_ob_out_pre[17]), .A(cceip1_im_din[49]));
Q_ASSIGN U1879 ( .B(kme_cceip1_ob_out_pre[18]), .A(cceip1_im_din[50]));
Q_ASSIGN U1880 ( .B(kme_cceip1_ob_out_pre[19]), .A(cceip1_im_din[51]));
Q_ASSIGN U1881 ( .B(kme_cceip1_ob_out_pre[20]), .A(cceip1_im_din[52]));
Q_ASSIGN U1882 ( .B(kme_cceip1_ob_out_pre[21]), .A(cceip1_im_din[53]));
Q_ASSIGN U1883 ( .B(kme_cceip1_ob_out_pre[22]), .A(cceip1_im_din[54]));
Q_ASSIGN U1884 ( .B(kme_cceip1_ob_out_pre[23]), .A(cceip1_im_din[55]));
Q_ASSIGN U1885 ( .B(kme_cceip1_ob_out_pre[24]), .A(cceip1_im_din[56]));
Q_ASSIGN U1886 ( .B(kme_cceip1_ob_out_pre[25]), .A(cceip1_im_din[57]));
Q_ASSIGN U1887 ( .B(kme_cceip1_ob_out_pre[26]), .A(cceip1_im_din[58]));
Q_ASSIGN U1888 ( .B(kme_cceip1_ob_out_pre[27]), .A(cceip1_im_din[59]));
Q_ASSIGN U1889 ( .B(kme_cceip1_ob_out_pre[28]), .A(cceip1_im_din[60]));
Q_ASSIGN U1890 ( .B(kme_cceip1_ob_out_pre[29]), .A(cceip1_im_din[61]));
Q_ASSIGN U1891 ( .B(kme_cceip1_ob_out_pre[30]), .A(cceip1_im_din[62]));
Q_ASSIGN U1892 ( .B(kme_cceip1_ob_out_pre[31]), .A(cceip1_im_din[63]));
Q_ASSIGN U1893 ( .B(kme_cceip1_ob_out_pre[32]), .A(cceip1_im_din[64]));
Q_ASSIGN U1894 ( .B(kme_cceip1_ob_out_pre[33]), .A(cceip1_im_din[65]));
Q_ASSIGN U1895 ( .B(kme_cceip1_ob_out_pre[34]), .A(cceip1_im_din[66]));
Q_ASSIGN U1896 ( .B(kme_cceip1_ob_out_pre[35]), .A(cceip1_im_din[67]));
Q_ASSIGN U1897 ( .B(kme_cceip1_ob_out_pre[36]), .A(cceip1_im_din[68]));
Q_ASSIGN U1898 ( .B(kme_cceip1_ob_out_pre[37]), .A(cceip1_im_din[69]));
Q_ASSIGN U1899 ( .B(kme_cceip1_ob_out_pre[38]), .A(cceip1_im_din[70]));
Q_ASSIGN U1900 ( .B(kme_cceip1_ob_out_pre[39]), .A(cceip1_im_din[71]));
Q_ASSIGN U1901 ( .B(kme_cceip1_ob_out_pre[40]), .A(cceip1_im_din[72]));
Q_ASSIGN U1902 ( .B(kme_cceip1_ob_out_pre[41]), .A(cceip1_im_din[73]));
Q_ASSIGN U1903 ( .B(kme_cceip1_ob_out_pre[42]), .A(cceip1_im_din[74]));
Q_ASSIGN U1904 ( .B(kme_cceip1_ob_out_pre[43]), .A(cceip1_im_din[75]));
Q_ASSIGN U1905 ( .B(kme_cceip1_ob_out_pre[44]), .A(cceip1_im_din[76]));
Q_ASSIGN U1906 ( .B(kme_cceip1_ob_out_pre[45]), .A(cceip1_im_din[77]));
Q_ASSIGN U1907 ( .B(kme_cceip1_ob_out_pre[46]), .A(cceip1_im_din[78]));
Q_ASSIGN U1908 ( .B(kme_cceip1_ob_out_pre[47]), .A(cceip1_im_din[79]));
Q_ASSIGN U1909 ( .B(kme_cceip1_ob_out_pre[48]), .A(cceip1_im_din[80]));
Q_ASSIGN U1910 ( .B(kme_cceip1_ob_out_pre[49]), .A(cceip1_im_din[81]));
Q_ASSIGN U1911 ( .B(kme_cceip1_ob_out_pre[50]), .A(cceip1_im_din[82]));
Q_ASSIGN U1912 ( .B(kme_cceip1_ob_out_pre[51]), .A(cceip1_im_din[83]));
Q_ASSIGN U1913 ( .B(kme_cceip1_ob_out_pre[52]), .A(cceip1_im_din[84]));
Q_ASSIGN U1914 ( .B(kme_cceip1_ob_out_pre[53]), .A(cceip1_im_din[85]));
Q_ASSIGN U1915 ( .B(kme_cceip1_ob_out_pre[54]), .A(cceip1_im_din[86]));
Q_ASSIGN U1916 ( .B(kme_cceip1_ob_out_pre[55]), .A(cceip1_im_din[87]));
Q_ASSIGN U1917 ( .B(kme_cceip1_ob_out_pre[56]), .A(cceip1_im_din[88]));
Q_ASSIGN U1918 ( .B(kme_cceip1_ob_out_pre[57]), .A(cceip1_im_din[89]));
Q_ASSIGN U1919 ( .B(kme_cceip1_ob_out_pre[58]), .A(cceip1_im_din[90]));
Q_ASSIGN U1920 ( .B(kme_cceip1_ob_out_pre[59]), .A(cceip1_im_din[91]));
Q_ASSIGN U1921 ( .B(kme_cceip1_ob_out_pre[60]), .A(cceip1_im_din[92]));
Q_ASSIGN U1922 ( .B(kme_cceip1_ob_out_pre[61]), .A(cceip1_im_din[93]));
Q_ASSIGN U1923 ( .B(kme_cceip1_ob_out_pre[62]), .A(cceip1_im_din[94]));
Q_ASSIGN U1924 ( .B(kme_cceip1_ob_out_pre[63]), .A(cceip1_im_din[95]));
Q_ASSIGN U1925 ( .B(kme_cddip0_ob_out_pre[64]), .A(cddip0_im_din[6]));
Q_ASSIGN U1926 ( .B(kme_cddip0_ob_out_pre[66]), .A(cddip0_im_din[8]));
Q_ASSIGN U1927 ( .B(kme_cddip0_ob_out_pre[67]), .A(cddip0_im_din[9]));
Q_ASSIGN U1928 ( .B(kme_cddip0_ob_out_pre[68]), .A(cddip0_im_din[10]));
Q_ASSIGN U1929 ( .B(kme_cddip0_ob_out_pre[69]), .A(cddip0_im_din[11]));
Q_ASSIGN U1930 ( .B(kme_cddip0_ob_out_pre[70]), .A(cddip0_im_din[12]));
Q_ASSIGN U1931 ( .B(kme_cddip0_ob_out_pre[71]), .A(cddip0_im_din[13]));
Q_ASSIGN U1932 ( .B(kme_cddip0_ob_out_pre[80]), .A(cddip0_im_din[14]));
Q_ASSIGN U1933 ( .B(kme_cddip0_ob_out_pre[72]), .A(cddip0_im_din[23]));
Q_ASSIGN U1934 ( .B(kme_cddip0_ob_out_pre[73]), .A(cddip0_im_din[24]));
Q_ASSIGN U1935 ( .B(kme_cddip0_ob_out_pre[74]), .A(cddip0_im_din[25]));
Q_ASSIGN U1936 ( .B(kme_cddip0_ob_out_pre[75]), .A(cddip0_im_din[26]));
Q_ASSIGN U1937 ( .B(kme_cddip0_ob_out_pre[76]), .A(cddip0_im_din[27]));
Q_ASSIGN U1938 ( .B(kme_cddip0_ob_out_pre[77]), .A(cddip0_im_din[28]));
Q_ASSIGN U1939 ( .B(kme_cddip0_ob_out_pre[78]), .A(cddip0_im_din[29]));
Q_ASSIGN U1940 ( .B(kme_cddip0_ob_out_pre[79]), .A(cddip0_im_din[30]));
Q_ASSIGN U1941 ( .B(kme_cddip0_ob_out_pre[65]), .A(cddip0_im_din[31]));
Q_ASSIGN U1942 ( .B(kme_cddip0_ob_out_pre[65]), .A(cddip0_im_din[7]));
Q_ASSIGN U1943 ( .B(kme_cddip0_ob_out_pre[0]), .A(cddip0_im_din[32]));
Q_ASSIGN U1944 ( .B(kme_cddip0_ob_out_pre[1]), .A(cddip0_im_din[33]));
Q_ASSIGN U1945 ( .B(kme_cddip0_ob_out_pre[2]), .A(cddip0_im_din[34]));
Q_ASSIGN U1946 ( .B(kme_cddip0_ob_out_pre[3]), .A(cddip0_im_din[35]));
Q_ASSIGN U1947 ( .B(kme_cddip0_ob_out_pre[4]), .A(cddip0_im_din[36]));
Q_ASSIGN U1948 ( .B(kme_cddip0_ob_out_pre[5]), .A(cddip0_im_din[37]));
Q_ASSIGN U1949 ( .B(kme_cddip0_ob_out_pre[6]), .A(cddip0_im_din[38]));
Q_ASSIGN U1950 ( .B(kme_cddip0_ob_out_pre[7]), .A(cddip0_im_din[39]));
Q_ASSIGN U1951 ( .B(kme_cddip0_ob_out_pre[8]), .A(cddip0_im_din[40]));
Q_ASSIGN U1952 ( .B(kme_cddip0_ob_out_pre[9]), .A(cddip0_im_din[41]));
Q_ASSIGN U1953 ( .B(kme_cddip0_ob_out_pre[10]), .A(cddip0_im_din[42]));
Q_ASSIGN U1954 ( .B(kme_cddip0_ob_out_pre[11]), .A(cddip0_im_din[43]));
Q_ASSIGN U1955 ( .B(kme_cddip0_ob_out_pre[12]), .A(cddip0_im_din[44]));
Q_ASSIGN U1956 ( .B(kme_cddip0_ob_out_pre[13]), .A(cddip0_im_din[45]));
Q_ASSIGN U1957 ( .B(kme_cddip0_ob_out_pre[14]), .A(cddip0_im_din[46]));
Q_ASSIGN U1958 ( .B(kme_cddip0_ob_out_pre[15]), .A(cddip0_im_din[47]));
Q_ASSIGN U1959 ( .B(kme_cddip0_ob_out_pre[16]), .A(cddip0_im_din[48]));
Q_ASSIGN U1960 ( .B(kme_cddip0_ob_out_pre[17]), .A(cddip0_im_din[49]));
Q_ASSIGN U1961 ( .B(kme_cddip0_ob_out_pre[18]), .A(cddip0_im_din[50]));
Q_ASSIGN U1962 ( .B(kme_cddip0_ob_out_pre[19]), .A(cddip0_im_din[51]));
Q_ASSIGN U1963 ( .B(kme_cddip0_ob_out_pre[20]), .A(cddip0_im_din[52]));
Q_ASSIGN U1964 ( .B(kme_cddip0_ob_out_pre[21]), .A(cddip0_im_din[53]));
Q_ASSIGN U1965 ( .B(kme_cddip0_ob_out_pre[22]), .A(cddip0_im_din[54]));
Q_ASSIGN U1966 ( .B(kme_cddip0_ob_out_pre[23]), .A(cddip0_im_din[55]));
Q_ASSIGN U1967 ( .B(kme_cddip0_ob_out_pre[24]), .A(cddip0_im_din[56]));
Q_ASSIGN U1968 ( .B(kme_cddip0_ob_out_pre[25]), .A(cddip0_im_din[57]));
Q_ASSIGN U1969 ( .B(kme_cddip0_ob_out_pre[26]), .A(cddip0_im_din[58]));
Q_ASSIGN U1970 ( .B(kme_cddip0_ob_out_pre[27]), .A(cddip0_im_din[59]));
Q_ASSIGN U1971 ( .B(kme_cddip0_ob_out_pre[28]), .A(cddip0_im_din[60]));
Q_ASSIGN U1972 ( .B(kme_cddip0_ob_out_pre[29]), .A(cddip0_im_din[61]));
Q_ASSIGN U1973 ( .B(kme_cddip0_ob_out_pre[30]), .A(cddip0_im_din[62]));
Q_ASSIGN U1974 ( .B(kme_cddip0_ob_out_pre[31]), .A(cddip0_im_din[63]));
Q_ASSIGN U1975 ( .B(kme_cddip0_ob_out_pre[32]), .A(cddip0_im_din[64]));
Q_ASSIGN U1976 ( .B(kme_cddip0_ob_out_pre[33]), .A(cddip0_im_din[65]));
Q_ASSIGN U1977 ( .B(kme_cddip0_ob_out_pre[34]), .A(cddip0_im_din[66]));
Q_ASSIGN U1978 ( .B(kme_cddip0_ob_out_pre[35]), .A(cddip0_im_din[67]));
Q_ASSIGN U1979 ( .B(kme_cddip0_ob_out_pre[36]), .A(cddip0_im_din[68]));
Q_ASSIGN U1980 ( .B(kme_cddip0_ob_out_pre[37]), .A(cddip0_im_din[69]));
Q_ASSIGN U1981 ( .B(kme_cddip0_ob_out_pre[38]), .A(cddip0_im_din[70]));
Q_ASSIGN U1982 ( .B(kme_cddip0_ob_out_pre[39]), .A(cddip0_im_din[71]));
Q_ASSIGN U1983 ( .B(kme_cddip0_ob_out_pre[40]), .A(cddip0_im_din[72]));
Q_ASSIGN U1984 ( .B(kme_cddip0_ob_out_pre[41]), .A(cddip0_im_din[73]));
Q_ASSIGN U1985 ( .B(kme_cddip0_ob_out_pre[42]), .A(cddip0_im_din[74]));
Q_ASSIGN U1986 ( .B(kme_cddip0_ob_out_pre[43]), .A(cddip0_im_din[75]));
Q_ASSIGN U1987 ( .B(kme_cddip0_ob_out_pre[44]), .A(cddip0_im_din[76]));
Q_ASSIGN U1988 ( .B(kme_cddip0_ob_out_pre[45]), .A(cddip0_im_din[77]));
Q_ASSIGN U1989 ( .B(kme_cddip0_ob_out_pre[46]), .A(cddip0_im_din[78]));
Q_ASSIGN U1990 ( .B(kme_cddip0_ob_out_pre[47]), .A(cddip0_im_din[79]));
Q_ASSIGN U1991 ( .B(kme_cddip0_ob_out_pre[48]), .A(cddip0_im_din[80]));
Q_ASSIGN U1992 ( .B(kme_cddip0_ob_out_pre[49]), .A(cddip0_im_din[81]));
Q_ASSIGN U1993 ( .B(kme_cddip0_ob_out_pre[50]), .A(cddip0_im_din[82]));
Q_ASSIGN U1994 ( .B(kme_cddip0_ob_out_pre[51]), .A(cddip0_im_din[83]));
Q_ASSIGN U1995 ( .B(kme_cddip0_ob_out_pre[52]), .A(cddip0_im_din[84]));
Q_ASSIGN U1996 ( .B(kme_cddip0_ob_out_pre[53]), .A(cddip0_im_din[85]));
Q_ASSIGN U1997 ( .B(kme_cddip0_ob_out_pre[54]), .A(cddip0_im_din[86]));
Q_ASSIGN U1998 ( .B(kme_cddip0_ob_out_pre[55]), .A(cddip0_im_din[87]));
Q_ASSIGN U1999 ( .B(kme_cddip0_ob_out_pre[56]), .A(cddip0_im_din[88]));
Q_ASSIGN U2000 ( .B(kme_cddip0_ob_out_pre[57]), .A(cddip0_im_din[89]));
Q_ASSIGN U2001 ( .B(kme_cddip0_ob_out_pre[58]), .A(cddip0_im_din[90]));
Q_ASSIGN U2002 ( .B(kme_cddip0_ob_out_pre[59]), .A(cddip0_im_din[91]));
Q_ASSIGN U2003 ( .B(kme_cddip0_ob_out_pre[60]), .A(cddip0_im_din[92]));
Q_ASSIGN U2004 ( .B(kme_cddip0_ob_out_pre[61]), .A(cddip0_im_din[93]));
Q_ASSIGN U2005 ( .B(kme_cddip0_ob_out_pre[62]), .A(cddip0_im_din[94]));
Q_ASSIGN U2006 ( .B(kme_cddip0_ob_out_pre[63]), .A(cddip0_im_din[95]));
Q_ASSIGN U2007 ( .B(kme_cceip0_ob_out_pre[64]), .A(cceip0_im_din[6]));
Q_ASSIGN U2008 ( .B(kme_cceip0_ob_out_pre[66]), .A(cceip0_im_din[8]));
Q_ASSIGN U2009 ( .B(kme_cceip0_ob_out_pre[67]), .A(cceip0_im_din[9]));
Q_ASSIGN U2010 ( .B(kme_cceip0_ob_out_pre[68]), .A(cceip0_im_din[10]));
Q_ASSIGN U2011 ( .B(kme_cceip0_ob_out_pre[69]), .A(cceip0_im_din[11]));
Q_ASSIGN U2012 ( .B(kme_cceip0_ob_out_pre[70]), .A(cceip0_im_din[12]));
Q_ASSIGN U2013 ( .B(kme_cceip0_ob_out_pre[71]), .A(cceip0_im_din[13]));
Q_ASSIGN U2014 ( .B(kme_cceip0_ob_out_pre[80]), .A(cceip0_im_din[14]));
Q_ASSIGN U2015 ( .B(kme_cceip0_ob_out_pre[72]), .A(cceip0_im_din[23]));
Q_ASSIGN U2016 ( .B(kme_cceip0_ob_out_pre[73]), .A(cceip0_im_din[24]));
Q_ASSIGN U2017 ( .B(kme_cceip0_ob_out_pre[74]), .A(cceip0_im_din[25]));
Q_ASSIGN U2018 ( .B(kme_cceip0_ob_out_pre[75]), .A(cceip0_im_din[26]));
Q_ASSIGN U2019 ( .B(kme_cceip0_ob_out_pre[76]), .A(cceip0_im_din[27]));
Q_ASSIGN U2020 ( .B(kme_cceip0_ob_out_pre[77]), .A(cceip0_im_din[28]));
Q_ASSIGN U2021 ( .B(kme_cceip0_ob_out_pre[78]), .A(cceip0_im_din[29]));
Q_ASSIGN U2022 ( .B(kme_cceip0_ob_out_pre[79]), .A(cceip0_im_din[30]));
Q_ASSIGN U2023 ( .B(kme_cceip0_ob_out_pre[65]), .A(cceip0_im_din[31]));
Q_ASSIGN U2024 ( .B(kme_cceip0_ob_out_pre[65]), .A(cceip0_im_din[7]));
Q_ASSIGN U2025 ( .B(kme_cceip0_ob_out_pre[0]), .A(cceip0_im_din[32]));
Q_ASSIGN U2026 ( .B(kme_cceip0_ob_out_pre[1]), .A(cceip0_im_din[33]));
Q_ASSIGN U2027 ( .B(kme_cceip0_ob_out_pre[2]), .A(cceip0_im_din[34]));
Q_ASSIGN U2028 ( .B(kme_cceip0_ob_out_pre[3]), .A(cceip0_im_din[35]));
Q_ASSIGN U2029 ( .B(kme_cceip0_ob_out_pre[4]), .A(cceip0_im_din[36]));
Q_ASSIGN U2030 ( .B(kme_cceip0_ob_out_pre[5]), .A(cceip0_im_din[37]));
Q_ASSIGN U2031 ( .B(kme_cceip0_ob_out_pre[6]), .A(cceip0_im_din[38]));
Q_ASSIGN U2032 ( .B(kme_cceip0_ob_out_pre[7]), .A(cceip0_im_din[39]));
Q_ASSIGN U2033 ( .B(kme_cceip0_ob_out_pre[8]), .A(cceip0_im_din[40]));
Q_ASSIGN U2034 ( .B(kme_cceip0_ob_out_pre[9]), .A(cceip0_im_din[41]));
Q_ASSIGN U2035 ( .B(kme_cceip0_ob_out_pre[10]), .A(cceip0_im_din[42]));
Q_ASSIGN U2036 ( .B(kme_cceip0_ob_out_pre[11]), .A(cceip0_im_din[43]));
Q_ASSIGN U2037 ( .B(kme_cceip0_ob_out_pre[12]), .A(cceip0_im_din[44]));
Q_ASSIGN U2038 ( .B(kme_cceip0_ob_out_pre[13]), .A(cceip0_im_din[45]));
Q_ASSIGN U2039 ( .B(kme_cceip0_ob_out_pre[14]), .A(cceip0_im_din[46]));
Q_ASSIGN U2040 ( .B(kme_cceip0_ob_out_pre[15]), .A(cceip0_im_din[47]));
Q_ASSIGN U2041 ( .B(kme_cceip0_ob_out_pre[16]), .A(cceip0_im_din[48]));
Q_ASSIGN U2042 ( .B(kme_cceip0_ob_out_pre[17]), .A(cceip0_im_din[49]));
Q_ASSIGN U2043 ( .B(kme_cceip0_ob_out_pre[18]), .A(cceip0_im_din[50]));
Q_ASSIGN U2044 ( .B(kme_cceip0_ob_out_pre[19]), .A(cceip0_im_din[51]));
Q_ASSIGN U2045 ( .B(kme_cceip0_ob_out_pre[20]), .A(cceip0_im_din[52]));
Q_ASSIGN U2046 ( .B(kme_cceip0_ob_out_pre[21]), .A(cceip0_im_din[53]));
Q_ASSIGN U2047 ( .B(kme_cceip0_ob_out_pre[22]), .A(cceip0_im_din[54]));
Q_ASSIGN U2048 ( .B(kme_cceip0_ob_out_pre[23]), .A(cceip0_im_din[55]));
Q_ASSIGN U2049 ( .B(kme_cceip0_ob_out_pre[24]), .A(cceip0_im_din[56]));
Q_ASSIGN U2050 ( .B(kme_cceip0_ob_out_pre[25]), .A(cceip0_im_din[57]));
Q_ASSIGN U2051 ( .B(kme_cceip0_ob_out_pre[26]), .A(cceip0_im_din[58]));
Q_ASSIGN U2052 ( .B(kme_cceip0_ob_out_pre[27]), .A(cceip0_im_din[59]));
Q_ASSIGN U2053 ( .B(kme_cceip0_ob_out_pre[28]), .A(cceip0_im_din[60]));
Q_ASSIGN U2054 ( .B(kme_cceip0_ob_out_pre[29]), .A(cceip0_im_din[61]));
Q_ASSIGN U2055 ( .B(kme_cceip0_ob_out_pre[30]), .A(cceip0_im_din[62]));
Q_ASSIGN U2056 ( .B(kme_cceip0_ob_out_pre[31]), .A(cceip0_im_din[63]));
Q_ASSIGN U2057 ( .B(kme_cceip0_ob_out_pre[32]), .A(cceip0_im_din[64]));
Q_ASSIGN U2058 ( .B(kme_cceip0_ob_out_pre[33]), .A(cceip0_im_din[65]));
Q_ASSIGN U2059 ( .B(kme_cceip0_ob_out_pre[34]), .A(cceip0_im_din[66]));
Q_ASSIGN U2060 ( .B(kme_cceip0_ob_out_pre[35]), .A(cceip0_im_din[67]));
Q_ASSIGN U2061 ( .B(kme_cceip0_ob_out_pre[36]), .A(cceip0_im_din[68]));
Q_ASSIGN U2062 ( .B(kme_cceip0_ob_out_pre[37]), .A(cceip0_im_din[69]));
Q_ASSIGN U2063 ( .B(kme_cceip0_ob_out_pre[38]), .A(cceip0_im_din[70]));
Q_ASSIGN U2064 ( .B(kme_cceip0_ob_out_pre[39]), .A(cceip0_im_din[71]));
Q_ASSIGN U2065 ( .B(kme_cceip0_ob_out_pre[40]), .A(cceip0_im_din[72]));
Q_ASSIGN U2066 ( .B(kme_cceip0_ob_out_pre[41]), .A(cceip0_im_din[73]));
Q_ASSIGN U2067 ( .B(kme_cceip0_ob_out_pre[42]), .A(cceip0_im_din[74]));
Q_ASSIGN U2068 ( .B(kme_cceip0_ob_out_pre[43]), .A(cceip0_im_din[75]));
Q_ASSIGN U2069 ( .B(kme_cceip0_ob_out_pre[44]), .A(cceip0_im_din[76]));
Q_ASSIGN U2070 ( .B(kme_cceip0_ob_out_pre[45]), .A(cceip0_im_din[77]));
Q_ASSIGN U2071 ( .B(kme_cceip0_ob_out_pre[46]), .A(cceip0_im_din[78]));
Q_ASSIGN U2072 ( .B(kme_cceip0_ob_out_pre[47]), .A(cceip0_im_din[79]));
Q_ASSIGN U2073 ( .B(kme_cceip0_ob_out_pre[48]), .A(cceip0_im_din[80]));
Q_ASSIGN U2074 ( .B(kme_cceip0_ob_out_pre[49]), .A(cceip0_im_din[81]));
Q_ASSIGN U2075 ( .B(kme_cceip0_ob_out_pre[50]), .A(cceip0_im_din[82]));
Q_ASSIGN U2076 ( .B(kme_cceip0_ob_out_pre[51]), .A(cceip0_im_din[83]));
Q_ASSIGN U2077 ( .B(kme_cceip0_ob_out_pre[52]), .A(cceip0_im_din[84]));
Q_ASSIGN U2078 ( .B(kme_cceip0_ob_out_pre[53]), .A(cceip0_im_din[85]));
Q_ASSIGN U2079 ( .B(kme_cceip0_ob_out_pre[54]), .A(cceip0_im_din[86]));
Q_ASSIGN U2080 ( .B(kme_cceip0_ob_out_pre[55]), .A(cceip0_im_din[87]));
Q_ASSIGN U2081 ( .B(kme_cceip0_ob_out_pre[56]), .A(cceip0_im_din[88]));
Q_ASSIGN U2082 ( .B(kme_cceip0_ob_out_pre[57]), .A(cceip0_im_din[89]));
Q_ASSIGN U2083 ( .B(kme_cceip0_ob_out_pre[58]), .A(cceip0_im_din[90]));
Q_ASSIGN U2084 ( .B(kme_cceip0_ob_out_pre[59]), .A(cceip0_im_din[91]));
Q_ASSIGN U2085 ( .B(kme_cceip0_ob_out_pre[60]), .A(cceip0_im_din[92]));
Q_ASSIGN U2086 ( .B(kme_cceip0_ob_out_pre[61]), .A(cceip0_im_din[93]));
Q_ASSIGN U2087 ( .B(kme_cceip0_ob_out_pre[62]), .A(cceip0_im_din[94]));
Q_ASSIGN U2088 ( .B(kme_cceip0_ob_out_pre[63]), .A(cceip0_im_din[95]));
ixc_assign _zz_strnp_35 ( o_send_kme_ib_beat, _zy_simnet_tvar_37);
ixc_assign _zz_strnp_34 ( o_disable_ckv_kim_ism_reads, _zy_simnet_tvar_36);
ixc_assign _zz_strnp_33 ( o_tready_override_val, _zy_simnet_tvar_35);
ixc_assign _zz_strnp_32 ( spare[3], _zy_simnet_tvar_34);
ixc_assign_25 _zz_strnp_31 ( spare[31:7], _zy_simnet_tvar_33[0:24]);
ixc_assign_84 _zz_strnp_0 ( _zy_simnet_rbus_ring_o_0_w$[0:83], 
	rbus_ring_o[83:0]);
nx_reg_indirect_access u_SA_CTRL ( .stat_code( 
	_zy_simnet_sa_ctrl_ia_status_794_w$[0:2]), .stat_datawords( 
	_zy_simnet_sa_ctrl_ia_status_795_w$[0:4]), .stat_addr( 
	_zy_simnet_sa_ctrl_ia_status_796_w$[0:4]), .capability_lst( 
	_zy_simnet_sa_ctrl_ia_capability_797_w$[0:15]), .capability_type( 
	_zy_simnet_sa_ctrl_ia_capability_798_w$[0:3]), .rd_dat( 
	_zy_simnet_sa_ctrl_ia_rdata_799_w$[0:31]), .mem_a( { \sa_ctrl[31][31] , 
	\sa_ctrl[31][30] , \sa_ctrl[31][29] , \sa_ctrl[31][28] , 
	\sa_ctrl[31][27] , \sa_ctrl[31][26] , \sa_ctrl[31][25] , 
	\sa_ctrl[31][24] , \sa_ctrl[31][23] , \sa_ctrl[31][22] , 
	\sa_ctrl[31][21] , \sa_ctrl[31][20] , \sa_ctrl[31][19] , 
	\sa_ctrl[31][18] , \sa_ctrl[31][17] , \sa_ctrl[31][16] , 
	\sa_ctrl[31][15] , \sa_ctrl[31][14] , \sa_ctrl[31][13] , 
	\sa_ctrl[31][12] , \sa_ctrl[31][11] , \sa_ctrl[31][10] , 
	\sa_ctrl[31][9] , \sa_ctrl[31][8] , \sa_ctrl[31][7] , 
	\sa_ctrl[31][6] , \sa_ctrl[31][5] , \sa_ctrl[31][4] , 
	\sa_ctrl[31][3] , \sa_ctrl[31][2] , \sa_ctrl[31][1] , 
	\sa_ctrl[31][0] , \sa_ctrl[30][31] , \sa_ctrl[30][30] , 
	\sa_ctrl[30][29] , \sa_ctrl[30][28] , \sa_ctrl[30][27] , 
	\sa_ctrl[30][26] , \sa_ctrl[30][25] , \sa_ctrl[30][24] , 
	\sa_ctrl[30][23] , \sa_ctrl[30][22] , \sa_ctrl[30][21] , 
	\sa_ctrl[30][20] , \sa_ctrl[30][19] , \sa_ctrl[30][18] , 
	\sa_ctrl[30][17] , \sa_ctrl[30][16] , \sa_ctrl[30][15] , 
	\sa_ctrl[30][14] , \sa_ctrl[30][13] , \sa_ctrl[30][12] , 
	\sa_ctrl[30][11] , \sa_ctrl[30][10] , \sa_ctrl[30][9] , 
	\sa_ctrl[30][8] , \sa_ctrl[30][7] , \sa_ctrl[30][6] , 
	\sa_ctrl[30][5] , \sa_ctrl[30][4] , \sa_ctrl[30][3] , 
	\sa_ctrl[30][2] , \sa_ctrl[30][1] , \sa_ctrl[30][0] , 
	\sa_ctrl[29][31] , \sa_ctrl[29][30] , \sa_ctrl[29][29] , 
	\sa_ctrl[29][28] , \sa_ctrl[29][27] , \sa_ctrl[29][26] , 
	\sa_ctrl[29][25] , \sa_ctrl[29][24] , \sa_ctrl[29][23] , 
	\sa_ctrl[29][22] , \sa_ctrl[29][21] , \sa_ctrl[29][20] , 
	\sa_ctrl[29][19] , \sa_ctrl[29][18] , \sa_ctrl[29][17] , 
	\sa_ctrl[29][16] , \sa_ctrl[29][15] , \sa_ctrl[29][14] , 
	\sa_ctrl[29][13] , \sa_ctrl[29][12] , \sa_ctrl[29][11] , 
	\sa_ctrl[29][10] , \sa_ctrl[29][9] , \sa_ctrl[29][8] , 
	\sa_ctrl[29][7] , \sa_ctrl[29][6] , \sa_ctrl[29][5] , 
	\sa_ctrl[29][4] , \sa_ctrl[29][3] , \sa_ctrl[29][2] , 
	\sa_ctrl[29][1] , \sa_ctrl[29][0] , \sa_ctrl[28][31] , 
	\sa_ctrl[28][30] , \sa_ctrl[28][29] , \sa_ctrl[28][28] , 
	\sa_ctrl[28][27] , \sa_ctrl[28][26] , \sa_ctrl[28][25] , 
	\sa_ctrl[28][24] , \sa_ctrl[28][23] , \sa_ctrl[28][22] , 
	\sa_ctrl[28][21] , \sa_ctrl[28][20] , \sa_ctrl[28][19] , 
	\sa_ctrl[28][18] , \sa_ctrl[28][17] , \sa_ctrl[28][16] , 
	\sa_ctrl[28][15] , \sa_ctrl[28][14] , \sa_ctrl[28][13] , 
	\sa_ctrl[28][12] , \sa_ctrl[28][11] , \sa_ctrl[28][10] , 
	\sa_ctrl[28][9] , \sa_ctrl[28][8] , \sa_ctrl[28][7] , 
	\sa_ctrl[28][6] , \sa_ctrl[28][5] , \sa_ctrl[28][4] , 
	\sa_ctrl[28][3] , \sa_ctrl[28][2] , \sa_ctrl[28][1] , 
	\sa_ctrl[28][0] , \sa_ctrl[27][31] , \sa_ctrl[27][30] , 
	\sa_ctrl[27][29] , \sa_ctrl[27][28] , \sa_ctrl[27][27] , 
	\sa_ctrl[27][26] , \sa_ctrl[27][25] , \sa_ctrl[27][24] , 
	\sa_ctrl[27][23] , \sa_ctrl[27][22] , \sa_ctrl[27][21] , 
	\sa_ctrl[27][20] , \sa_ctrl[27][19] , \sa_ctrl[27][18] , 
	\sa_ctrl[27][17] , \sa_ctrl[27][16] , \sa_ctrl[27][15] , 
	\sa_ctrl[27][14] , \sa_ctrl[27][13] , \sa_ctrl[27][12] , 
	\sa_ctrl[27][11] , \sa_ctrl[27][10] , \sa_ctrl[27][9] , 
	\sa_ctrl[27][8] , \sa_ctrl[27][7] , \sa_ctrl[27][6] , 
	\sa_ctrl[27][5] , \sa_ctrl[27][4] , \sa_ctrl[27][3] , 
	\sa_ctrl[27][2] , \sa_ctrl[27][1] , \sa_ctrl[27][0] , 
	\sa_ctrl[26][31] , \sa_ctrl[26][30] , \sa_ctrl[26][29] , 
	\sa_ctrl[26][28] , \sa_ctrl[26][27] , \sa_ctrl[26][26] , 
	\sa_ctrl[26][25] , \sa_ctrl[26][24] , \sa_ctrl[26][23] , 
	\sa_ctrl[26][22] , \sa_ctrl[26][21] , \sa_ctrl[26][20] , 
	\sa_ctrl[26][19] , \sa_ctrl[26][18] , \sa_ctrl[26][17] , 
	\sa_ctrl[26][16] , \sa_ctrl[26][15] , \sa_ctrl[26][14] , 
	\sa_ctrl[26][13] , \sa_ctrl[26][12] , \sa_ctrl[26][11] , 
	\sa_ctrl[26][10] , \sa_ctrl[26][9] , \sa_ctrl[26][8] , 
	\sa_ctrl[26][7] , \sa_ctrl[26][6] , \sa_ctrl[26][5] , 
	\sa_ctrl[26][4] , \sa_ctrl[26][3] , \sa_ctrl[26][2] , 
	\sa_ctrl[26][1] , \sa_ctrl[26][0] , \sa_ctrl[25][31] , 
	\sa_ctrl[25][30] , \sa_ctrl[25][29] , \sa_ctrl[25][28] , 
	\sa_ctrl[25][27] , \sa_ctrl[25][26] , \sa_ctrl[25][25] , 
	\sa_ctrl[25][24] , \sa_ctrl[25][23] , \sa_ctrl[25][22] , 
	\sa_ctrl[25][21] , \sa_ctrl[25][20] , \sa_ctrl[25][19] , 
	\sa_ctrl[25][18] , \sa_ctrl[25][17] , \sa_ctrl[25][16] , 
	\sa_ctrl[25][15] , \sa_ctrl[25][14] , \sa_ctrl[25][13] , 
	\sa_ctrl[25][12] , \sa_ctrl[25][11] , \sa_ctrl[25][10] , 
	\sa_ctrl[25][9] , \sa_ctrl[25][8] , \sa_ctrl[25][7] , 
	\sa_ctrl[25][6] , \sa_ctrl[25][5] , \sa_ctrl[25][4] , 
	\sa_ctrl[25][3] , \sa_ctrl[25][2] , \sa_ctrl[25][1] , 
	\sa_ctrl[25][0] , \sa_ctrl[24][31] , \sa_ctrl[24][30] , 
	\sa_ctrl[24][29] , \sa_ctrl[24][28] , \sa_ctrl[24][27] , 
	\sa_ctrl[24][26] , \sa_ctrl[24][25] , \sa_ctrl[24][24] , 
	\sa_ctrl[24][23] , \sa_ctrl[24][22] , \sa_ctrl[24][21] , 
	\sa_ctrl[24][20] , \sa_ctrl[24][19] , \sa_ctrl[24][18] , 
	\sa_ctrl[24][17] , \sa_ctrl[24][16] , \sa_ctrl[24][15] , 
	\sa_ctrl[24][14] , \sa_ctrl[24][13] , \sa_ctrl[24][12] , 
	\sa_ctrl[24][11] , \sa_ctrl[24][10] , \sa_ctrl[24][9] , 
	\sa_ctrl[24][8] , \sa_ctrl[24][7] , \sa_ctrl[24][6] , 
	\sa_ctrl[24][5] , \sa_ctrl[24][4] , \sa_ctrl[24][3] , 
	\sa_ctrl[24][2] , \sa_ctrl[24][1] , \sa_ctrl[24][0] , 
	\sa_ctrl[23][31] , \sa_ctrl[23][30] , \sa_ctrl[23][29] , 
	\sa_ctrl[23][28] , \sa_ctrl[23][27] , \sa_ctrl[23][26] , 
	\sa_ctrl[23][25] , \sa_ctrl[23][24] , \sa_ctrl[23][23] , 
	\sa_ctrl[23][22] , \sa_ctrl[23][21] , \sa_ctrl[23][20] , 
	\sa_ctrl[23][19] , \sa_ctrl[23][18] , \sa_ctrl[23][17] , 
	\sa_ctrl[23][16] , \sa_ctrl[23][15] , \sa_ctrl[23][14] , 
	\sa_ctrl[23][13] , \sa_ctrl[23][12] , \sa_ctrl[23][11] , 
	\sa_ctrl[23][10] , \sa_ctrl[23][9] , \sa_ctrl[23][8] , 
	\sa_ctrl[23][7] , \sa_ctrl[23][6] , \sa_ctrl[23][5] , 
	\sa_ctrl[23][4] , \sa_ctrl[23][3] , \sa_ctrl[23][2] , 
	\sa_ctrl[23][1] , \sa_ctrl[23][0] , \sa_ctrl[22][31] , 
	\sa_ctrl[22][30] , \sa_ctrl[22][29] , \sa_ctrl[22][28] , 
	\sa_ctrl[22][27] , \sa_ctrl[22][26] , \sa_ctrl[22][25] , 
	\sa_ctrl[22][24] , \sa_ctrl[22][23] , \sa_ctrl[22][22] , 
	\sa_ctrl[22][21] , \sa_ctrl[22][20] , \sa_ctrl[22][19] , 
	\sa_ctrl[22][18] , \sa_ctrl[22][17] , \sa_ctrl[22][16] , 
	\sa_ctrl[22][15] , \sa_ctrl[22][14] , \sa_ctrl[22][13] , 
	\sa_ctrl[22][12] , \sa_ctrl[22][11] , \sa_ctrl[22][10] , 
	\sa_ctrl[22][9] , \sa_ctrl[22][8] , \sa_ctrl[22][7] , 
	\sa_ctrl[22][6] , \sa_ctrl[22][5] , \sa_ctrl[22][4] , 
	\sa_ctrl[22][3] , \sa_ctrl[22][2] , \sa_ctrl[22][1] , 
	\sa_ctrl[22][0] , \sa_ctrl[21][31] , \sa_ctrl[21][30] , 
	\sa_ctrl[21][29] , \sa_ctrl[21][28] , \sa_ctrl[21][27] , 
	\sa_ctrl[21][26] , \sa_ctrl[21][25] , \sa_ctrl[21][24] , 
	\sa_ctrl[21][23] , \sa_ctrl[21][22] , \sa_ctrl[21][21] , 
	\sa_ctrl[21][20] , \sa_ctrl[21][19] , \sa_ctrl[21][18] , 
	\sa_ctrl[21][17] , \sa_ctrl[21][16] , \sa_ctrl[21][15] , 
	\sa_ctrl[21][14] , \sa_ctrl[21][13] , \sa_ctrl[21][12] , 
	\sa_ctrl[21][11] , \sa_ctrl[21][10] , \sa_ctrl[21][9] , 
	\sa_ctrl[21][8] , \sa_ctrl[21][7] , \sa_ctrl[21][6] , 
	\sa_ctrl[21][5] , \sa_ctrl[21][4] , \sa_ctrl[21][3] , 
	\sa_ctrl[21][2] , \sa_ctrl[21][1] , \sa_ctrl[21][0] , 
	\sa_ctrl[20][31] , \sa_ctrl[20][30] , \sa_ctrl[20][29] , 
	\sa_ctrl[20][28] , \sa_ctrl[20][27] , \sa_ctrl[20][26] , 
	\sa_ctrl[20][25] , \sa_ctrl[20][24] , \sa_ctrl[20][23] , 
	\sa_ctrl[20][22] , \sa_ctrl[20][21] , \sa_ctrl[20][20] , 
	\sa_ctrl[20][19] , \sa_ctrl[20][18] , \sa_ctrl[20][17] , 
	\sa_ctrl[20][16] , \sa_ctrl[20][15] , \sa_ctrl[20][14] , 
	\sa_ctrl[20][13] , \sa_ctrl[20][12] , \sa_ctrl[20][11] , 
	\sa_ctrl[20][10] , \sa_ctrl[20][9] , \sa_ctrl[20][8] , 
	\sa_ctrl[20][7] , \sa_ctrl[20][6] , \sa_ctrl[20][5] , 
	\sa_ctrl[20][4] , \sa_ctrl[20][3] , \sa_ctrl[20][2] , 
	\sa_ctrl[20][1] , \sa_ctrl[20][0] , \sa_ctrl[19][31] , 
	\sa_ctrl[19][30] , \sa_ctrl[19][29] , \sa_ctrl[19][28] , 
	\sa_ctrl[19][27] , \sa_ctrl[19][26] , \sa_ctrl[19][25] , 
	\sa_ctrl[19][24] , \sa_ctrl[19][23] , \sa_ctrl[19][22] , 
	\sa_ctrl[19][21] , \sa_ctrl[19][20] , \sa_ctrl[19][19] , 
	\sa_ctrl[19][18] , \sa_ctrl[19][17] , \sa_ctrl[19][16] , 
	\sa_ctrl[19][15] , \sa_ctrl[19][14] , \sa_ctrl[19][13] , 
	\sa_ctrl[19][12] , \sa_ctrl[19][11] , \sa_ctrl[19][10] , 
	\sa_ctrl[19][9] , \sa_ctrl[19][8] , \sa_ctrl[19][7] , 
	\sa_ctrl[19][6] , \sa_ctrl[19][5] , \sa_ctrl[19][4] , 
	\sa_ctrl[19][3] , \sa_ctrl[19][2] , \sa_ctrl[19][1] , 
	\sa_ctrl[19][0] , \sa_ctrl[18][31] , \sa_ctrl[18][30] , 
	\sa_ctrl[18][29] , \sa_ctrl[18][28] , \sa_ctrl[18][27] , 
	\sa_ctrl[18][26] , \sa_ctrl[18][25] , \sa_ctrl[18][24] , 
	\sa_ctrl[18][23] , \sa_ctrl[18][22] , \sa_ctrl[18][21] , 
	\sa_ctrl[18][20] , \sa_ctrl[18][19] , \sa_ctrl[18][18] , 
	\sa_ctrl[18][17] , \sa_ctrl[18][16] , \sa_ctrl[18][15] , 
	\sa_ctrl[18][14] , \sa_ctrl[18][13] , \sa_ctrl[18][12] , 
	\sa_ctrl[18][11] , \sa_ctrl[18][10] , \sa_ctrl[18][9] , 
	\sa_ctrl[18][8] , \sa_ctrl[18][7] , \sa_ctrl[18][6] , 
	\sa_ctrl[18][5] , \sa_ctrl[18][4] , \sa_ctrl[18][3] , 
	\sa_ctrl[18][2] , \sa_ctrl[18][1] , \sa_ctrl[18][0] , 
	\sa_ctrl[17][31] , \sa_ctrl[17][30] , \sa_ctrl[17][29] , 
	\sa_ctrl[17][28] , \sa_ctrl[17][27] , \sa_ctrl[17][26] , 
	\sa_ctrl[17][25] , \sa_ctrl[17][24] , \sa_ctrl[17][23] , 
	\sa_ctrl[17][22] , \sa_ctrl[17][21] , \sa_ctrl[17][20] , 
	\sa_ctrl[17][19] , \sa_ctrl[17][18] , \sa_ctrl[17][17] , 
	\sa_ctrl[17][16] , \sa_ctrl[17][15] , \sa_ctrl[17][14] , 
	\sa_ctrl[17][13] , \sa_ctrl[17][12] , \sa_ctrl[17][11] , 
	\sa_ctrl[17][10] , \sa_ctrl[17][9] , \sa_ctrl[17][8] , 
	\sa_ctrl[17][7] , \sa_ctrl[17][6] , \sa_ctrl[17][5] , 
	\sa_ctrl[17][4] , \sa_ctrl[17][3] , \sa_ctrl[17][2] , 
	\sa_ctrl[17][1] , \sa_ctrl[17][0] , \sa_ctrl[16][31] , 
	\sa_ctrl[16][30] , \sa_ctrl[16][29] , \sa_ctrl[16][28] , 
	\sa_ctrl[16][27] , \sa_ctrl[16][26] , \sa_ctrl[16][25] , 
	\sa_ctrl[16][24] , \sa_ctrl[16][23] , \sa_ctrl[16][22] , 
	\sa_ctrl[16][21] , \sa_ctrl[16][20] , \sa_ctrl[16][19] , 
	\sa_ctrl[16][18] , \sa_ctrl[16][17] , \sa_ctrl[16][16] , 
	\sa_ctrl[16][15] , \sa_ctrl[16][14] , \sa_ctrl[16][13] , 
	\sa_ctrl[16][12] , \sa_ctrl[16][11] , \sa_ctrl[16][10] , 
	\sa_ctrl[16][9] , \sa_ctrl[16][8] , \sa_ctrl[16][7] , 
	\sa_ctrl[16][6] , \sa_ctrl[16][5] , \sa_ctrl[16][4] , 
	\sa_ctrl[16][3] , \sa_ctrl[16][2] , \sa_ctrl[16][1] , 
	\sa_ctrl[16][0] , \sa_ctrl[15][31] , \sa_ctrl[15][30] , 
	\sa_ctrl[15][29] , \sa_ctrl[15][28] , \sa_ctrl[15][27] , 
	\sa_ctrl[15][26] , \sa_ctrl[15][25] , \sa_ctrl[15][24] , 
	\sa_ctrl[15][23] , \sa_ctrl[15][22] , \sa_ctrl[15][21] , 
	\sa_ctrl[15][20] , \sa_ctrl[15][19] , \sa_ctrl[15][18] , 
	\sa_ctrl[15][17] , \sa_ctrl[15][16] , \sa_ctrl[15][15] , 
	\sa_ctrl[15][14] , \sa_ctrl[15][13] , \sa_ctrl[15][12] , 
	\sa_ctrl[15][11] , \sa_ctrl[15][10] , \sa_ctrl[15][9] , 
	\sa_ctrl[15][8] , \sa_ctrl[15][7] , \sa_ctrl[15][6] , 
	\sa_ctrl[15][5] , \sa_ctrl[15][4] , \sa_ctrl[15][3] , 
	\sa_ctrl[15][2] , \sa_ctrl[15][1] , \sa_ctrl[15][0] , 
	\sa_ctrl[14][31] , \sa_ctrl[14][30] , \sa_ctrl[14][29] , 
	\sa_ctrl[14][28] , \sa_ctrl[14][27] , \sa_ctrl[14][26] , 
	\sa_ctrl[14][25] , \sa_ctrl[14][24] , \sa_ctrl[14][23] , 
	\sa_ctrl[14][22] , \sa_ctrl[14][21] , \sa_ctrl[14][20] , 
	\sa_ctrl[14][19] , \sa_ctrl[14][18] , \sa_ctrl[14][17] , 
	\sa_ctrl[14][16] , \sa_ctrl[14][15] , \sa_ctrl[14][14] , 
	\sa_ctrl[14][13] , \sa_ctrl[14][12] , \sa_ctrl[14][11] , 
	\sa_ctrl[14][10] , \sa_ctrl[14][9] , \sa_ctrl[14][8] , 
	\sa_ctrl[14][7] , \sa_ctrl[14][6] , \sa_ctrl[14][5] , 
	\sa_ctrl[14][4] , \sa_ctrl[14][3] , \sa_ctrl[14][2] , 
	\sa_ctrl[14][1] , \sa_ctrl[14][0] , \sa_ctrl[13][31] , 
	\sa_ctrl[13][30] , \sa_ctrl[13][29] , \sa_ctrl[13][28] , 
	\sa_ctrl[13][27] , \sa_ctrl[13][26] , \sa_ctrl[13][25] , 
	\sa_ctrl[13][24] , \sa_ctrl[13][23] , \sa_ctrl[13][22] , 
	\sa_ctrl[13][21] , \sa_ctrl[13][20] , \sa_ctrl[13][19] , 
	\sa_ctrl[13][18] , \sa_ctrl[13][17] , \sa_ctrl[13][16] , 
	\sa_ctrl[13][15] , \sa_ctrl[13][14] , \sa_ctrl[13][13] , 
	\sa_ctrl[13][12] , \sa_ctrl[13][11] , \sa_ctrl[13][10] , 
	\sa_ctrl[13][9] , \sa_ctrl[13][8] , \sa_ctrl[13][7] , 
	\sa_ctrl[13][6] , \sa_ctrl[13][5] , \sa_ctrl[13][4] , 
	\sa_ctrl[13][3] , \sa_ctrl[13][2] , \sa_ctrl[13][1] , 
	\sa_ctrl[13][0] , \sa_ctrl[12][31] , \sa_ctrl[12][30] , 
	\sa_ctrl[12][29] , \sa_ctrl[12][28] , \sa_ctrl[12][27] , 
	\sa_ctrl[12][26] , \sa_ctrl[12][25] , \sa_ctrl[12][24] , 
	\sa_ctrl[12][23] , \sa_ctrl[12][22] , \sa_ctrl[12][21] , 
	\sa_ctrl[12][20] , \sa_ctrl[12][19] , \sa_ctrl[12][18] , 
	\sa_ctrl[12][17] , \sa_ctrl[12][16] , \sa_ctrl[12][15] , 
	\sa_ctrl[12][14] , \sa_ctrl[12][13] , \sa_ctrl[12][12] , 
	\sa_ctrl[12][11] , \sa_ctrl[12][10] , \sa_ctrl[12][9] , 
	\sa_ctrl[12][8] , \sa_ctrl[12][7] , \sa_ctrl[12][6] , 
	\sa_ctrl[12][5] , \sa_ctrl[12][4] , \sa_ctrl[12][3] , 
	\sa_ctrl[12][2] , \sa_ctrl[12][1] , \sa_ctrl[12][0] , 
	\sa_ctrl[11][31] , \sa_ctrl[11][30] , \sa_ctrl[11][29] , 
	\sa_ctrl[11][28] , \sa_ctrl[11][27] , \sa_ctrl[11][26] , 
	\sa_ctrl[11][25] , \sa_ctrl[11][24] , \sa_ctrl[11][23] , 
	\sa_ctrl[11][22] , \sa_ctrl[11][21] , \sa_ctrl[11][20] , 
	\sa_ctrl[11][19] , \sa_ctrl[11][18] , \sa_ctrl[11][17] , 
	\sa_ctrl[11][16] , \sa_ctrl[11][15] , \sa_ctrl[11][14] , 
	\sa_ctrl[11][13] , \sa_ctrl[11][12] , \sa_ctrl[11][11] , 
	\sa_ctrl[11][10] , \sa_ctrl[11][9] , \sa_ctrl[11][8] , 
	\sa_ctrl[11][7] , \sa_ctrl[11][6] , \sa_ctrl[11][5] , 
	\sa_ctrl[11][4] , \sa_ctrl[11][3] , \sa_ctrl[11][2] , 
	\sa_ctrl[11][1] , \sa_ctrl[11][0] , \sa_ctrl[10][31] , 
	\sa_ctrl[10][30] , \sa_ctrl[10][29] , \sa_ctrl[10][28] , 
	\sa_ctrl[10][27] , \sa_ctrl[10][26] , \sa_ctrl[10][25] , 
	\sa_ctrl[10][24] , \sa_ctrl[10][23] , \sa_ctrl[10][22] , 
	\sa_ctrl[10][21] , \sa_ctrl[10][20] , \sa_ctrl[10][19] , 
	\sa_ctrl[10][18] , \sa_ctrl[10][17] , \sa_ctrl[10][16] , 
	\sa_ctrl[10][15] , \sa_ctrl[10][14] , \sa_ctrl[10][13] , 
	\sa_ctrl[10][12] , \sa_ctrl[10][11] , \sa_ctrl[10][10] , 
	\sa_ctrl[10][9] , \sa_ctrl[10][8] , \sa_ctrl[10][7] , 
	\sa_ctrl[10][6] , \sa_ctrl[10][5] , \sa_ctrl[10][4] , 
	\sa_ctrl[10][3] , \sa_ctrl[10][2] , \sa_ctrl[10][1] , 
	\sa_ctrl[10][0] , \sa_ctrl[9][31] , \sa_ctrl[9][30] , 
	\sa_ctrl[9][29] , \sa_ctrl[9][28] , \sa_ctrl[9][27] , 
	\sa_ctrl[9][26] , \sa_ctrl[9][25] , \sa_ctrl[9][24] , 
	\sa_ctrl[9][23] , \sa_ctrl[9][22] , \sa_ctrl[9][21] , 
	\sa_ctrl[9][20] , \sa_ctrl[9][19] , \sa_ctrl[9][18] , 
	\sa_ctrl[9][17] , \sa_ctrl[9][16] , \sa_ctrl[9][15] , 
	\sa_ctrl[9][14] , \sa_ctrl[9][13] , \sa_ctrl[9][12] , 
	\sa_ctrl[9][11] , \sa_ctrl[9][10] , \sa_ctrl[9][9] , \sa_ctrl[9][8] , 
	\sa_ctrl[9][7] , \sa_ctrl[9][6] , \sa_ctrl[9][5] , \sa_ctrl[9][4] , 
	\sa_ctrl[9][3] , \sa_ctrl[9][2] , \sa_ctrl[9][1] , \sa_ctrl[9][0] , 
	\sa_ctrl[8][31] , \sa_ctrl[8][30] , \sa_ctrl[8][29] , 
	\sa_ctrl[8][28] , \sa_ctrl[8][27] , \sa_ctrl[8][26] , 
	\sa_ctrl[8][25] , \sa_ctrl[8][24] , \sa_ctrl[8][23] , 
	\sa_ctrl[8][22] , \sa_ctrl[8][21] , \sa_ctrl[8][20] , 
	\sa_ctrl[8][19] , \sa_ctrl[8][18] , \sa_ctrl[8][17] , 
	\sa_ctrl[8][16] , \sa_ctrl[8][15] , \sa_ctrl[8][14] , 
	\sa_ctrl[8][13] , \sa_ctrl[8][12] , \sa_ctrl[8][11] , 
	\sa_ctrl[8][10] , \sa_ctrl[8][9] , \sa_ctrl[8][8] , \sa_ctrl[8][7] , 
	\sa_ctrl[8][6] , \sa_ctrl[8][5] , \sa_ctrl[8][4] , \sa_ctrl[8][3] , 
	\sa_ctrl[8][2] , \sa_ctrl[8][1] , \sa_ctrl[8][0] , \sa_ctrl[7][31] , 
	\sa_ctrl[7][30] , \sa_ctrl[7][29] , \sa_ctrl[7][28] , 
	\sa_ctrl[7][27] , \sa_ctrl[7][26] , \sa_ctrl[7][25] , 
	\sa_ctrl[7][24] , \sa_ctrl[7][23] , \sa_ctrl[7][22] , 
	\sa_ctrl[7][21] , \sa_ctrl[7][20] , \sa_ctrl[7][19] , 
	\sa_ctrl[7][18] , \sa_ctrl[7][17] , \sa_ctrl[7][16] , 
	\sa_ctrl[7][15] , \sa_ctrl[7][14] , \sa_ctrl[7][13] , 
	\sa_ctrl[7][12] , \sa_ctrl[7][11] , \sa_ctrl[7][10] , 
	\sa_ctrl[7][9] , \sa_ctrl[7][8] , \sa_ctrl[7][7] , \sa_ctrl[7][6] , 
	\sa_ctrl[7][5] , \sa_ctrl[7][4] , \sa_ctrl[7][3] , \sa_ctrl[7][2] , 
	\sa_ctrl[7][1] , \sa_ctrl[7][0] , \sa_ctrl[6][31] , \sa_ctrl[6][30] , 
	\sa_ctrl[6][29] , \sa_ctrl[6][28] , \sa_ctrl[6][27] , 
	\sa_ctrl[6][26] , \sa_ctrl[6][25] , \sa_ctrl[6][24] , 
	\sa_ctrl[6][23] , \sa_ctrl[6][22] , \sa_ctrl[6][21] , 
	\sa_ctrl[6][20] , \sa_ctrl[6][19] , \sa_ctrl[6][18] , 
	\sa_ctrl[6][17] , \sa_ctrl[6][16] , \sa_ctrl[6][15] , 
	\sa_ctrl[6][14] , \sa_ctrl[6][13] , \sa_ctrl[6][12] , 
	\sa_ctrl[6][11] , \sa_ctrl[6][10] , \sa_ctrl[6][9] , \sa_ctrl[6][8] , 
	\sa_ctrl[6][7] , \sa_ctrl[6][6] , \sa_ctrl[6][5] , \sa_ctrl[6][4] , 
	\sa_ctrl[6][3] , \sa_ctrl[6][2] , \sa_ctrl[6][1] , \sa_ctrl[6][0] , 
	\sa_ctrl[5][31] , \sa_ctrl[5][30] , \sa_ctrl[5][29] , 
	\sa_ctrl[5][28] , \sa_ctrl[5][27] , \sa_ctrl[5][26] , 
	\sa_ctrl[5][25] , \sa_ctrl[5][24] , \sa_ctrl[5][23] , 
	\sa_ctrl[5][22] , \sa_ctrl[5][21] , \sa_ctrl[5][20] , 
	\sa_ctrl[5][19] , \sa_ctrl[5][18] , \sa_ctrl[5][17] , 
	\sa_ctrl[5][16] , \sa_ctrl[5][15] , \sa_ctrl[5][14] , 
	\sa_ctrl[5][13] , \sa_ctrl[5][12] , \sa_ctrl[5][11] , 
	\sa_ctrl[5][10] , \sa_ctrl[5][9] , \sa_ctrl[5][8] , \sa_ctrl[5][7] , 
	\sa_ctrl[5][6] , \sa_ctrl[5][5] , \sa_ctrl[5][4] , \sa_ctrl[5][3] , 
	\sa_ctrl[5][2] , \sa_ctrl[5][1] , \sa_ctrl[5][0] , \sa_ctrl[4][31] , 
	\sa_ctrl[4][30] , \sa_ctrl[4][29] , \sa_ctrl[4][28] , 
	\sa_ctrl[4][27] , \sa_ctrl[4][26] , \sa_ctrl[4][25] , 
	\sa_ctrl[4][24] , \sa_ctrl[4][23] , \sa_ctrl[4][22] , 
	\sa_ctrl[4][21] , \sa_ctrl[4][20] , \sa_ctrl[4][19] , 
	\sa_ctrl[4][18] , \sa_ctrl[4][17] , \sa_ctrl[4][16] , 
	\sa_ctrl[4][15] , \sa_ctrl[4][14] , \sa_ctrl[4][13] , 
	\sa_ctrl[4][12] , \sa_ctrl[4][11] , \sa_ctrl[4][10] , 
	\sa_ctrl[4][9] , \sa_ctrl[4][8] , \sa_ctrl[4][7] , \sa_ctrl[4][6] , 
	\sa_ctrl[4][5] , \sa_ctrl[4][4] , \sa_ctrl[4][3] , \sa_ctrl[4][2] , 
	\sa_ctrl[4][1] , \sa_ctrl[4][0] , \sa_ctrl[3][31] , \sa_ctrl[3][30] , 
	\sa_ctrl[3][29] , \sa_ctrl[3][28] , \sa_ctrl[3][27] , 
	\sa_ctrl[3][26] , \sa_ctrl[3][25] , \sa_ctrl[3][24] , 
	\sa_ctrl[3][23] , \sa_ctrl[3][22] , \sa_ctrl[3][21] , 
	\sa_ctrl[3][20] , \sa_ctrl[3][19] , \sa_ctrl[3][18] , 
	\sa_ctrl[3][17] , \sa_ctrl[3][16] , \sa_ctrl[3][15] , 
	\sa_ctrl[3][14] , \sa_ctrl[3][13] , \sa_ctrl[3][12] , 
	\sa_ctrl[3][11] , \sa_ctrl[3][10] , \sa_ctrl[3][9] , \sa_ctrl[3][8] , 
	\sa_ctrl[3][7] , \sa_ctrl[3][6] , \sa_ctrl[3][5] , \sa_ctrl[3][4] , 
	\sa_ctrl[3][3] , \sa_ctrl[3][2] , \sa_ctrl[3][1] , \sa_ctrl[3][0] , 
	\sa_ctrl[2][31] , \sa_ctrl[2][30] , \sa_ctrl[2][29] , 
	\sa_ctrl[2][28] , \sa_ctrl[2][27] , \sa_ctrl[2][26] , 
	\sa_ctrl[2][25] , \sa_ctrl[2][24] , \sa_ctrl[2][23] , 
	\sa_ctrl[2][22] , \sa_ctrl[2][21] , \sa_ctrl[2][20] , 
	\sa_ctrl[2][19] , \sa_ctrl[2][18] , \sa_ctrl[2][17] , 
	\sa_ctrl[2][16] , \sa_ctrl[2][15] , \sa_ctrl[2][14] , 
	\sa_ctrl[2][13] , \sa_ctrl[2][12] , \sa_ctrl[2][11] , 
	\sa_ctrl[2][10] , \sa_ctrl[2][9] , \sa_ctrl[2][8] , \sa_ctrl[2][7] , 
	\sa_ctrl[2][6] , \sa_ctrl[2][5] , \sa_ctrl[2][4] , \sa_ctrl[2][3] , 
	\sa_ctrl[2][2] , \sa_ctrl[2][1] , \sa_ctrl[2][0] , \sa_ctrl[1][31] , 
	\sa_ctrl[1][30] , \sa_ctrl[1][29] , \sa_ctrl[1][28] , 
	\sa_ctrl[1][27] , \sa_ctrl[1][26] , \sa_ctrl[1][25] , 
	\sa_ctrl[1][24] , \sa_ctrl[1][23] , \sa_ctrl[1][22] , 
	\sa_ctrl[1][21] , \sa_ctrl[1][20] , \sa_ctrl[1][19] , 
	\sa_ctrl[1][18] , \sa_ctrl[1][17] , \sa_ctrl[1][16] , 
	\sa_ctrl[1][15] , \sa_ctrl[1][14] , \sa_ctrl[1][13] , 
	\sa_ctrl[1][12] , \sa_ctrl[1][11] , \sa_ctrl[1][10] , 
	\sa_ctrl[1][9] , \sa_ctrl[1][8] , \sa_ctrl[1][7] , \sa_ctrl[1][6] , 
	\sa_ctrl[1][5] , \sa_ctrl[1][4] , \sa_ctrl[1][3] , \sa_ctrl[1][2] , 
	\sa_ctrl[1][1] , \sa_ctrl[1][0] , \sa_ctrl[0][31] , \sa_ctrl[0][30] , 
	\sa_ctrl[0][29] , \sa_ctrl[0][28] , \sa_ctrl[0][27] , 
	\sa_ctrl[0][26] , \sa_ctrl[0][25] , \sa_ctrl[0][24] , 
	\sa_ctrl[0][23] , \sa_ctrl[0][22] , \sa_ctrl[0][21] , 
	\sa_ctrl[0][20] , \sa_ctrl[0][19] , \sa_ctrl[0][18] , 
	\sa_ctrl[0][17] , \sa_ctrl[0][16] , \sa_ctrl[0][15] , 
	\sa_ctrl[0][14] , \sa_ctrl[0][13] , \sa_ctrl[0][12] , 
	\sa_ctrl[0][11] , \sa_ctrl[0][10] , \sa_ctrl[0][9] , \sa_ctrl[0][8] , 
	\sa_ctrl[0][7] , \sa_ctrl[0][6] , \sa_ctrl[0][5] , \sa_ctrl[0][4] , 
	\sa_ctrl[0][3] , \sa_ctrl[0][2] , \sa_ctrl[0][1] , \sa_ctrl[0][0] }), 
	.clk( clk), .rst_n( rst_n), .addr( 
	_zy_simnet_reg_addr_800_w$[0:10]), .cmnd_op( 
	_zy_simnet_sa_ctrl_ia_config_801_w$[0:3]), .cmnd_addr( 
	_zy_simnet_sa_ctrl_ia_config_802_w$[0:4]), .wr_stb( 
	_zy_simnet_wr_stb_803_w$), .wr_dat( 
	_zy_simnet_sa_ctrl_ia_wdata_804_w$[0:31]), .rst_dat( { 
	\sa_ctrl_rst_dat[31][31] , \sa_ctrl_rst_dat[31][30] , 
	\sa_ctrl_rst_dat[31][29] , \sa_ctrl_rst_dat[31][28] , 
	\sa_ctrl_rst_dat[31][27] , \sa_ctrl_rst_dat[31][26] , 
	\sa_ctrl_rst_dat[31][25] , \sa_ctrl_rst_dat[31][24] , 
	\sa_ctrl_rst_dat[31][23] , \sa_ctrl_rst_dat[31][22] , 
	\sa_ctrl_rst_dat[31][21] , \sa_ctrl_rst_dat[31][20] , 
	\sa_ctrl_rst_dat[31][19] , \sa_ctrl_rst_dat[31][18] , 
	\sa_ctrl_rst_dat[31][17] , \sa_ctrl_rst_dat[31][16] , 
	\sa_ctrl_rst_dat[31][15] , \sa_ctrl_rst_dat[31][14] , 
	\sa_ctrl_rst_dat[31][13] , \sa_ctrl_rst_dat[31][12] , 
	\sa_ctrl_rst_dat[31][11] , \sa_ctrl_rst_dat[31][10] , 
	\sa_ctrl_rst_dat[31][9] , \sa_ctrl_rst_dat[31][8] , 
	\sa_ctrl_rst_dat[31][7] , \sa_ctrl_rst_dat[31][6] , 
	\sa_ctrl_rst_dat[31][5] , \sa_ctrl_rst_dat[31][4] , 
	\sa_ctrl_rst_dat[31][3] , \sa_ctrl_rst_dat[31][2] , 
	\sa_ctrl_rst_dat[31][1] , \sa_ctrl_rst_dat[31][0] , 
	\sa_ctrl_rst_dat[30][31] , \sa_ctrl_rst_dat[30][30] , 
	\sa_ctrl_rst_dat[30][29] , \sa_ctrl_rst_dat[30][28] , 
	\sa_ctrl_rst_dat[30][27] , \sa_ctrl_rst_dat[30][26] , 
	\sa_ctrl_rst_dat[30][25] , \sa_ctrl_rst_dat[30][24] , 
	\sa_ctrl_rst_dat[30][23] , \sa_ctrl_rst_dat[30][22] , 
	\sa_ctrl_rst_dat[30][21] , \sa_ctrl_rst_dat[30][20] , 
	\sa_ctrl_rst_dat[30][19] , \sa_ctrl_rst_dat[30][18] , 
	\sa_ctrl_rst_dat[30][17] , \sa_ctrl_rst_dat[30][16] , 
	\sa_ctrl_rst_dat[30][15] , \sa_ctrl_rst_dat[30][14] , 
	\sa_ctrl_rst_dat[30][13] , \sa_ctrl_rst_dat[30][12] , 
	\sa_ctrl_rst_dat[30][11] , \sa_ctrl_rst_dat[30][10] , 
	\sa_ctrl_rst_dat[30][9] , \sa_ctrl_rst_dat[30][8] , 
	\sa_ctrl_rst_dat[30][7] , \sa_ctrl_rst_dat[30][6] , 
	\sa_ctrl_rst_dat[30][5] , \sa_ctrl_rst_dat[30][4] , 
	\sa_ctrl_rst_dat[30][3] , \sa_ctrl_rst_dat[30][2] , 
	\sa_ctrl_rst_dat[30][1] , \sa_ctrl_rst_dat[30][0] , 
	\sa_ctrl_rst_dat[29][31] , \sa_ctrl_rst_dat[29][30] , 
	\sa_ctrl_rst_dat[29][29] , \sa_ctrl_rst_dat[29][28] , 
	\sa_ctrl_rst_dat[29][27] , \sa_ctrl_rst_dat[29][26] , 
	\sa_ctrl_rst_dat[29][25] , \sa_ctrl_rst_dat[29][24] , 
	\sa_ctrl_rst_dat[29][23] , \sa_ctrl_rst_dat[29][22] , 
	\sa_ctrl_rst_dat[29][21] , \sa_ctrl_rst_dat[29][20] , 
	\sa_ctrl_rst_dat[29][19] , \sa_ctrl_rst_dat[29][18] , 
	\sa_ctrl_rst_dat[29][17] , \sa_ctrl_rst_dat[29][16] , 
	\sa_ctrl_rst_dat[29][15] , \sa_ctrl_rst_dat[29][14] , 
	\sa_ctrl_rst_dat[29][13] , \sa_ctrl_rst_dat[29][12] , 
	\sa_ctrl_rst_dat[29][11] , \sa_ctrl_rst_dat[29][10] , 
	\sa_ctrl_rst_dat[29][9] , \sa_ctrl_rst_dat[29][8] , 
	\sa_ctrl_rst_dat[29][7] , \sa_ctrl_rst_dat[29][6] , 
	\sa_ctrl_rst_dat[29][5] , \sa_ctrl_rst_dat[29][4] , 
	\sa_ctrl_rst_dat[29][3] , \sa_ctrl_rst_dat[29][2] , 
	\sa_ctrl_rst_dat[29][1] , \sa_ctrl_rst_dat[29][0] , 
	\sa_ctrl_rst_dat[28][31] , \sa_ctrl_rst_dat[28][30] , 
	\sa_ctrl_rst_dat[28][29] , \sa_ctrl_rst_dat[28][28] , 
	\sa_ctrl_rst_dat[28][27] , \sa_ctrl_rst_dat[28][26] , 
	\sa_ctrl_rst_dat[28][25] , \sa_ctrl_rst_dat[28][24] , 
	\sa_ctrl_rst_dat[28][23] , \sa_ctrl_rst_dat[28][22] , 
	\sa_ctrl_rst_dat[28][21] , \sa_ctrl_rst_dat[28][20] , 
	\sa_ctrl_rst_dat[28][19] , \sa_ctrl_rst_dat[28][18] , 
	\sa_ctrl_rst_dat[28][17] , \sa_ctrl_rst_dat[28][16] , 
	\sa_ctrl_rst_dat[28][15] , \sa_ctrl_rst_dat[28][14] , 
	\sa_ctrl_rst_dat[28][13] , \sa_ctrl_rst_dat[28][12] , 
	\sa_ctrl_rst_dat[28][11] , \sa_ctrl_rst_dat[28][10] , 
	\sa_ctrl_rst_dat[28][9] , \sa_ctrl_rst_dat[28][8] , 
	\sa_ctrl_rst_dat[28][7] , \sa_ctrl_rst_dat[28][6] , 
	\sa_ctrl_rst_dat[28][5] , \sa_ctrl_rst_dat[28][4] , 
	\sa_ctrl_rst_dat[28][3] , \sa_ctrl_rst_dat[28][2] , 
	\sa_ctrl_rst_dat[28][1] , \sa_ctrl_rst_dat[28][0] , 
	\sa_ctrl_rst_dat[27][31] , \sa_ctrl_rst_dat[27][30] , 
	\sa_ctrl_rst_dat[27][29] , \sa_ctrl_rst_dat[27][28] , 
	\sa_ctrl_rst_dat[27][27] , \sa_ctrl_rst_dat[27][26] , 
	\sa_ctrl_rst_dat[27][25] , \sa_ctrl_rst_dat[27][24] , 
	\sa_ctrl_rst_dat[27][23] , \sa_ctrl_rst_dat[27][22] , 
	\sa_ctrl_rst_dat[27][21] , \sa_ctrl_rst_dat[27][20] , 
	\sa_ctrl_rst_dat[27][19] , \sa_ctrl_rst_dat[27][18] , 
	\sa_ctrl_rst_dat[27][17] , \sa_ctrl_rst_dat[27][16] , 
	\sa_ctrl_rst_dat[27][15] , \sa_ctrl_rst_dat[27][14] , 
	\sa_ctrl_rst_dat[27][13] , \sa_ctrl_rst_dat[27][12] , 
	\sa_ctrl_rst_dat[27][11] , \sa_ctrl_rst_dat[27][10] , 
	\sa_ctrl_rst_dat[27][9] , \sa_ctrl_rst_dat[27][8] , 
	\sa_ctrl_rst_dat[27][7] , \sa_ctrl_rst_dat[27][6] , 
	\sa_ctrl_rst_dat[27][5] , \sa_ctrl_rst_dat[27][4] , 
	\sa_ctrl_rst_dat[27][3] , \sa_ctrl_rst_dat[27][2] , 
	\sa_ctrl_rst_dat[27][1] , \sa_ctrl_rst_dat[27][0] , 
	\sa_ctrl_rst_dat[26][31] , \sa_ctrl_rst_dat[26][30] , 
	\sa_ctrl_rst_dat[26][29] , \sa_ctrl_rst_dat[26][28] , 
	\sa_ctrl_rst_dat[26][27] , \sa_ctrl_rst_dat[26][26] , 
	\sa_ctrl_rst_dat[26][25] , \sa_ctrl_rst_dat[26][24] , 
	\sa_ctrl_rst_dat[26][23] , \sa_ctrl_rst_dat[26][22] , 
	\sa_ctrl_rst_dat[26][21] , \sa_ctrl_rst_dat[26][20] , 
	\sa_ctrl_rst_dat[26][19] , \sa_ctrl_rst_dat[26][18] , 
	\sa_ctrl_rst_dat[26][17] , \sa_ctrl_rst_dat[26][16] , 
	\sa_ctrl_rst_dat[26][15] , \sa_ctrl_rst_dat[26][14] , 
	\sa_ctrl_rst_dat[26][13] , \sa_ctrl_rst_dat[26][12] , 
	\sa_ctrl_rst_dat[26][11] , \sa_ctrl_rst_dat[26][10] , 
	\sa_ctrl_rst_dat[26][9] , \sa_ctrl_rst_dat[26][8] , 
	\sa_ctrl_rst_dat[26][7] , \sa_ctrl_rst_dat[26][6] , 
	\sa_ctrl_rst_dat[26][5] , \sa_ctrl_rst_dat[26][4] , 
	\sa_ctrl_rst_dat[26][3] , \sa_ctrl_rst_dat[26][2] , 
	\sa_ctrl_rst_dat[26][1] , \sa_ctrl_rst_dat[26][0] , 
	\sa_ctrl_rst_dat[25][31] , \sa_ctrl_rst_dat[25][30] , 
	\sa_ctrl_rst_dat[25][29] , \sa_ctrl_rst_dat[25][28] , 
	\sa_ctrl_rst_dat[25][27] , \sa_ctrl_rst_dat[25][26] , 
	\sa_ctrl_rst_dat[25][25] , \sa_ctrl_rst_dat[25][24] , 
	\sa_ctrl_rst_dat[25][23] , \sa_ctrl_rst_dat[25][22] , 
	\sa_ctrl_rst_dat[25][21] , \sa_ctrl_rst_dat[25][20] , 
	\sa_ctrl_rst_dat[25][19] , \sa_ctrl_rst_dat[25][18] , 
	\sa_ctrl_rst_dat[25][17] , \sa_ctrl_rst_dat[25][16] , 
	\sa_ctrl_rst_dat[25][15] , \sa_ctrl_rst_dat[25][14] , 
	\sa_ctrl_rst_dat[25][13] , \sa_ctrl_rst_dat[25][12] , 
	\sa_ctrl_rst_dat[25][11] , \sa_ctrl_rst_dat[25][10] , 
	\sa_ctrl_rst_dat[25][9] , \sa_ctrl_rst_dat[25][8] , 
	\sa_ctrl_rst_dat[25][7] , \sa_ctrl_rst_dat[25][6] , 
	\sa_ctrl_rst_dat[25][5] , \sa_ctrl_rst_dat[25][4] , 
	\sa_ctrl_rst_dat[25][3] , \sa_ctrl_rst_dat[25][2] , 
	\sa_ctrl_rst_dat[25][1] , \sa_ctrl_rst_dat[25][0] , 
	\sa_ctrl_rst_dat[24][31] , \sa_ctrl_rst_dat[24][30] , 
	\sa_ctrl_rst_dat[24][29] , \sa_ctrl_rst_dat[24][28] , 
	\sa_ctrl_rst_dat[24][27] , \sa_ctrl_rst_dat[24][26] , 
	\sa_ctrl_rst_dat[24][25] , \sa_ctrl_rst_dat[24][24] , 
	\sa_ctrl_rst_dat[24][23] , \sa_ctrl_rst_dat[24][22] , 
	\sa_ctrl_rst_dat[24][21] , \sa_ctrl_rst_dat[24][20] , 
	\sa_ctrl_rst_dat[24][19] , \sa_ctrl_rst_dat[24][18] , 
	\sa_ctrl_rst_dat[24][17] , \sa_ctrl_rst_dat[24][16] , 
	\sa_ctrl_rst_dat[24][15] , \sa_ctrl_rst_dat[24][14] , 
	\sa_ctrl_rst_dat[24][13] , \sa_ctrl_rst_dat[24][12] , 
	\sa_ctrl_rst_dat[24][11] , \sa_ctrl_rst_dat[24][10] , 
	\sa_ctrl_rst_dat[24][9] , \sa_ctrl_rst_dat[24][8] , 
	\sa_ctrl_rst_dat[24][7] , \sa_ctrl_rst_dat[24][6] , 
	\sa_ctrl_rst_dat[24][5] , \sa_ctrl_rst_dat[24][4] , 
	\sa_ctrl_rst_dat[24][3] , \sa_ctrl_rst_dat[24][2] , 
	\sa_ctrl_rst_dat[24][1] , \sa_ctrl_rst_dat[24][0] , 
	\sa_ctrl_rst_dat[23][31] , \sa_ctrl_rst_dat[23][30] , 
	\sa_ctrl_rst_dat[23][29] , \sa_ctrl_rst_dat[23][28] , 
	\sa_ctrl_rst_dat[23][27] , \sa_ctrl_rst_dat[23][26] , 
	\sa_ctrl_rst_dat[23][25] , \sa_ctrl_rst_dat[23][24] , 
	\sa_ctrl_rst_dat[23][23] , \sa_ctrl_rst_dat[23][22] , 
	\sa_ctrl_rst_dat[23][21] , \sa_ctrl_rst_dat[23][20] , 
	\sa_ctrl_rst_dat[23][19] , \sa_ctrl_rst_dat[23][18] , 
	\sa_ctrl_rst_dat[23][17] , \sa_ctrl_rst_dat[23][16] , 
	\sa_ctrl_rst_dat[23][15] , \sa_ctrl_rst_dat[23][14] , 
	\sa_ctrl_rst_dat[23][13] , \sa_ctrl_rst_dat[23][12] , 
	\sa_ctrl_rst_dat[23][11] , \sa_ctrl_rst_dat[23][10] , 
	\sa_ctrl_rst_dat[23][9] , \sa_ctrl_rst_dat[23][8] , 
	\sa_ctrl_rst_dat[23][7] , \sa_ctrl_rst_dat[23][6] , 
	\sa_ctrl_rst_dat[23][5] , \sa_ctrl_rst_dat[23][4] , 
	\sa_ctrl_rst_dat[23][3] , \sa_ctrl_rst_dat[23][2] , 
	\sa_ctrl_rst_dat[23][1] , \sa_ctrl_rst_dat[23][0] , 
	\sa_ctrl_rst_dat[22][31] , \sa_ctrl_rst_dat[22][30] , 
	\sa_ctrl_rst_dat[22][29] , \sa_ctrl_rst_dat[22][28] , 
	\sa_ctrl_rst_dat[22][27] , \sa_ctrl_rst_dat[22][26] , 
	\sa_ctrl_rst_dat[22][25] , \sa_ctrl_rst_dat[22][24] , 
	\sa_ctrl_rst_dat[22][23] , \sa_ctrl_rst_dat[22][22] , 
	\sa_ctrl_rst_dat[22][21] , \sa_ctrl_rst_dat[22][20] , 
	\sa_ctrl_rst_dat[22][19] , \sa_ctrl_rst_dat[22][18] , 
	\sa_ctrl_rst_dat[22][17] , \sa_ctrl_rst_dat[22][16] , 
	\sa_ctrl_rst_dat[22][15] , \sa_ctrl_rst_dat[22][14] , 
	\sa_ctrl_rst_dat[22][13] , \sa_ctrl_rst_dat[22][12] , 
	\sa_ctrl_rst_dat[22][11] , \sa_ctrl_rst_dat[22][10] , 
	\sa_ctrl_rst_dat[22][9] , \sa_ctrl_rst_dat[22][8] , 
	\sa_ctrl_rst_dat[22][7] , \sa_ctrl_rst_dat[22][6] , 
	\sa_ctrl_rst_dat[22][5] , \sa_ctrl_rst_dat[22][4] , 
	\sa_ctrl_rst_dat[22][3] , \sa_ctrl_rst_dat[22][2] , 
	\sa_ctrl_rst_dat[22][1] , \sa_ctrl_rst_dat[22][0] , 
	\sa_ctrl_rst_dat[21][31] , \sa_ctrl_rst_dat[21][30] , 
	\sa_ctrl_rst_dat[21][29] , \sa_ctrl_rst_dat[21][28] , 
	\sa_ctrl_rst_dat[21][27] , \sa_ctrl_rst_dat[21][26] , 
	\sa_ctrl_rst_dat[21][25] , \sa_ctrl_rst_dat[21][24] , 
	\sa_ctrl_rst_dat[21][23] , \sa_ctrl_rst_dat[21][22] , 
	\sa_ctrl_rst_dat[21][21] , \sa_ctrl_rst_dat[21][20] , 
	\sa_ctrl_rst_dat[21][19] , \sa_ctrl_rst_dat[21][18] , 
	\sa_ctrl_rst_dat[21][17] , \sa_ctrl_rst_dat[21][16] , 
	\sa_ctrl_rst_dat[21][15] , \sa_ctrl_rst_dat[21][14] , 
	\sa_ctrl_rst_dat[21][13] , \sa_ctrl_rst_dat[21][12] , 
	\sa_ctrl_rst_dat[21][11] , \sa_ctrl_rst_dat[21][10] , 
	\sa_ctrl_rst_dat[21][9] , \sa_ctrl_rst_dat[21][8] , 
	\sa_ctrl_rst_dat[21][7] , \sa_ctrl_rst_dat[21][6] , 
	\sa_ctrl_rst_dat[21][5] , \sa_ctrl_rst_dat[21][4] , 
	\sa_ctrl_rst_dat[21][3] , \sa_ctrl_rst_dat[21][2] , 
	\sa_ctrl_rst_dat[21][1] , \sa_ctrl_rst_dat[21][0] , 
	\sa_ctrl_rst_dat[20][31] , \sa_ctrl_rst_dat[20][30] , 
	\sa_ctrl_rst_dat[20][29] , \sa_ctrl_rst_dat[20][28] , 
	\sa_ctrl_rst_dat[20][27] , \sa_ctrl_rst_dat[20][26] , 
	\sa_ctrl_rst_dat[20][25] , \sa_ctrl_rst_dat[20][24] , 
	\sa_ctrl_rst_dat[20][23] , \sa_ctrl_rst_dat[20][22] , 
	\sa_ctrl_rst_dat[20][21] , \sa_ctrl_rst_dat[20][20] , 
	\sa_ctrl_rst_dat[20][19] , \sa_ctrl_rst_dat[20][18] , 
	\sa_ctrl_rst_dat[20][17] , \sa_ctrl_rst_dat[20][16] , 
	\sa_ctrl_rst_dat[20][15] , \sa_ctrl_rst_dat[20][14] , 
	\sa_ctrl_rst_dat[20][13] , \sa_ctrl_rst_dat[20][12] , 
	\sa_ctrl_rst_dat[20][11] , \sa_ctrl_rst_dat[20][10] , 
	\sa_ctrl_rst_dat[20][9] , \sa_ctrl_rst_dat[20][8] , 
	\sa_ctrl_rst_dat[20][7] , \sa_ctrl_rst_dat[20][6] , 
	\sa_ctrl_rst_dat[20][5] , \sa_ctrl_rst_dat[20][4] , 
	\sa_ctrl_rst_dat[20][3] , \sa_ctrl_rst_dat[20][2] , 
	\sa_ctrl_rst_dat[20][1] , \sa_ctrl_rst_dat[20][0] , 
	\sa_ctrl_rst_dat[19][31] , \sa_ctrl_rst_dat[19][30] , 
	\sa_ctrl_rst_dat[19][29] , \sa_ctrl_rst_dat[19][28] , 
	\sa_ctrl_rst_dat[19][27] , \sa_ctrl_rst_dat[19][26] , 
	\sa_ctrl_rst_dat[19][25] , \sa_ctrl_rst_dat[19][24] , 
	\sa_ctrl_rst_dat[19][23] , \sa_ctrl_rst_dat[19][22] , 
	\sa_ctrl_rst_dat[19][21] , \sa_ctrl_rst_dat[19][20] , 
	\sa_ctrl_rst_dat[19][19] , \sa_ctrl_rst_dat[19][18] , 
	\sa_ctrl_rst_dat[19][17] , \sa_ctrl_rst_dat[19][16] , 
	\sa_ctrl_rst_dat[19][15] , \sa_ctrl_rst_dat[19][14] , 
	\sa_ctrl_rst_dat[19][13] , \sa_ctrl_rst_dat[19][12] , 
	\sa_ctrl_rst_dat[19][11] , \sa_ctrl_rst_dat[19][10] , 
	\sa_ctrl_rst_dat[19][9] , \sa_ctrl_rst_dat[19][8] , 
	\sa_ctrl_rst_dat[19][7] , \sa_ctrl_rst_dat[19][6] , 
	\sa_ctrl_rst_dat[19][5] , \sa_ctrl_rst_dat[19][4] , 
	\sa_ctrl_rst_dat[19][3] , \sa_ctrl_rst_dat[19][2] , 
	\sa_ctrl_rst_dat[19][1] , \sa_ctrl_rst_dat[19][0] , 
	\sa_ctrl_rst_dat[18][31] , \sa_ctrl_rst_dat[18][30] , 
	\sa_ctrl_rst_dat[18][29] , \sa_ctrl_rst_dat[18][28] , 
	\sa_ctrl_rst_dat[18][27] , \sa_ctrl_rst_dat[18][26] , 
	\sa_ctrl_rst_dat[18][25] , \sa_ctrl_rst_dat[18][24] , 
	\sa_ctrl_rst_dat[18][23] , \sa_ctrl_rst_dat[18][22] , 
	\sa_ctrl_rst_dat[18][21] , \sa_ctrl_rst_dat[18][20] , 
	\sa_ctrl_rst_dat[18][19] , \sa_ctrl_rst_dat[18][18] , 
	\sa_ctrl_rst_dat[18][17] , \sa_ctrl_rst_dat[18][16] , 
	\sa_ctrl_rst_dat[18][15] , \sa_ctrl_rst_dat[18][14] , 
	\sa_ctrl_rst_dat[18][13] , \sa_ctrl_rst_dat[18][12] , 
	\sa_ctrl_rst_dat[18][11] , \sa_ctrl_rst_dat[18][10] , 
	\sa_ctrl_rst_dat[18][9] , \sa_ctrl_rst_dat[18][8] , 
	\sa_ctrl_rst_dat[18][7] , \sa_ctrl_rst_dat[18][6] , 
	\sa_ctrl_rst_dat[18][5] , \sa_ctrl_rst_dat[18][4] , 
	\sa_ctrl_rst_dat[18][3] , \sa_ctrl_rst_dat[18][2] , 
	\sa_ctrl_rst_dat[18][1] , \sa_ctrl_rst_dat[18][0] , 
	\sa_ctrl_rst_dat[17][31] , \sa_ctrl_rst_dat[17][30] , 
	\sa_ctrl_rst_dat[17][29] , \sa_ctrl_rst_dat[17][28] , 
	\sa_ctrl_rst_dat[17][27] , \sa_ctrl_rst_dat[17][26] , 
	\sa_ctrl_rst_dat[17][25] , \sa_ctrl_rst_dat[17][24] , 
	\sa_ctrl_rst_dat[17][23] , \sa_ctrl_rst_dat[17][22] , 
	\sa_ctrl_rst_dat[17][21] , \sa_ctrl_rst_dat[17][20] , 
	\sa_ctrl_rst_dat[17][19] , \sa_ctrl_rst_dat[17][18] , 
	\sa_ctrl_rst_dat[17][17] , \sa_ctrl_rst_dat[17][16] , 
	\sa_ctrl_rst_dat[17][15] , \sa_ctrl_rst_dat[17][14] , 
	\sa_ctrl_rst_dat[17][13] , \sa_ctrl_rst_dat[17][12] , 
	\sa_ctrl_rst_dat[17][11] , \sa_ctrl_rst_dat[17][10] , 
	\sa_ctrl_rst_dat[17][9] , \sa_ctrl_rst_dat[17][8] , 
	\sa_ctrl_rst_dat[17][7] , \sa_ctrl_rst_dat[17][6] , 
	\sa_ctrl_rst_dat[17][5] , \sa_ctrl_rst_dat[17][4] , 
	\sa_ctrl_rst_dat[17][3] , \sa_ctrl_rst_dat[17][2] , 
	\sa_ctrl_rst_dat[17][1] , \sa_ctrl_rst_dat[17][0] , 
	\sa_ctrl_rst_dat[16][31] , \sa_ctrl_rst_dat[16][30] , 
	\sa_ctrl_rst_dat[16][29] , \sa_ctrl_rst_dat[16][28] , 
	\sa_ctrl_rst_dat[16][27] , \sa_ctrl_rst_dat[16][26] , 
	\sa_ctrl_rst_dat[16][25] , \sa_ctrl_rst_dat[16][24] , 
	\sa_ctrl_rst_dat[16][23] , \sa_ctrl_rst_dat[16][22] , 
	\sa_ctrl_rst_dat[16][21] , \sa_ctrl_rst_dat[16][20] , 
	\sa_ctrl_rst_dat[16][19] , \sa_ctrl_rst_dat[16][18] , 
	\sa_ctrl_rst_dat[16][17] , \sa_ctrl_rst_dat[16][16] , 
	\sa_ctrl_rst_dat[16][15] , \sa_ctrl_rst_dat[16][14] , 
	\sa_ctrl_rst_dat[16][13] , \sa_ctrl_rst_dat[16][12] , 
	\sa_ctrl_rst_dat[16][11] , \sa_ctrl_rst_dat[16][10] , 
	\sa_ctrl_rst_dat[16][9] , \sa_ctrl_rst_dat[16][8] , 
	\sa_ctrl_rst_dat[16][7] , \sa_ctrl_rst_dat[16][6] , 
	\sa_ctrl_rst_dat[16][5] , \sa_ctrl_rst_dat[16][4] , 
	\sa_ctrl_rst_dat[16][3] , \sa_ctrl_rst_dat[16][2] , 
	\sa_ctrl_rst_dat[16][1] , \sa_ctrl_rst_dat[16][0] , 
	\sa_ctrl_rst_dat[15][31] , \sa_ctrl_rst_dat[15][30] , 
	\sa_ctrl_rst_dat[15][29] , \sa_ctrl_rst_dat[15][28] , 
	\sa_ctrl_rst_dat[15][27] , \sa_ctrl_rst_dat[15][26] , 
	\sa_ctrl_rst_dat[15][25] , \sa_ctrl_rst_dat[15][24] , 
	\sa_ctrl_rst_dat[15][23] , \sa_ctrl_rst_dat[15][22] , 
	\sa_ctrl_rst_dat[15][21] , \sa_ctrl_rst_dat[15][20] , 
	\sa_ctrl_rst_dat[15][19] , \sa_ctrl_rst_dat[15][18] , 
	\sa_ctrl_rst_dat[15][17] , \sa_ctrl_rst_dat[15][16] , 
	\sa_ctrl_rst_dat[15][15] , \sa_ctrl_rst_dat[15][14] , 
	\sa_ctrl_rst_dat[15][13] , \sa_ctrl_rst_dat[15][12] , 
	\sa_ctrl_rst_dat[15][11] , \sa_ctrl_rst_dat[15][10] , 
	\sa_ctrl_rst_dat[15][9] , \sa_ctrl_rst_dat[15][8] , 
	\sa_ctrl_rst_dat[15][7] , \sa_ctrl_rst_dat[15][6] , 
	\sa_ctrl_rst_dat[15][5] , \sa_ctrl_rst_dat[15][4] , 
	\sa_ctrl_rst_dat[15][3] , \sa_ctrl_rst_dat[15][2] , 
	\sa_ctrl_rst_dat[15][1] , \sa_ctrl_rst_dat[15][0] , 
	\sa_ctrl_rst_dat[14][31] , \sa_ctrl_rst_dat[14][30] , 
	\sa_ctrl_rst_dat[14][29] , \sa_ctrl_rst_dat[14][28] , 
	\sa_ctrl_rst_dat[14][27] , \sa_ctrl_rst_dat[14][26] , 
	\sa_ctrl_rst_dat[14][25] , \sa_ctrl_rst_dat[14][24] , 
	\sa_ctrl_rst_dat[14][23] , \sa_ctrl_rst_dat[14][22] , 
	\sa_ctrl_rst_dat[14][21] , \sa_ctrl_rst_dat[14][20] , 
	\sa_ctrl_rst_dat[14][19] , \sa_ctrl_rst_dat[14][18] , 
	\sa_ctrl_rst_dat[14][17] , \sa_ctrl_rst_dat[14][16] , 
	\sa_ctrl_rst_dat[14][15] , \sa_ctrl_rst_dat[14][14] , 
	\sa_ctrl_rst_dat[14][13] , \sa_ctrl_rst_dat[14][12] , 
	\sa_ctrl_rst_dat[14][11] , \sa_ctrl_rst_dat[14][10] , 
	\sa_ctrl_rst_dat[14][9] , \sa_ctrl_rst_dat[14][8] , 
	\sa_ctrl_rst_dat[14][7] , \sa_ctrl_rst_dat[14][6] , 
	\sa_ctrl_rst_dat[14][5] , \sa_ctrl_rst_dat[14][4] , 
	\sa_ctrl_rst_dat[14][3] , \sa_ctrl_rst_dat[14][2] , 
	\sa_ctrl_rst_dat[14][1] , \sa_ctrl_rst_dat[14][0] , 
	\sa_ctrl_rst_dat[13][31] , \sa_ctrl_rst_dat[13][30] , 
	\sa_ctrl_rst_dat[13][29] , \sa_ctrl_rst_dat[13][28] , 
	\sa_ctrl_rst_dat[13][27] , \sa_ctrl_rst_dat[13][26] , 
	\sa_ctrl_rst_dat[13][25] , \sa_ctrl_rst_dat[13][24] , 
	\sa_ctrl_rst_dat[13][23] , \sa_ctrl_rst_dat[13][22] , 
	\sa_ctrl_rst_dat[13][21] , \sa_ctrl_rst_dat[13][20] , 
	\sa_ctrl_rst_dat[13][19] , \sa_ctrl_rst_dat[13][18] , 
	\sa_ctrl_rst_dat[13][17] , \sa_ctrl_rst_dat[13][16] , 
	\sa_ctrl_rst_dat[13][15] , \sa_ctrl_rst_dat[13][14] , 
	\sa_ctrl_rst_dat[13][13] , \sa_ctrl_rst_dat[13][12] , 
	\sa_ctrl_rst_dat[13][11] , \sa_ctrl_rst_dat[13][10] , 
	\sa_ctrl_rst_dat[13][9] , \sa_ctrl_rst_dat[13][8] , 
	\sa_ctrl_rst_dat[13][7] , \sa_ctrl_rst_dat[13][6] , 
	\sa_ctrl_rst_dat[13][5] , \sa_ctrl_rst_dat[13][4] , 
	\sa_ctrl_rst_dat[13][3] , \sa_ctrl_rst_dat[13][2] , 
	\sa_ctrl_rst_dat[13][1] , \sa_ctrl_rst_dat[13][0] , 
	\sa_ctrl_rst_dat[12][31] , \sa_ctrl_rst_dat[12][30] , 
	\sa_ctrl_rst_dat[12][29] , \sa_ctrl_rst_dat[12][28] , 
	\sa_ctrl_rst_dat[12][27] , \sa_ctrl_rst_dat[12][26] , 
	\sa_ctrl_rst_dat[12][25] , \sa_ctrl_rst_dat[12][24] , 
	\sa_ctrl_rst_dat[12][23] , \sa_ctrl_rst_dat[12][22] , 
	\sa_ctrl_rst_dat[12][21] , \sa_ctrl_rst_dat[12][20] , 
	\sa_ctrl_rst_dat[12][19] , \sa_ctrl_rst_dat[12][18] , 
	\sa_ctrl_rst_dat[12][17] , \sa_ctrl_rst_dat[12][16] , 
	\sa_ctrl_rst_dat[12][15] , \sa_ctrl_rst_dat[12][14] , 
	\sa_ctrl_rst_dat[12][13] , \sa_ctrl_rst_dat[12][12] , 
	\sa_ctrl_rst_dat[12][11] , \sa_ctrl_rst_dat[12][10] , 
	\sa_ctrl_rst_dat[12][9] , \sa_ctrl_rst_dat[12][8] , 
	\sa_ctrl_rst_dat[12][7] , \sa_ctrl_rst_dat[12][6] , 
	\sa_ctrl_rst_dat[12][5] , \sa_ctrl_rst_dat[12][4] , 
	\sa_ctrl_rst_dat[12][3] , \sa_ctrl_rst_dat[12][2] , 
	\sa_ctrl_rst_dat[12][1] , \sa_ctrl_rst_dat[12][0] , 
	\sa_ctrl_rst_dat[11][31] , \sa_ctrl_rst_dat[11][30] , 
	\sa_ctrl_rst_dat[11][29] , \sa_ctrl_rst_dat[11][28] , 
	\sa_ctrl_rst_dat[11][27] , \sa_ctrl_rst_dat[11][26] , 
	\sa_ctrl_rst_dat[11][25] , \sa_ctrl_rst_dat[11][24] , 
	\sa_ctrl_rst_dat[11][23] , \sa_ctrl_rst_dat[11][22] , 
	\sa_ctrl_rst_dat[11][21] , \sa_ctrl_rst_dat[11][20] , 
	\sa_ctrl_rst_dat[11][19] , \sa_ctrl_rst_dat[11][18] , 
	\sa_ctrl_rst_dat[11][17] , \sa_ctrl_rst_dat[11][16] , 
	\sa_ctrl_rst_dat[11][15] , \sa_ctrl_rst_dat[11][14] , 
	\sa_ctrl_rst_dat[11][13] , \sa_ctrl_rst_dat[11][12] , 
	\sa_ctrl_rst_dat[11][11] , \sa_ctrl_rst_dat[11][10] , 
	\sa_ctrl_rst_dat[11][9] , \sa_ctrl_rst_dat[11][8] , 
	\sa_ctrl_rst_dat[11][7] , \sa_ctrl_rst_dat[11][6] , 
	\sa_ctrl_rst_dat[11][5] , \sa_ctrl_rst_dat[11][4] , 
	\sa_ctrl_rst_dat[11][3] , \sa_ctrl_rst_dat[11][2] , 
	\sa_ctrl_rst_dat[11][1] , \sa_ctrl_rst_dat[11][0] , 
	\sa_ctrl_rst_dat[10][31] , \sa_ctrl_rst_dat[10][30] , 
	\sa_ctrl_rst_dat[10][29] , \sa_ctrl_rst_dat[10][28] , 
	\sa_ctrl_rst_dat[10][27] , \sa_ctrl_rst_dat[10][26] , 
	\sa_ctrl_rst_dat[10][25] , \sa_ctrl_rst_dat[10][24] , 
	\sa_ctrl_rst_dat[10][23] , \sa_ctrl_rst_dat[10][22] , 
	\sa_ctrl_rst_dat[10][21] , \sa_ctrl_rst_dat[10][20] , 
	\sa_ctrl_rst_dat[10][19] , \sa_ctrl_rst_dat[10][18] , 
	\sa_ctrl_rst_dat[10][17] , \sa_ctrl_rst_dat[10][16] , 
	\sa_ctrl_rst_dat[10][15] , \sa_ctrl_rst_dat[10][14] , 
	\sa_ctrl_rst_dat[10][13] , \sa_ctrl_rst_dat[10][12] , 
	\sa_ctrl_rst_dat[10][11] , \sa_ctrl_rst_dat[10][10] , 
	\sa_ctrl_rst_dat[10][9] , \sa_ctrl_rst_dat[10][8] , 
	\sa_ctrl_rst_dat[10][7] , \sa_ctrl_rst_dat[10][6] , 
	\sa_ctrl_rst_dat[10][5] , \sa_ctrl_rst_dat[10][4] , 
	\sa_ctrl_rst_dat[10][3] , \sa_ctrl_rst_dat[10][2] , 
	\sa_ctrl_rst_dat[10][1] , \sa_ctrl_rst_dat[10][0] , 
	\sa_ctrl_rst_dat[9][31] , \sa_ctrl_rst_dat[9][30] , 
	\sa_ctrl_rst_dat[9][29] , \sa_ctrl_rst_dat[9][28] , 
	\sa_ctrl_rst_dat[9][27] , \sa_ctrl_rst_dat[9][26] , 
	\sa_ctrl_rst_dat[9][25] , \sa_ctrl_rst_dat[9][24] , 
	\sa_ctrl_rst_dat[9][23] , \sa_ctrl_rst_dat[9][22] , 
	\sa_ctrl_rst_dat[9][21] , \sa_ctrl_rst_dat[9][20] , 
	\sa_ctrl_rst_dat[9][19] , \sa_ctrl_rst_dat[9][18] , 
	\sa_ctrl_rst_dat[9][17] , \sa_ctrl_rst_dat[9][16] , 
	\sa_ctrl_rst_dat[9][15] , \sa_ctrl_rst_dat[9][14] , 
	\sa_ctrl_rst_dat[9][13] , \sa_ctrl_rst_dat[9][12] , 
	\sa_ctrl_rst_dat[9][11] , \sa_ctrl_rst_dat[9][10] , 
	\sa_ctrl_rst_dat[9][9] , \sa_ctrl_rst_dat[9][8] , 
	\sa_ctrl_rst_dat[9][7] , \sa_ctrl_rst_dat[9][6] , 
	\sa_ctrl_rst_dat[9][5] , \sa_ctrl_rst_dat[9][4] , 
	\sa_ctrl_rst_dat[9][3] , \sa_ctrl_rst_dat[9][2] , 
	\sa_ctrl_rst_dat[9][1] , \sa_ctrl_rst_dat[9][0] , 
	\sa_ctrl_rst_dat[8][31] , \sa_ctrl_rst_dat[8][30] , 
	\sa_ctrl_rst_dat[8][29] , \sa_ctrl_rst_dat[8][28] , 
	\sa_ctrl_rst_dat[8][27] , \sa_ctrl_rst_dat[8][26] , 
	\sa_ctrl_rst_dat[8][25] , \sa_ctrl_rst_dat[8][24] , 
	\sa_ctrl_rst_dat[8][23] , \sa_ctrl_rst_dat[8][22] , 
	\sa_ctrl_rst_dat[8][21] , \sa_ctrl_rst_dat[8][20] , 
	\sa_ctrl_rst_dat[8][19] , \sa_ctrl_rst_dat[8][18] , 
	\sa_ctrl_rst_dat[8][17] , \sa_ctrl_rst_dat[8][16] , 
	\sa_ctrl_rst_dat[8][15] , \sa_ctrl_rst_dat[8][14] , 
	\sa_ctrl_rst_dat[8][13] , \sa_ctrl_rst_dat[8][12] , 
	\sa_ctrl_rst_dat[8][11] , \sa_ctrl_rst_dat[8][10] , 
	\sa_ctrl_rst_dat[8][9] , \sa_ctrl_rst_dat[8][8] , 
	\sa_ctrl_rst_dat[8][7] , \sa_ctrl_rst_dat[8][6] , 
	\sa_ctrl_rst_dat[8][5] , \sa_ctrl_rst_dat[8][4] , 
	\sa_ctrl_rst_dat[8][3] , \sa_ctrl_rst_dat[8][2] , 
	\sa_ctrl_rst_dat[8][1] , \sa_ctrl_rst_dat[8][0] , 
	\sa_ctrl_rst_dat[7][31] , \sa_ctrl_rst_dat[7][30] , 
	\sa_ctrl_rst_dat[7][29] , \sa_ctrl_rst_dat[7][28] , 
	\sa_ctrl_rst_dat[7][27] , \sa_ctrl_rst_dat[7][26] , 
	\sa_ctrl_rst_dat[7][25] , \sa_ctrl_rst_dat[7][24] , 
	\sa_ctrl_rst_dat[7][23] , \sa_ctrl_rst_dat[7][22] , 
	\sa_ctrl_rst_dat[7][21] , \sa_ctrl_rst_dat[7][20] , 
	\sa_ctrl_rst_dat[7][19] , \sa_ctrl_rst_dat[7][18] , 
	\sa_ctrl_rst_dat[7][17] , \sa_ctrl_rst_dat[7][16] , 
	\sa_ctrl_rst_dat[7][15] , \sa_ctrl_rst_dat[7][14] , 
	\sa_ctrl_rst_dat[7][13] , \sa_ctrl_rst_dat[7][12] , 
	\sa_ctrl_rst_dat[7][11] , \sa_ctrl_rst_dat[7][10] , 
	\sa_ctrl_rst_dat[7][9] , \sa_ctrl_rst_dat[7][8] , 
	\sa_ctrl_rst_dat[7][7] , \sa_ctrl_rst_dat[7][6] , 
	\sa_ctrl_rst_dat[7][5] , \sa_ctrl_rst_dat[7][4] , 
	\sa_ctrl_rst_dat[7][3] , \sa_ctrl_rst_dat[7][2] , 
	\sa_ctrl_rst_dat[7][1] , \sa_ctrl_rst_dat[7][0] , 
	\sa_ctrl_rst_dat[6][31] , \sa_ctrl_rst_dat[6][30] , 
	\sa_ctrl_rst_dat[6][29] , \sa_ctrl_rst_dat[6][28] , 
	\sa_ctrl_rst_dat[6][27] , \sa_ctrl_rst_dat[6][26] , 
	\sa_ctrl_rst_dat[6][25] , \sa_ctrl_rst_dat[6][24] , 
	\sa_ctrl_rst_dat[6][23] , \sa_ctrl_rst_dat[6][22] , 
	\sa_ctrl_rst_dat[6][21] , \sa_ctrl_rst_dat[6][20] , 
	\sa_ctrl_rst_dat[6][19] , \sa_ctrl_rst_dat[6][18] , 
	\sa_ctrl_rst_dat[6][17] , \sa_ctrl_rst_dat[6][16] , 
	\sa_ctrl_rst_dat[6][15] , \sa_ctrl_rst_dat[6][14] , 
	\sa_ctrl_rst_dat[6][13] , \sa_ctrl_rst_dat[6][12] , 
	\sa_ctrl_rst_dat[6][11] , \sa_ctrl_rst_dat[6][10] , 
	\sa_ctrl_rst_dat[6][9] , \sa_ctrl_rst_dat[6][8] , 
	\sa_ctrl_rst_dat[6][7] , \sa_ctrl_rst_dat[6][6] , 
	\sa_ctrl_rst_dat[6][5] , \sa_ctrl_rst_dat[6][4] , 
	\sa_ctrl_rst_dat[6][3] , \sa_ctrl_rst_dat[6][2] , 
	\sa_ctrl_rst_dat[6][1] , \sa_ctrl_rst_dat[6][0] , 
	\sa_ctrl_rst_dat[5][31] , \sa_ctrl_rst_dat[5][30] , 
	\sa_ctrl_rst_dat[5][29] , \sa_ctrl_rst_dat[5][28] , 
	\sa_ctrl_rst_dat[5][27] , \sa_ctrl_rst_dat[5][26] , 
	\sa_ctrl_rst_dat[5][25] , \sa_ctrl_rst_dat[5][24] , 
	\sa_ctrl_rst_dat[5][23] , \sa_ctrl_rst_dat[5][22] , 
	\sa_ctrl_rst_dat[5][21] , \sa_ctrl_rst_dat[5][20] , 
	\sa_ctrl_rst_dat[5][19] , \sa_ctrl_rst_dat[5][18] , 
	\sa_ctrl_rst_dat[5][17] , \sa_ctrl_rst_dat[5][16] , 
	\sa_ctrl_rst_dat[5][15] , \sa_ctrl_rst_dat[5][14] , 
	\sa_ctrl_rst_dat[5][13] , \sa_ctrl_rst_dat[5][12] , 
	\sa_ctrl_rst_dat[5][11] , \sa_ctrl_rst_dat[5][10] , 
	\sa_ctrl_rst_dat[5][9] , \sa_ctrl_rst_dat[5][8] , 
	\sa_ctrl_rst_dat[5][7] , \sa_ctrl_rst_dat[5][6] , 
	\sa_ctrl_rst_dat[5][5] , \sa_ctrl_rst_dat[5][4] , 
	\sa_ctrl_rst_dat[5][3] , \sa_ctrl_rst_dat[5][2] , 
	\sa_ctrl_rst_dat[5][1] , \sa_ctrl_rst_dat[5][0] , 
	\sa_ctrl_rst_dat[4][31] , \sa_ctrl_rst_dat[4][30] , 
	\sa_ctrl_rst_dat[4][29] , \sa_ctrl_rst_dat[4][28] , 
	\sa_ctrl_rst_dat[4][27] , \sa_ctrl_rst_dat[4][26] , 
	\sa_ctrl_rst_dat[4][25] , \sa_ctrl_rst_dat[4][24] , 
	\sa_ctrl_rst_dat[4][23] , \sa_ctrl_rst_dat[4][22] , 
	\sa_ctrl_rst_dat[4][21] , \sa_ctrl_rst_dat[4][20] , 
	\sa_ctrl_rst_dat[4][19] , \sa_ctrl_rst_dat[4][18] , 
	\sa_ctrl_rst_dat[4][17] , \sa_ctrl_rst_dat[4][16] , 
	\sa_ctrl_rst_dat[4][15] , \sa_ctrl_rst_dat[4][14] , 
	\sa_ctrl_rst_dat[4][13] , \sa_ctrl_rst_dat[4][12] , 
	\sa_ctrl_rst_dat[4][11] , \sa_ctrl_rst_dat[4][10] , 
	\sa_ctrl_rst_dat[4][9] , \sa_ctrl_rst_dat[4][8] , 
	\sa_ctrl_rst_dat[4][7] , \sa_ctrl_rst_dat[4][6] , 
	\sa_ctrl_rst_dat[4][5] , \sa_ctrl_rst_dat[4][4] , 
	\sa_ctrl_rst_dat[4][3] , \sa_ctrl_rst_dat[4][2] , 
	\sa_ctrl_rst_dat[4][1] , \sa_ctrl_rst_dat[4][0] , 
	\sa_ctrl_rst_dat[3][31] , \sa_ctrl_rst_dat[3][30] , 
	\sa_ctrl_rst_dat[3][29] , \sa_ctrl_rst_dat[3][28] , 
	\sa_ctrl_rst_dat[3][27] , \sa_ctrl_rst_dat[3][26] , 
	\sa_ctrl_rst_dat[3][25] , \sa_ctrl_rst_dat[3][24] , 
	\sa_ctrl_rst_dat[3][23] , \sa_ctrl_rst_dat[3][22] , 
	\sa_ctrl_rst_dat[3][21] , \sa_ctrl_rst_dat[3][20] , 
	\sa_ctrl_rst_dat[3][19] , \sa_ctrl_rst_dat[3][18] , 
	\sa_ctrl_rst_dat[3][17] , \sa_ctrl_rst_dat[3][16] , 
	\sa_ctrl_rst_dat[3][15] , \sa_ctrl_rst_dat[3][14] , 
	\sa_ctrl_rst_dat[3][13] , \sa_ctrl_rst_dat[3][12] , 
	\sa_ctrl_rst_dat[3][11] , \sa_ctrl_rst_dat[3][10] , 
	\sa_ctrl_rst_dat[3][9] , \sa_ctrl_rst_dat[3][8] , 
	\sa_ctrl_rst_dat[3][7] , \sa_ctrl_rst_dat[3][6] , 
	\sa_ctrl_rst_dat[3][5] , \sa_ctrl_rst_dat[3][4] , 
	\sa_ctrl_rst_dat[3][3] , \sa_ctrl_rst_dat[3][2] , 
	\sa_ctrl_rst_dat[3][1] , \sa_ctrl_rst_dat[3][0] , 
	\sa_ctrl_rst_dat[2][31] , \sa_ctrl_rst_dat[2][30] , 
	\sa_ctrl_rst_dat[2][29] , \sa_ctrl_rst_dat[2][28] , 
	\sa_ctrl_rst_dat[2][27] , \sa_ctrl_rst_dat[2][26] , 
	\sa_ctrl_rst_dat[2][25] , \sa_ctrl_rst_dat[2][24] , 
	\sa_ctrl_rst_dat[2][23] , \sa_ctrl_rst_dat[2][22] , 
	\sa_ctrl_rst_dat[2][21] , \sa_ctrl_rst_dat[2][20] , 
	\sa_ctrl_rst_dat[2][19] , \sa_ctrl_rst_dat[2][18] , 
	\sa_ctrl_rst_dat[2][17] , \sa_ctrl_rst_dat[2][16] , 
	\sa_ctrl_rst_dat[2][15] , \sa_ctrl_rst_dat[2][14] , 
	\sa_ctrl_rst_dat[2][13] , \sa_ctrl_rst_dat[2][12] , 
	\sa_ctrl_rst_dat[2][11] , \sa_ctrl_rst_dat[2][10] , 
	\sa_ctrl_rst_dat[2][9] , \sa_ctrl_rst_dat[2][8] , 
	\sa_ctrl_rst_dat[2][7] , \sa_ctrl_rst_dat[2][6] , 
	\sa_ctrl_rst_dat[2][5] , \sa_ctrl_rst_dat[2][4] , 
	\sa_ctrl_rst_dat[2][3] , \sa_ctrl_rst_dat[2][2] , 
	\sa_ctrl_rst_dat[2][1] , \sa_ctrl_rst_dat[2][0] , 
	\sa_ctrl_rst_dat[1][31] , \sa_ctrl_rst_dat[1][30] , 
	\sa_ctrl_rst_dat[1][29] , \sa_ctrl_rst_dat[1][28] , 
	\sa_ctrl_rst_dat[1][27] , \sa_ctrl_rst_dat[1][26] , 
	\sa_ctrl_rst_dat[1][25] , \sa_ctrl_rst_dat[1][24] , 
	\sa_ctrl_rst_dat[1][23] , \sa_ctrl_rst_dat[1][22] , 
	\sa_ctrl_rst_dat[1][21] , \sa_ctrl_rst_dat[1][20] , 
	\sa_ctrl_rst_dat[1][19] , \sa_ctrl_rst_dat[1][18] , 
	\sa_ctrl_rst_dat[1][17] , \sa_ctrl_rst_dat[1][16] , 
	\sa_ctrl_rst_dat[1][15] , \sa_ctrl_rst_dat[1][14] , 
	\sa_ctrl_rst_dat[1][13] , \sa_ctrl_rst_dat[1][12] , 
	\sa_ctrl_rst_dat[1][11] , \sa_ctrl_rst_dat[1][10] , 
	\sa_ctrl_rst_dat[1][9] , \sa_ctrl_rst_dat[1][8] , 
	\sa_ctrl_rst_dat[1][7] , \sa_ctrl_rst_dat[1][6] , 
	\sa_ctrl_rst_dat[1][5] , \sa_ctrl_rst_dat[1][4] , 
	\sa_ctrl_rst_dat[1][3] , \sa_ctrl_rst_dat[1][2] , 
	\sa_ctrl_rst_dat[1][1] , \sa_ctrl_rst_dat[1][0] , 
	\sa_ctrl_rst_dat[0][31] , \sa_ctrl_rst_dat[0][30] , 
	\sa_ctrl_rst_dat[0][29] , \sa_ctrl_rst_dat[0][28] , 
	\sa_ctrl_rst_dat[0][27] , \sa_ctrl_rst_dat[0][26] , 
	\sa_ctrl_rst_dat[0][25] , \sa_ctrl_rst_dat[0][24] , 
	\sa_ctrl_rst_dat[0][23] , \sa_ctrl_rst_dat[0][22] , 
	\sa_ctrl_rst_dat[0][21] , \sa_ctrl_rst_dat[0][20] , 
	\sa_ctrl_rst_dat[0][19] , \sa_ctrl_rst_dat[0][18] , 
	\sa_ctrl_rst_dat[0][17] , \sa_ctrl_rst_dat[0][16] , 
	\sa_ctrl_rst_dat[0][15] , \sa_ctrl_rst_dat[0][14] , 
	\sa_ctrl_rst_dat[0][13] , \sa_ctrl_rst_dat[0][12] , 
	\sa_ctrl_rst_dat[0][11] , \sa_ctrl_rst_dat[0][10] , 
	\sa_ctrl_rst_dat[0][9] , \sa_ctrl_rst_dat[0][8] , 
	\sa_ctrl_rst_dat[0][7] , \sa_ctrl_rst_dat[0][6] , 
	\sa_ctrl_rst_dat[0][5] , \sa_ctrl_rst_dat[0][4] , 
	\sa_ctrl_rst_dat[0][3] , \sa_ctrl_rst_dat[0][2] , 
	\sa_ctrl_rst_dat[0][1] , \sa_ctrl_rst_dat[0][0] }));
nx_roreg_indirect_access_xcm129 u_SA_COUNT ( .stat_code( 
	_zy_simnet_sa_count_ia_status_783_w$[0:2]), .stat_datawords( 
	_zy_simnet_sa_count_ia_status_784_w$[0:4]), .stat_addr( 
	_zy_simnet_sa_count_ia_status_785_w$[0:4]), .capability_lst( 
	_zy_simnet_sa_count_ia_capability_786_w$[0:15]), .capability_type( 
	_zy_simnet_sa_count_ia_capability_787_w$[0:3]), .rd_dat( 
	_zy_simnet_sa_count_ia_rdata_788_w$[0:63]), .clk( clk), .rst_n( rst_n), 
	.addr( _zy_simnet_reg_addr_789_w$[0:10]), .cmnd_op( 
	_zy_simnet_sa_count_ia_config_790_w$[0:3]), .cmnd_addr( 
	_zy_simnet_sa_count_ia_config_791_w$[0:4]), .wr_stb( 
	_zy_simnet_wr_stb_792_w$), .wr_dat( 
	_zy_simnet_sa_count_ia_wdata_793_w$[0:63]), .mem_a( { 
	\sa_count[31][63] , \sa_count[31][62] , \sa_count[31][61] , 
	\sa_count[31][60] , \sa_count[31][59] , \sa_count[31][58] , 
	\sa_count[31][57] , \sa_count[31][56] , \sa_count[31][55] , 
	\sa_count[31][54] , \sa_count[31][53] , \sa_count[31][52] , 
	\sa_count[31][51] , \sa_count[31][50] , \sa_count[31][49] , 
	\sa_count[31][48] , \sa_count[31][47] , \sa_count[31][46] , 
	\sa_count[31][45] , \sa_count[31][44] , \sa_count[31][43] , 
	\sa_count[31][42] , \sa_count[31][41] , \sa_count[31][40] , 
	\sa_count[31][39] , \sa_count[31][38] , \sa_count[31][37] , 
	\sa_count[31][36] , \sa_count[31][35] , \sa_count[31][34] , 
	\sa_count[31][33] , \sa_count[31][32] , \sa_count[31][31] , 
	\sa_count[31][30] , \sa_count[31][29] , \sa_count[31][28] , 
	\sa_count[31][27] , \sa_count[31][26] , \sa_count[31][25] , 
	\sa_count[31][24] , \sa_count[31][23] , \sa_count[31][22] , 
	\sa_count[31][21] , \sa_count[31][20] , \sa_count[31][19] , 
	\sa_count[31][18] , \sa_count[31][17] , \sa_count[31][16] , 
	\sa_count[31][15] , \sa_count[31][14] , \sa_count[31][13] , 
	\sa_count[31][12] , \sa_count[31][11] , \sa_count[31][10] , 
	\sa_count[31][9] , \sa_count[31][8] , \sa_count[31][7] , 
	\sa_count[31][6] , \sa_count[31][5] , \sa_count[31][4] , 
	\sa_count[31][3] , \sa_count[31][2] , \sa_count[31][1] , 
	\sa_count[31][0] , \sa_count[30][63] , \sa_count[30][62] , 
	\sa_count[30][61] , \sa_count[30][60] , \sa_count[30][59] , 
	\sa_count[30][58] , \sa_count[30][57] , \sa_count[30][56] , 
	\sa_count[30][55] , \sa_count[30][54] , \sa_count[30][53] , 
	\sa_count[30][52] , \sa_count[30][51] , \sa_count[30][50] , 
	\sa_count[30][49] , \sa_count[30][48] , \sa_count[30][47] , 
	\sa_count[30][46] , \sa_count[30][45] , \sa_count[30][44] , 
	\sa_count[30][43] , \sa_count[30][42] , \sa_count[30][41] , 
	\sa_count[30][40] , \sa_count[30][39] , \sa_count[30][38] , 
	\sa_count[30][37] , \sa_count[30][36] , \sa_count[30][35] , 
	\sa_count[30][34] , \sa_count[30][33] , \sa_count[30][32] , 
	\sa_count[30][31] , \sa_count[30][30] , \sa_count[30][29] , 
	\sa_count[30][28] , \sa_count[30][27] , \sa_count[30][26] , 
	\sa_count[30][25] , \sa_count[30][24] , \sa_count[30][23] , 
	\sa_count[30][22] , \sa_count[30][21] , \sa_count[30][20] , 
	\sa_count[30][19] , \sa_count[30][18] , \sa_count[30][17] , 
	\sa_count[30][16] , \sa_count[30][15] , \sa_count[30][14] , 
	\sa_count[30][13] , \sa_count[30][12] , \sa_count[30][11] , 
	\sa_count[30][10] , \sa_count[30][9] , \sa_count[30][8] , 
	\sa_count[30][7] , \sa_count[30][6] , \sa_count[30][5] , 
	\sa_count[30][4] , \sa_count[30][3] , \sa_count[30][2] , 
	\sa_count[30][1] , \sa_count[30][0] , \sa_count[29][63] , 
	\sa_count[29][62] , \sa_count[29][61] , \sa_count[29][60] , 
	\sa_count[29][59] , \sa_count[29][58] , \sa_count[29][57] , 
	\sa_count[29][56] , \sa_count[29][55] , \sa_count[29][54] , 
	\sa_count[29][53] , \sa_count[29][52] , \sa_count[29][51] , 
	\sa_count[29][50] , \sa_count[29][49] , \sa_count[29][48] , 
	\sa_count[29][47] , \sa_count[29][46] , \sa_count[29][45] , 
	\sa_count[29][44] , \sa_count[29][43] , \sa_count[29][42] , 
	\sa_count[29][41] , \sa_count[29][40] , \sa_count[29][39] , 
	\sa_count[29][38] , \sa_count[29][37] , \sa_count[29][36] , 
	\sa_count[29][35] , \sa_count[29][34] , \sa_count[29][33] , 
	\sa_count[29][32] , \sa_count[29][31] , \sa_count[29][30] , 
	\sa_count[29][29] , \sa_count[29][28] , \sa_count[29][27] , 
	\sa_count[29][26] , \sa_count[29][25] , \sa_count[29][24] , 
	\sa_count[29][23] , \sa_count[29][22] , \sa_count[29][21] , 
	\sa_count[29][20] , \sa_count[29][19] , \sa_count[29][18] , 
	\sa_count[29][17] , \sa_count[29][16] , \sa_count[29][15] , 
	\sa_count[29][14] , \sa_count[29][13] , \sa_count[29][12] , 
	\sa_count[29][11] , \sa_count[29][10] , \sa_count[29][9] , 
	\sa_count[29][8] , \sa_count[29][7] , \sa_count[29][6] , 
	\sa_count[29][5] , \sa_count[29][4] , \sa_count[29][3] , 
	\sa_count[29][2] , \sa_count[29][1] , \sa_count[29][0] , 
	\sa_count[28][63] , \sa_count[28][62] , \sa_count[28][61] , 
	\sa_count[28][60] , \sa_count[28][59] , \sa_count[28][58] , 
	\sa_count[28][57] , \sa_count[28][56] , \sa_count[28][55] , 
	\sa_count[28][54] , \sa_count[28][53] , \sa_count[28][52] , 
	\sa_count[28][51] , \sa_count[28][50] , \sa_count[28][49] , 
	\sa_count[28][48] , \sa_count[28][47] , \sa_count[28][46] , 
	\sa_count[28][45] , \sa_count[28][44] , \sa_count[28][43] , 
	\sa_count[28][42] , \sa_count[28][41] , \sa_count[28][40] , 
	\sa_count[28][39] , \sa_count[28][38] , \sa_count[28][37] , 
	\sa_count[28][36] , \sa_count[28][35] , \sa_count[28][34] , 
	\sa_count[28][33] , \sa_count[28][32] , \sa_count[28][31] , 
	\sa_count[28][30] , \sa_count[28][29] , \sa_count[28][28] , 
	\sa_count[28][27] , \sa_count[28][26] , \sa_count[28][25] , 
	\sa_count[28][24] , \sa_count[28][23] , \sa_count[28][22] , 
	\sa_count[28][21] , \sa_count[28][20] , \sa_count[28][19] , 
	\sa_count[28][18] , \sa_count[28][17] , \sa_count[28][16] , 
	\sa_count[28][15] , \sa_count[28][14] , \sa_count[28][13] , 
	\sa_count[28][12] , \sa_count[28][11] , \sa_count[28][10] , 
	\sa_count[28][9] , \sa_count[28][8] , \sa_count[28][7] , 
	\sa_count[28][6] , \sa_count[28][5] , \sa_count[28][4] , 
	\sa_count[28][3] , \sa_count[28][2] , \sa_count[28][1] , 
	\sa_count[28][0] , \sa_count[27][63] , \sa_count[27][62] , 
	\sa_count[27][61] , \sa_count[27][60] , \sa_count[27][59] , 
	\sa_count[27][58] , \sa_count[27][57] , \sa_count[27][56] , 
	\sa_count[27][55] , \sa_count[27][54] , \sa_count[27][53] , 
	\sa_count[27][52] , \sa_count[27][51] , \sa_count[27][50] , 
	\sa_count[27][49] , \sa_count[27][48] , \sa_count[27][47] , 
	\sa_count[27][46] , \sa_count[27][45] , \sa_count[27][44] , 
	\sa_count[27][43] , \sa_count[27][42] , \sa_count[27][41] , 
	\sa_count[27][40] , \sa_count[27][39] , \sa_count[27][38] , 
	\sa_count[27][37] , \sa_count[27][36] , \sa_count[27][35] , 
	\sa_count[27][34] , \sa_count[27][33] , \sa_count[27][32] , 
	\sa_count[27][31] , \sa_count[27][30] , \sa_count[27][29] , 
	\sa_count[27][28] , \sa_count[27][27] , \sa_count[27][26] , 
	\sa_count[27][25] , \sa_count[27][24] , \sa_count[27][23] , 
	\sa_count[27][22] , \sa_count[27][21] , \sa_count[27][20] , 
	\sa_count[27][19] , \sa_count[27][18] , \sa_count[27][17] , 
	\sa_count[27][16] , \sa_count[27][15] , \sa_count[27][14] , 
	\sa_count[27][13] , \sa_count[27][12] , \sa_count[27][11] , 
	\sa_count[27][10] , \sa_count[27][9] , \sa_count[27][8] , 
	\sa_count[27][7] , \sa_count[27][6] , \sa_count[27][5] , 
	\sa_count[27][4] , \sa_count[27][3] , \sa_count[27][2] , 
	\sa_count[27][1] , \sa_count[27][0] , \sa_count[26][63] , 
	\sa_count[26][62] , \sa_count[26][61] , \sa_count[26][60] , 
	\sa_count[26][59] , \sa_count[26][58] , \sa_count[26][57] , 
	\sa_count[26][56] , \sa_count[26][55] , \sa_count[26][54] , 
	\sa_count[26][53] , \sa_count[26][52] , \sa_count[26][51] , 
	\sa_count[26][50] , \sa_count[26][49] , \sa_count[26][48] , 
	\sa_count[26][47] , \sa_count[26][46] , \sa_count[26][45] , 
	\sa_count[26][44] , \sa_count[26][43] , \sa_count[26][42] , 
	\sa_count[26][41] , \sa_count[26][40] , \sa_count[26][39] , 
	\sa_count[26][38] , \sa_count[26][37] , \sa_count[26][36] , 
	\sa_count[26][35] , \sa_count[26][34] , \sa_count[26][33] , 
	\sa_count[26][32] , \sa_count[26][31] , \sa_count[26][30] , 
	\sa_count[26][29] , \sa_count[26][28] , \sa_count[26][27] , 
	\sa_count[26][26] , \sa_count[26][25] , \sa_count[26][24] , 
	\sa_count[26][23] , \sa_count[26][22] , \sa_count[26][21] , 
	\sa_count[26][20] , \sa_count[26][19] , \sa_count[26][18] , 
	\sa_count[26][17] , \sa_count[26][16] , \sa_count[26][15] , 
	\sa_count[26][14] , \sa_count[26][13] , \sa_count[26][12] , 
	\sa_count[26][11] , \sa_count[26][10] , \sa_count[26][9] , 
	\sa_count[26][8] , \sa_count[26][7] , \sa_count[26][6] , 
	\sa_count[26][5] , \sa_count[26][4] , \sa_count[26][3] , 
	\sa_count[26][2] , \sa_count[26][1] , \sa_count[26][0] , 
	\sa_count[25][63] , \sa_count[25][62] , \sa_count[25][61] , 
	\sa_count[25][60] , \sa_count[25][59] , \sa_count[25][58] , 
	\sa_count[25][57] , \sa_count[25][56] , \sa_count[25][55] , 
	\sa_count[25][54] , \sa_count[25][53] , \sa_count[25][52] , 
	\sa_count[25][51] , \sa_count[25][50] , \sa_count[25][49] , 
	\sa_count[25][48] , \sa_count[25][47] , \sa_count[25][46] , 
	\sa_count[25][45] , \sa_count[25][44] , \sa_count[25][43] , 
	\sa_count[25][42] , \sa_count[25][41] , \sa_count[25][40] , 
	\sa_count[25][39] , \sa_count[25][38] , \sa_count[25][37] , 
	\sa_count[25][36] , \sa_count[25][35] , \sa_count[25][34] , 
	\sa_count[25][33] , \sa_count[25][32] , \sa_count[25][31] , 
	\sa_count[25][30] , \sa_count[25][29] , \sa_count[25][28] , 
	\sa_count[25][27] , \sa_count[25][26] , \sa_count[25][25] , 
	\sa_count[25][24] , \sa_count[25][23] , \sa_count[25][22] , 
	\sa_count[25][21] , \sa_count[25][20] , \sa_count[25][19] , 
	\sa_count[25][18] , \sa_count[25][17] , \sa_count[25][16] , 
	\sa_count[25][15] , \sa_count[25][14] , \sa_count[25][13] , 
	\sa_count[25][12] , \sa_count[25][11] , \sa_count[25][10] , 
	\sa_count[25][9] , \sa_count[25][8] , \sa_count[25][7] , 
	\sa_count[25][6] , \sa_count[25][5] , \sa_count[25][4] , 
	\sa_count[25][3] , \sa_count[25][2] , \sa_count[25][1] , 
	\sa_count[25][0] , \sa_count[24][63] , \sa_count[24][62] , 
	\sa_count[24][61] , \sa_count[24][60] , \sa_count[24][59] , 
	\sa_count[24][58] , \sa_count[24][57] , \sa_count[24][56] , 
	\sa_count[24][55] , \sa_count[24][54] , \sa_count[24][53] , 
	\sa_count[24][52] , \sa_count[24][51] , \sa_count[24][50] , 
	\sa_count[24][49] , \sa_count[24][48] , \sa_count[24][47] , 
	\sa_count[24][46] , \sa_count[24][45] , \sa_count[24][44] , 
	\sa_count[24][43] , \sa_count[24][42] , \sa_count[24][41] , 
	\sa_count[24][40] , \sa_count[24][39] , \sa_count[24][38] , 
	\sa_count[24][37] , \sa_count[24][36] , \sa_count[24][35] , 
	\sa_count[24][34] , \sa_count[24][33] , \sa_count[24][32] , 
	\sa_count[24][31] , \sa_count[24][30] , \sa_count[24][29] , 
	\sa_count[24][28] , \sa_count[24][27] , \sa_count[24][26] , 
	\sa_count[24][25] , \sa_count[24][24] , \sa_count[24][23] , 
	\sa_count[24][22] , \sa_count[24][21] , \sa_count[24][20] , 
	\sa_count[24][19] , \sa_count[24][18] , \sa_count[24][17] , 
	\sa_count[24][16] , \sa_count[24][15] , \sa_count[24][14] , 
	\sa_count[24][13] , \sa_count[24][12] , \sa_count[24][11] , 
	\sa_count[24][10] , \sa_count[24][9] , \sa_count[24][8] , 
	\sa_count[24][7] , \sa_count[24][6] , \sa_count[24][5] , 
	\sa_count[24][4] , \sa_count[24][3] , \sa_count[24][2] , 
	\sa_count[24][1] , \sa_count[24][0] , \sa_count[23][63] , 
	\sa_count[23][62] , \sa_count[23][61] , \sa_count[23][60] , 
	\sa_count[23][59] , \sa_count[23][58] , \sa_count[23][57] , 
	\sa_count[23][56] , \sa_count[23][55] , \sa_count[23][54] , 
	\sa_count[23][53] , \sa_count[23][52] , \sa_count[23][51] , 
	\sa_count[23][50] , \sa_count[23][49] , \sa_count[23][48] , 
	\sa_count[23][47] , \sa_count[23][46] , \sa_count[23][45] , 
	\sa_count[23][44] , \sa_count[23][43] , \sa_count[23][42] , 
	\sa_count[23][41] , \sa_count[23][40] , \sa_count[23][39] , 
	\sa_count[23][38] , \sa_count[23][37] , \sa_count[23][36] , 
	\sa_count[23][35] , \sa_count[23][34] , \sa_count[23][33] , 
	\sa_count[23][32] , \sa_count[23][31] , \sa_count[23][30] , 
	\sa_count[23][29] , \sa_count[23][28] , \sa_count[23][27] , 
	\sa_count[23][26] , \sa_count[23][25] , \sa_count[23][24] , 
	\sa_count[23][23] , \sa_count[23][22] , \sa_count[23][21] , 
	\sa_count[23][20] , \sa_count[23][19] , \sa_count[23][18] , 
	\sa_count[23][17] , \sa_count[23][16] , \sa_count[23][15] , 
	\sa_count[23][14] , \sa_count[23][13] , \sa_count[23][12] , 
	\sa_count[23][11] , \sa_count[23][10] , \sa_count[23][9] , 
	\sa_count[23][8] , \sa_count[23][7] , \sa_count[23][6] , 
	\sa_count[23][5] , \sa_count[23][4] , \sa_count[23][3] , 
	\sa_count[23][2] , \sa_count[23][1] , \sa_count[23][0] , 
	\sa_count[22][63] , \sa_count[22][62] , \sa_count[22][61] , 
	\sa_count[22][60] , \sa_count[22][59] , \sa_count[22][58] , 
	\sa_count[22][57] , \sa_count[22][56] , \sa_count[22][55] , 
	\sa_count[22][54] , \sa_count[22][53] , \sa_count[22][52] , 
	\sa_count[22][51] , \sa_count[22][50] , \sa_count[22][49] , 
	\sa_count[22][48] , \sa_count[22][47] , \sa_count[22][46] , 
	\sa_count[22][45] , \sa_count[22][44] , \sa_count[22][43] , 
	\sa_count[22][42] , \sa_count[22][41] , \sa_count[22][40] , 
	\sa_count[22][39] , \sa_count[22][38] , \sa_count[22][37] , 
	\sa_count[22][36] , \sa_count[22][35] , \sa_count[22][34] , 
	\sa_count[22][33] , \sa_count[22][32] , \sa_count[22][31] , 
	\sa_count[22][30] , \sa_count[22][29] , \sa_count[22][28] , 
	\sa_count[22][27] , \sa_count[22][26] , \sa_count[22][25] , 
	\sa_count[22][24] , \sa_count[22][23] , \sa_count[22][22] , 
	\sa_count[22][21] , \sa_count[22][20] , \sa_count[22][19] , 
	\sa_count[22][18] , \sa_count[22][17] , \sa_count[22][16] , 
	\sa_count[22][15] , \sa_count[22][14] , \sa_count[22][13] , 
	\sa_count[22][12] , \sa_count[22][11] , \sa_count[22][10] , 
	\sa_count[22][9] , \sa_count[22][8] , \sa_count[22][7] , 
	\sa_count[22][6] , \sa_count[22][5] , \sa_count[22][4] , 
	\sa_count[22][3] , \sa_count[22][2] , \sa_count[22][1] , 
	\sa_count[22][0] , \sa_count[21][63] , \sa_count[21][62] , 
	\sa_count[21][61] , \sa_count[21][60] , \sa_count[21][59] , 
	\sa_count[21][58] , \sa_count[21][57] , \sa_count[21][56] , 
	\sa_count[21][55] , \sa_count[21][54] , \sa_count[21][53] , 
	\sa_count[21][52] , \sa_count[21][51] , \sa_count[21][50] , 
	\sa_count[21][49] , \sa_count[21][48] , \sa_count[21][47] , 
	\sa_count[21][46] , \sa_count[21][45] , \sa_count[21][44] , 
	\sa_count[21][43] , \sa_count[21][42] , \sa_count[21][41] , 
	\sa_count[21][40] , \sa_count[21][39] , \sa_count[21][38] , 
	\sa_count[21][37] , \sa_count[21][36] , \sa_count[21][35] , 
	\sa_count[21][34] , \sa_count[21][33] , \sa_count[21][32] , 
	\sa_count[21][31] , \sa_count[21][30] , \sa_count[21][29] , 
	\sa_count[21][28] , \sa_count[21][27] , \sa_count[21][26] , 
	\sa_count[21][25] , \sa_count[21][24] , \sa_count[21][23] , 
	\sa_count[21][22] , \sa_count[21][21] , \sa_count[21][20] , 
	\sa_count[21][19] , \sa_count[21][18] , \sa_count[21][17] , 
	\sa_count[21][16] , \sa_count[21][15] , \sa_count[21][14] , 
	\sa_count[21][13] , \sa_count[21][12] , \sa_count[21][11] , 
	\sa_count[21][10] , \sa_count[21][9] , \sa_count[21][8] , 
	\sa_count[21][7] , \sa_count[21][6] , \sa_count[21][5] , 
	\sa_count[21][4] , \sa_count[21][3] , \sa_count[21][2] , 
	\sa_count[21][1] , \sa_count[21][0] , \sa_count[20][63] , 
	\sa_count[20][62] , \sa_count[20][61] , \sa_count[20][60] , 
	\sa_count[20][59] , \sa_count[20][58] , \sa_count[20][57] , 
	\sa_count[20][56] , \sa_count[20][55] , \sa_count[20][54] , 
	\sa_count[20][53] , \sa_count[20][52] , \sa_count[20][51] , 
	\sa_count[20][50] , \sa_count[20][49] , \sa_count[20][48] , 
	\sa_count[20][47] , \sa_count[20][46] , \sa_count[20][45] , 
	\sa_count[20][44] , \sa_count[20][43] , \sa_count[20][42] , 
	\sa_count[20][41] , \sa_count[20][40] , \sa_count[20][39] , 
	\sa_count[20][38] , \sa_count[20][37] , \sa_count[20][36] , 
	\sa_count[20][35] , \sa_count[20][34] , \sa_count[20][33] , 
	\sa_count[20][32] , \sa_count[20][31] , \sa_count[20][30] , 
	\sa_count[20][29] , \sa_count[20][28] , \sa_count[20][27] , 
	\sa_count[20][26] , \sa_count[20][25] , \sa_count[20][24] , 
	\sa_count[20][23] , \sa_count[20][22] , \sa_count[20][21] , 
	\sa_count[20][20] , \sa_count[20][19] , \sa_count[20][18] , 
	\sa_count[20][17] , \sa_count[20][16] , \sa_count[20][15] , 
	\sa_count[20][14] , \sa_count[20][13] , \sa_count[20][12] , 
	\sa_count[20][11] , \sa_count[20][10] , \sa_count[20][9] , 
	\sa_count[20][8] , \sa_count[20][7] , \sa_count[20][6] , 
	\sa_count[20][5] , \sa_count[20][4] , \sa_count[20][3] , 
	\sa_count[20][2] , \sa_count[20][1] , \sa_count[20][0] , 
	\sa_count[19][63] , \sa_count[19][62] , \sa_count[19][61] , 
	\sa_count[19][60] , \sa_count[19][59] , \sa_count[19][58] , 
	\sa_count[19][57] , \sa_count[19][56] , \sa_count[19][55] , 
	\sa_count[19][54] , \sa_count[19][53] , \sa_count[19][52] , 
	\sa_count[19][51] , \sa_count[19][50] , \sa_count[19][49] , 
	\sa_count[19][48] , \sa_count[19][47] , \sa_count[19][46] , 
	\sa_count[19][45] , \sa_count[19][44] , \sa_count[19][43] , 
	\sa_count[19][42] , \sa_count[19][41] , \sa_count[19][40] , 
	\sa_count[19][39] , \sa_count[19][38] , \sa_count[19][37] , 
	\sa_count[19][36] , \sa_count[19][35] , \sa_count[19][34] , 
	\sa_count[19][33] , \sa_count[19][32] , \sa_count[19][31] , 
	\sa_count[19][30] , \sa_count[19][29] , \sa_count[19][28] , 
	\sa_count[19][27] , \sa_count[19][26] , \sa_count[19][25] , 
	\sa_count[19][24] , \sa_count[19][23] , \sa_count[19][22] , 
	\sa_count[19][21] , \sa_count[19][20] , \sa_count[19][19] , 
	\sa_count[19][18] , \sa_count[19][17] , \sa_count[19][16] , 
	\sa_count[19][15] , \sa_count[19][14] , \sa_count[19][13] , 
	\sa_count[19][12] , \sa_count[19][11] , \sa_count[19][10] , 
	\sa_count[19][9] , \sa_count[19][8] , \sa_count[19][7] , 
	\sa_count[19][6] , \sa_count[19][5] , \sa_count[19][4] , 
	\sa_count[19][3] , \sa_count[19][2] , \sa_count[19][1] , 
	\sa_count[19][0] , \sa_count[18][63] , \sa_count[18][62] , 
	\sa_count[18][61] , \sa_count[18][60] , \sa_count[18][59] , 
	\sa_count[18][58] , \sa_count[18][57] , \sa_count[18][56] , 
	\sa_count[18][55] , \sa_count[18][54] , \sa_count[18][53] , 
	\sa_count[18][52] , \sa_count[18][51] , \sa_count[18][50] , 
	\sa_count[18][49] , \sa_count[18][48] , \sa_count[18][47] , 
	\sa_count[18][46] , \sa_count[18][45] , \sa_count[18][44] , 
	\sa_count[18][43] , \sa_count[18][42] , \sa_count[18][41] , 
	\sa_count[18][40] , \sa_count[18][39] , \sa_count[18][38] , 
	\sa_count[18][37] , \sa_count[18][36] , \sa_count[18][35] , 
	\sa_count[18][34] , \sa_count[18][33] , \sa_count[18][32] , 
	\sa_count[18][31] , \sa_count[18][30] , \sa_count[18][29] , 
	\sa_count[18][28] , \sa_count[18][27] , \sa_count[18][26] , 
	\sa_count[18][25] , \sa_count[18][24] , \sa_count[18][23] , 
	\sa_count[18][22] , \sa_count[18][21] , \sa_count[18][20] , 
	\sa_count[18][19] , \sa_count[18][18] , \sa_count[18][17] , 
	\sa_count[18][16] , \sa_count[18][15] , \sa_count[18][14] , 
	\sa_count[18][13] , \sa_count[18][12] , \sa_count[18][11] , 
	\sa_count[18][10] , \sa_count[18][9] , \sa_count[18][8] , 
	\sa_count[18][7] , \sa_count[18][6] , \sa_count[18][5] , 
	\sa_count[18][4] , \sa_count[18][3] , \sa_count[18][2] , 
	\sa_count[18][1] , \sa_count[18][0] , \sa_count[17][63] , 
	\sa_count[17][62] , \sa_count[17][61] , \sa_count[17][60] , 
	\sa_count[17][59] , \sa_count[17][58] , \sa_count[17][57] , 
	\sa_count[17][56] , \sa_count[17][55] , \sa_count[17][54] , 
	\sa_count[17][53] , \sa_count[17][52] , \sa_count[17][51] , 
	\sa_count[17][50] , \sa_count[17][49] , \sa_count[17][48] , 
	\sa_count[17][47] , \sa_count[17][46] , \sa_count[17][45] , 
	\sa_count[17][44] , \sa_count[17][43] , \sa_count[17][42] , 
	\sa_count[17][41] , \sa_count[17][40] , \sa_count[17][39] , 
	\sa_count[17][38] , \sa_count[17][37] , \sa_count[17][36] , 
	\sa_count[17][35] , \sa_count[17][34] , \sa_count[17][33] , 
	\sa_count[17][32] , \sa_count[17][31] , \sa_count[17][30] , 
	\sa_count[17][29] , \sa_count[17][28] , \sa_count[17][27] , 
	\sa_count[17][26] , \sa_count[17][25] , \sa_count[17][24] , 
	\sa_count[17][23] , \sa_count[17][22] , \sa_count[17][21] , 
	\sa_count[17][20] , \sa_count[17][19] , \sa_count[17][18] , 
	\sa_count[17][17] , \sa_count[17][16] , \sa_count[17][15] , 
	\sa_count[17][14] , \sa_count[17][13] , \sa_count[17][12] , 
	\sa_count[17][11] , \sa_count[17][10] , \sa_count[17][9] , 
	\sa_count[17][8] , \sa_count[17][7] , \sa_count[17][6] , 
	\sa_count[17][5] , \sa_count[17][4] , \sa_count[17][3] , 
	\sa_count[17][2] , \sa_count[17][1] , \sa_count[17][0] , 
	\sa_count[16][63] , \sa_count[16][62] , \sa_count[16][61] , 
	\sa_count[16][60] , \sa_count[16][59] , \sa_count[16][58] , 
	\sa_count[16][57] , \sa_count[16][56] , \sa_count[16][55] , 
	\sa_count[16][54] , \sa_count[16][53] , \sa_count[16][52] , 
	\sa_count[16][51] , \sa_count[16][50] , \sa_count[16][49] , 
	\sa_count[16][48] , \sa_count[16][47] , \sa_count[16][46] , 
	\sa_count[16][45] , \sa_count[16][44] , \sa_count[16][43] , 
	\sa_count[16][42] , \sa_count[16][41] , \sa_count[16][40] , 
	\sa_count[16][39] , \sa_count[16][38] , \sa_count[16][37] , 
	\sa_count[16][36] , \sa_count[16][35] , \sa_count[16][34] , 
	\sa_count[16][33] , \sa_count[16][32] , \sa_count[16][31] , 
	\sa_count[16][30] , \sa_count[16][29] , \sa_count[16][28] , 
	\sa_count[16][27] , \sa_count[16][26] , \sa_count[16][25] , 
	\sa_count[16][24] , \sa_count[16][23] , \sa_count[16][22] , 
	\sa_count[16][21] , \sa_count[16][20] , \sa_count[16][19] , 
	\sa_count[16][18] , \sa_count[16][17] , \sa_count[16][16] , 
	\sa_count[16][15] , \sa_count[16][14] , \sa_count[16][13] , 
	\sa_count[16][12] , \sa_count[16][11] , \sa_count[16][10] , 
	\sa_count[16][9] , \sa_count[16][8] , \sa_count[16][7] , 
	\sa_count[16][6] , \sa_count[16][5] , \sa_count[16][4] , 
	\sa_count[16][3] , \sa_count[16][2] , \sa_count[16][1] , 
	\sa_count[16][0] , \sa_count[15][63] , \sa_count[15][62] , 
	\sa_count[15][61] , \sa_count[15][60] , \sa_count[15][59] , 
	\sa_count[15][58] , \sa_count[15][57] , \sa_count[15][56] , 
	\sa_count[15][55] , \sa_count[15][54] , \sa_count[15][53] , 
	\sa_count[15][52] , \sa_count[15][51] , \sa_count[15][50] , 
	\sa_count[15][49] , \sa_count[15][48] , \sa_count[15][47] , 
	\sa_count[15][46] , \sa_count[15][45] , \sa_count[15][44] , 
	\sa_count[15][43] , \sa_count[15][42] , \sa_count[15][41] , 
	\sa_count[15][40] , \sa_count[15][39] , \sa_count[15][38] , 
	\sa_count[15][37] , \sa_count[15][36] , \sa_count[15][35] , 
	\sa_count[15][34] , \sa_count[15][33] , \sa_count[15][32] , 
	\sa_count[15][31] , \sa_count[15][30] , \sa_count[15][29] , 
	\sa_count[15][28] , \sa_count[15][27] , \sa_count[15][26] , 
	\sa_count[15][25] , \sa_count[15][24] , \sa_count[15][23] , 
	\sa_count[15][22] , \sa_count[15][21] , \sa_count[15][20] , 
	\sa_count[15][19] , \sa_count[15][18] , \sa_count[15][17] , 
	\sa_count[15][16] , \sa_count[15][15] , \sa_count[15][14] , 
	\sa_count[15][13] , \sa_count[15][12] , \sa_count[15][11] , 
	\sa_count[15][10] , \sa_count[15][9] , \sa_count[15][8] , 
	\sa_count[15][7] , \sa_count[15][6] , \sa_count[15][5] , 
	\sa_count[15][4] , \sa_count[15][3] , \sa_count[15][2] , 
	\sa_count[15][1] , \sa_count[15][0] , \sa_count[14][63] , 
	\sa_count[14][62] , \sa_count[14][61] , \sa_count[14][60] , 
	\sa_count[14][59] , \sa_count[14][58] , \sa_count[14][57] , 
	\sa_count[14][56] , \sa_count[14][55] , \sa_count[14][54] , 
	\sa_count[14][53] , \sa_count[14][52] , \sa_count[14][51] , 
	\sa_count[14][50] , \sa_count[14][49] , \sa_count[14][48] , 
	\sa_count[14][47] , \sa_count[14][46] , \sa_count[14][45] , 
	\sa_count[14][44] , \sa_count[14][43] , \sa_count[14][42] , 
	\sa_count[14][41] , \sa_count[14][40] , \sa_count[14][39] , 
	\sa_count[14][38] , \sa_count[14][37] , \sa_count[14][36] , 
	\sa_count[14][35] , \sa_count[14][34] , \sa_count[14][33] , 
	\sa_count[14][32] , \sa_count[14][31] , \sa_count[14][30] , 
	\sa_count[14][29] , \sa_count[14][28] , \sa_count[14][27] , 
	\sa_count[14][26] , \sa_count[14][25] , \sa_count[14][24] , 
	\sa_count[14][23] , \sa_count[14][22] , \sa_count[14][21] , 
	\sa_count[14][20] , \sa_count[14][19] , \sa_count[14][18] , 
	\sa_count[14][17] , \sa_count[14][16] , \sa_count[14][15] , 
	\sa_count[14][14] , \sa_count[14][13] , \sa_count[14][12] , 
	\sa_count[14][11] , \sa_count[14][10] , \sa_count[14][9] , 
	\sa_count[14][8] , \sa_count[14][7] , \sa_count[14][6] , 
	\sa_count[14][5] , \sa_count[14][4] , \sa_count[14][3] , 
	\sa_count[14][2] , \sa_count[14][1] , \sa_count[14][0] , 
	\sa_count[13][63] , \sa_count[13][62] , \sa_count[13][61] , 
	\sa_count[13][60] , \sa_count[13][59] , \sa_count[13][58] , 
	\sa_count[13][57] , \sa_count[13][56] , \sa_count[13][55] , 
	\sa_count[13][54] , \sa_count[13][53] , \sa_count[13][52] , 
	\sa_count[13][51] , \sa_count[13][50] , \sa_count[13][49] , 
	\sa_count[13][48] , \sa_count[13][47] , \sa_count[13][46] , 
	\sa_count[13][45] , \sa_count[13][44] , \sa_count[13][43] , 
	\sa_count[13][42] , \sa_count[13][41] , \sa_count[13][40] , 
	\sa_count[13][39] , \sa_count[13][38] , \sa_count[13][37] , 
	\sa_count[13][36] , \sa_count[13][35] , \sa_count[13][34] , 
	\sa_count[13][33] , \sa_count[13][32] , \sa_count[13][31] , 
	\sa_count[13][30] , \sa_count[13][29] , \sa_count[13][28] , 
	\sa_count[13][27] , \sa_count[13][26] , \sa_count[13][25] , 
	\sa_count[13][24] , \sa_count[13][23] , \sa_count[13][22] , 
	\sa_count[13][21] , \sa_count[13][20] , \sa_count[13][19] , 
	\sa_count[13][18] , \sa_count[13][17] , \sa_count[13][16] , 
	\sa_count[13][15] , \sa_count[13][14] , \sa_count[13][13] , 
	\sa_count[13][12] , \sa_count[13][11] , \sa_count[13][10] , 
	\sa_count[13][9] , \sa_count[13][8] , \sa_count[13][7] , 
	\sa_count[13][6] , \sa_count[13][5] , \sa_count[13][4] , 
	\sa_count[13][3] , \sa_count[13][2] , \sa_count[13][1] , 
	\sa_count[13][0] , \sa_count[12][63] , \sa_count[12][62] , 
	\sa_count[12][61] , \sa_count[12][60] , \sa_count[12][59] , 
	\sa_count[12][58] , \sa_count[12][57] , \sa_count[12][56] , 
	\sa_count[12][55] , \sa_count[12][54] , \sa_count[12][53] , 
	\sa_count[12][52] , \sa_count[12][51] , \sa_count[12][50] , 
	\sa_count[12][49] , \sa_count[12][48] , \sa_count[12][47] , 
	\sa_count[12][46] , \sa_count[12][45] , \sa_count[12][44] , 
	\sa_count[12][43] , \sa_count[12][42] , \sa_count[12][41] , 
	\sa_count[12][40] , \sa_count[12][39] , \sa_count[12][38] , 
	\sa_count[12][37] , \sa_count[12][36] , \sa_count[12][35] , 
	\sa_count[12][34] , \sa_count[12][33] , \sa_count[12][32] , 
	\sa_count[12][31] , \sa_count[12][30] , \sa_count[12][29] , 
	\sa_count[12][28] , \sa_count[12][27] , \sa_count[12][26] , 
	\sa_count[12][25] , \sa_count[12][24] , \sa_count[12][23] , 
	\sa_count[12][22] , \sa_count[12][21] , \sa_count[12][20] , 
	\sa_count[12][19] , \sa_count[12][18] , \sa_count[12][17] , 
	\sa_count[12][16] , \sa_count[12][15] , \sa_count[12][14] , 
	\sa_count[12][13] , \sa_count[12][12] , \sa_count[12][11] , 
	\sa_count[12][10] , \sa_count[12][9] , \sa_count[12][8] , 
	\sa_count[12][7] , \sa_count[12][6] , \sa_count[12][5] , 
	\sa_count[12][4] , \sa_count[12][3] , \sa_count[12][2] , 
	\sa_count[12][1] , \sa_count[12][0] , \sa_count[11][63] , 
	\sa_count[11][62] , \sa_count[11][61] , \sa_count[11][60] , 
	\sa_count[11][59] , \sa_count[11][58] , \sa_count[11][57] , 
	\sa_count[11][56] , \sa_count[11][55] , \sa_count[11][54] , 
	\sa_count[11][53] , \sa_count[11][52] , \sa_count[11][51] , 
	\sa_count[11][50] , \sa_count[11][49] , \sa_count[11][48] , 
	\sa_count[11][47] , \sa_count[11][46] , \sa_count[11][45] , 
	\sa_count[11][44] , \sa_count[11][43] , \sa_count[11][42] , 
	\sa_count[11][41] , \sa_count[11][40] , \sa_count[11][39] , 
	\sa_count[11][38] , \sa_count[11][37] , \sa_count[11][36] , 
	\sa_count[11][35] , \sa_count[11][34] , \sa_count[11][33] , 
	\sa_count[11][32] , \sa_count[11][31] , \sa_count[11][30] , 
	\sa_count[11][29] , \sa_count[11][28] , \sa_count[11][27] , 
	\sa_count[11][26] , \sa_count[11][25] , \sa_count[11][24] , 
	\sa_count[11][23] , \sa_count[11][22] , \sa_count[11][21] , 
	\sa_count[11][20] , \sa_count[11][19] , \sa_count[11][18] , 
	\sa_count[11][17] , \sa_count[11][16] , \sa_count[11][15] , 
	\sa_count[11][14] , \sa_count[11][13] , \sa_count[11][12] , 
	\sa_count[11][11] , \sa_count[11][10] , \sa_count[11][9] , 
	\sa_count[11][8] , \sa_count[11][7] , \sa_count[11][6] , 
	\sa_count[11][5] , \sa_count[11][4] , \sa_count[11][3] , 
	\sa_count[11][2] , \sa_count[11][1] , \sa_count[11][0] , 
	\sa_count[10][63] , \sa_count[10][62] , \sa_count[10][61] , 
	\sa_count[10][60] , \sa_count[10][59] , \sa_count[10][58] , 
	\sa_count[10][57] , \sa_count[10][56] , \sa_count[10][55] , 
	\sa_count[10][54] , \sa_count[10][53] , \sa_count[10][52] , 
	\sa_count[10][51] , \sa_count[10][50] , \sa_count[10][49] , 
	\sa_count[10][48] , \sa_count[10][47] , \sa_count[10][46] , 
	\sa_count[10][45] , \sa_count[10][44] , \sa_count[10][43] , 
	\sa_count[10][42] , \sa_count[10][41] , \sa_count[10][40] , 
	\sa_count[10][39] , \sa_count[10][38] , \sa_count[10][37] , 
	\sa_count[10][36] , \sa_count[10][35] , \sa_count[10][34] , 
	\sa_count[10][33] , \sa_count[10][32] , \sa_count[10][31] , 
	\sa_count[10][30] , \sa_count[10][29] , \sa_count[10][28] , 
	\sa_count[10][27] , \sa_count[10][26] , \sa_count[10][25] , 
	\sa_count[10][24] , \sa_count[10][23] , \sa_count[10][22] , 
	\sa_count[10][21] , \sa_count[10][20] , \sa_count[10][19] , 
	\sa_count[10][18] , \sa_count[10][17] , \sa_count[10][16] , 
	\sa_count[10][15] , \sa_count[10][14] , \sa_count[10][13] , 
	\sa_count[10][12] , \sa_count[10][11] , \sa_count[10][10] , 
	\sa_count[10][9] , \sa_count[10][8] , \sa_count[10][7] , 
	\sa_count[10][6] , \sa_count[10][5] , \sa_count[10][4] , 
	\sa_count[10][3] , \sa_count[10][2] , \sa_count[10][1] , 
	\sa_count[10][0] , \sa_count[9][63] , \sa_count[9][62] , 
	\sa_count[9][61] , \sa_count[9][60] , \sa_count[9][59] , 
	\sa_count[9][58] , \sa_count[9][57] , \sa_count[9][56] , 
	\sa_count[9][55] , \sa_count[9][54] , \sa_count[9][53] , 
	\sa_count[9][52] , \sa_count[9][51] , \sa_count[9][50] , 
	\sa_count[9][49] , \sa_count[9][48] , \sa_count[9][47] , 
	\sa_count[9][46] , \sa_count[9][45] , \sa_count[9][44] , 
	\sa_count[9][43] , \sa_count[9][42] , \sa_count[9][41] , 
	\sa_count[9][40] , \sa_count[9][39] , \sa_count[9][38] , 
	\sa_count[9][37] , \sa_count[9][36] , \sa_count[9][35] , 
	\sa_count[9][34] , \sa_count[9][33] , \sa_count[9][32] , 
	\sa_count[9][31] , \sa_count[9][30] , \sa_count[9][29] , 
	\sa_count[9][28] , \sa_count[9][27] , \sa_count[9][26] , 
	\sa_count[9][25] , \sa_count[9][24] , \sa_count[9][23] , 
	\sa_count[9][22] , \sa_count[9][21] , \sa_count[9][20] , 
	\sa_count[9][19] , \sa_count[9][18] , \sa_count[9][17] , 
	\sa_count[9][16] , \sa_count[9][15] , \sa_count[9][14] , 
	\sa_count[9][13] , \sa_count[9][12] , \sa_count[9][11] , 
	\sa_count[9][10] , \sa_count[9][9] , \sa_count[9][8] , 
	\sa_count[9][7] , \sa_count[9][6] , \sa_count[9][5] , 
	\sa_count[9][4] , \sa_count[9][3] , \sa_count[9][2] , 
	\sa_count[9][1] , \sa_count[9][0] , \sa_count[8][63] , 
	\sa_count[8][62] , \sa_count[8][61] , \sa_count[8][60] , 
	\sa_count[8][59] , \sa_count[8][58] , \sa_count[8][57] , 
	\sa_count[8][56] , \sa_count[8][55] , \sa_count[8][54] , 
	\sa_count[8][53] , \sa_count[8][52] , \sa_count[8][51] , 
	\sa_count[8][50] , \sa_count[8][49] , \sa_count[8][48] , 
	\sa_count[8][47] , \sa_count[8][46] , \sa_count[8][45] , 
	\sa_count[8][44] , \sa_count[8][43] , \sa_count[8][42] , 
	\sa_count[8][41] , \sa_count[8][40] , \sa_count[8][39] , 
	\sa_count[8][38] , \sa_count[8][37] , \sa_count[8][36] , 
	\sa_count[8][35] , \sa_count[8][34] , \sa_count[8][33] , 
	\sa_count[8][32] , \sa_count[8][31] , \sa_count[8][30] , 
	\sa_count[8][29] , \sa_count[8][28] , \sa_count[8][27] , 
	\sa_count[8][26] , \sa_count[8][25] , \sa_count[8][24] , 
	\sa_count[8][23] , \sa_count[8][22] , \sa_count[8][21] , 
	\sa_count[8][20] , \sa_count[8][19] , \sa_count[8][18] , 
	\sa_count[8][17] , \sa_count[8][16] , \sa_count[8][15] , 
	\sa_count[8][14] , \sa_count[8][13] , \sa_count[8][12] , 
	\sa_count[8][11] , \sa_count[8][10] , \sa_count[8][9] , 
	\sa_count[8][8] , \sa_count[8][7] , \sa_count[8][6] , 
	\sa_count[8][5] , \sa_count[8][4] , \sa_count[8][3] , 
	\sa_count[8][2] , \sa_count[8][1] , \sa_count[8][0] , 
	\sa_count[7][63] , \sa_count[7][62] , \sa_count[7][61] , 
	\sa_count[7][60] , \sa_count[7][59] , \sa_count[7][58] , 
	\sa_count[7][57] , \sa_count[7][56] , \sa_count[7][55] , 
	\sa_count[7][54] , \sa_count[7][53] , \sa_count[7][52] , 
	\sa_count[7][51] , \sa_count[7][50] , \sa_count[7][49] , 
	\sa_count[7][48] , \sa_count[7][47] , \sa_count[7][46] , 
	\sa_count[7][45] , \sa_count[7][44] , \sa_count[7][43] , 
	\sa_count[7][42] , \sa_count[7][41] , \sa_count[7][40] , 
	\sa_count[7][39] , \sa_count[7][38] , \sa_count[7][37] , 
	\sa_count[7][36] , \sa_count[7][35] , \sa_count[7][34] , 
	\sa_count[7][33] , \sa_count[7][32] , \sa_count[7][31] , 
	\sa_count[7][30] , \sa_count[7][29] , \sa_count[7][28] , 
	\sa_count[7][27] , \sa_count[7][26] , \sa_count[7][25] , 
	\sa_count[7][24] , \sa_count[7][23] , \sa_count[7][22] , 
	\sa_count[7][21] , \sa_count[7][20] , \sa_count[7][19] , 
	\sa_count[7][18] , \sa_count[7][17] , \sa_count[7][16] , 
	\sa_count[7][15] , \sa_count[7][14] , \sa_count[7][13] , 
	\sa_count[7][12] , \sa_count[7][11] , \sa_count[7][10] , 
	\sa_count[7][9] , \sa_count[7][8] , \sa_count[7][7] , 
	\sa_count[7][6] , \sa_count[7][5] , \sa_count[7][4] , 
	\sa_count[7][3] , \sa_count[7][2] , \sa_count[7][1] , 
	\sa_count[7][0] , \sa_count[6][63] , \sa_count[6][62] , 
	\sa_count[6][61] , \sa_count[6][60] , \sa_count[6][59] , 
	\sa_count[6][58] , \sa_count[6][57] , \sa_count[6][56] , 
	\sa_count[6][55] , \sa_count[6][54] , \sa_count[6][53] , 
	\sa_count[6][52] , \sa_count[6][51] , \sa_count[6][50] , 
	\sa_count[6][49] , \sa_count[6][48] , \sa_count[6][47] , 
	\sa_count[6][46] , \sa_count[6][45] , \sa_count[6][44] , 
	\sa_count[6][43] , \sa_count[6][42] , \sa_count[6][41] , 
	\sa_count[6][40] , \sa_count[6][39] , \sa_count[6][38] , 
	\sa_count[6][37] , \sa_count[6][36] , \sa_count[6][35] , 
	\sa_count[6][34] , \sa_count[6][33] , \sa_count[6][32] , 
	\sa_count[6][31] , \sa_count[6][30] , \sa_count[6][29] , 
	\sa_count[6][28] , \sa_count[6][27] , \sa_count[6][26] , 
	\sa_count[6][25] , \sa_count[6][24] , \sa_count[6][23] , 
	\sa_count[6][22] , \sa_count[6][21] , \sa_count[6][20] , 
	\sa_count[6][19] , \sa_count[6][18] , \sa_count[6][17] , 
	\sa_count[6][16] , \sa_count[6][15] , \sa_count[6][14] , 
	\sa_count[6][13] , \sa_count[6][12] , \sa_count[6][11] , 
	\sa_count[6][10] , \sa_count[6][9] , \sa_count[6][8] , 
	\sa_count[6][7] , \sa_count[6][6] , \sa_count[6][5] , 
	\sa_count[6][4] , \sa_count[6][3] , \sa_count[6][2] , 
	\sa_count[6][1] , \sa_count[6][0] , \sa_count[5][63] , 
	\sa_count[5][62] , \sa_count[5][61] , \sa_count[5][60] , 
	\sa_count[5][59] , \sa_count[5][58] , \sa_count[5][57] , 
	\sa_count[5][56] , \sa_count[5][55] , \sa_count[5][54] , 
	\sa_count[5][53] , \sa_count[5][52] , \sa_count[5][51] , 
	\sa_count[5][50] , \sa_count[5][49] , \sa_count[5][48] , 
	\sa_count[5][47] , \sa_count[5][46] , \sa_count[5][45] , 
	\sa_count[5][44] , \sa_count[5][43] , \sa_count[5][42] , 
	\sa_count[5][41] , \sa_count[5][40] , \sa_count[5][39] , 
	\sa_count[5][38] , \sa_count[5][37] , \sa_count[5][36] , 
	\sa_count[5][35] , \sa_count[5][34] , \sa_count[5][33] , 
	\sa_count[5][32] , \sa_count[5][31] , \sa_count[5][30] , 
	\sa_count[5][29] , \sa_count[5][28] , \sa_count[5][27] , 
	\sa_count[5][26] , \sa_count[5][25] , \sa_count[5][24] , 
	\sa_count[5][23] , \sa_count[5][22] , \sa_count[5][21] , 
	\sa_count[5][20] , \sa_count[5][19] , \sa_count[5][18] , 
	\sa_count[5][17] , \sa_count[5][16] , \sa_count[5][15] , 
	\sa_count[5][14] , \sa_count[5][13] , \sa_count[5][12] , 
	\sa_count[5][11] , \sa_count[5][10] , \sa_count[5][9] , 
	\sa_count[5][8] , \sa_count[5][7] , \sa_count[5][6] , 
	\sa_count[5][5] , \sa_count[5][4] , \sa_count[5][3] , 
	\sa_count[5][2] , \sa_count[5][1] , \sa_count[5][0] , 
	\sa_count[4][63] , \sa_count[4][62] , \sa_count[4][61] , 
	\sa_count[4][60] , \sa_count[4][59] , \sa_count[4][58] , 
	\sa_count[4][57] , \sa_count[4][56] , \sa_count[4][55] , 
	\sa_count[4][54] , \sa_count[4][53] , \sa_count[4][52] , 
	\sa_count[4][51] , \sa_count[4][50] , \sa_count[4][49] , 
	\sa_count[4][48] , \sa_count[4][47] , \sa_count[4][46] , 
	\sa_count[4][45] , \sa_count[4][44] , \sa_count[4][43] , 
	\sa_count[4][42] , \sa_count[4][41] , \sa_count[4][40] , 
	\sa_count[4][39] , \sa_count[4][38] , \sa_count[4][37] , 
	\sa_count[4][36] , \sa_count[4][35] , \sa_count[4][34] , 
	\sa_count[4][33] , \sa_count[4][32] , \sa_count[4][31] , 
	\sa_count[4][30] , \sa_count[4][29] , \sa_count[4][28] , 
	\sa_count[4][27] , \sa_count[4][26] , \sa_count[4][25] , 
	\sa_count[4][24] , \sa_count[4][23] , \sa_count[4][22] , 
	\sa_count[4][21] , \sa_count[4][20] , \sa_count[4][19] , 
	\sa_count[4][18] , \sa_count[4][17] , \sa_count[4][16] , 
	\sa_count[4][15] , \sa_count[4][14] , \sa_count[4][13] , 
	\sa_count[4][12] , \sa_count[4][11] , \sa_count[4][10] , 
	\sa_count[4][9] , \sa_count[4][8] , \sa_count[4][7] , 
	\sa_count[4][6] , \sa_count[4][5] , \sa_count[4][4] , 
	\sa_count[4][3] , \sa_count[4][2] , \sa_count[4][1] , 
	\sa_count[4][0] , \sa_count[3][63] , \sa_count[3][62] , 
	\sa_count[3][61] , \sa_count[3][60] , \sa_count[3][59] , 
	\sa_count[3][58] , \sa_count[3][57] , \sa_count[3][56] , 
	\sa_count[3][55] , \sa_count[3][54] , \sa_count[3][53] , 
	\sa_count[3][52] , \sa_count[3][51] , \sa_count[3][50] , 
	\sa_count[3][49] , \sa_count[3][48] , \sa_count[3][47] , 
	\sa_count[3][46] , \sa_count[3][45] , \sa_count[3][44] , 
	\sa_count[3][43] , \sa_count[3][42] , \sa_count[3][41] , 
	\sa_count[3][40] , \sa_count[3][39] , \sa_count[3][38] , 
	\sa_count[3][37] , \sa_count[3][36] , \sa_count[3][35] , 
	\sa_count[3][34] , \sa_count[3][33] , \sa_count[3][32] , 
	\sa_count[3][31] , \sa_count[3][30] , \sa_count[3][29] , 
	\sa_count[3][28] , \sa_count[3][27] , \sa_count[3][26] , 
	\sa_count[3][25] , \sa_count[3][24] , \sa_count[3][23] , 
	\sa_count[3][22] , \sa_count[3][21] , \sa_count[3][20] , 
	\sa_count[3][19] , \sa_count[3][18] , \sa_count[3][17] , 
	\sa_count[3][16] , \sa_count[3][15] , \sa_count[3][14] , 
	\sa_count[3][13] , \sa_count[3][12] , \sa_count[3][11] , 
	\sa_count[3][10] , \sa_count[3][9] , \sa_count[3][8] , 
	\sa_count[3][7] , \sa_count[3][6] , \sa_count[3][5] , 
	\sa_count[3][4] , \sa_count[3][3] , \sa_count[3][2] , 
	\sa_count[3][1] , \sa_count[3][0] , \sa_count[2][63] , 
	\sa_count[2][62] , \sa_count[2][61] , \sa_count[2][60] , 
	\sa_count[2][59] , \sa_count[2][58] , \sa_count[2][57] , 
	\sa_count[2][56] , \sa_count[2][55] , \sa_count[2][54] , 
	\sa_count[2][53] , \sa_count[2][52] , \sa_count[2][51] , 
	\sa_count[2][50] , \sa_count[2][49] , \sa_count[2][48] , 
	\sa_count[2][47] , \sa_count[2][46] , \sa_count[2][45] , 
	\sa_count[2][44] , \sa_count[2][43] , \sa_count[2][42] , 
	\sa_count[2][41] , \sa_count[2][40] , \sa_count[2][39] , 
	\sa_count[2][38] , \sa_count[2][37] , \sa_count[2][36] , 
	\sa_count[2][35] , \sa_count[2][34] , \sa_count[2][33] , 
	\sa_count[2][32] , \sa_count[2][31] , \sa_count[2][30] , 
	\sa_count[2][29] , \sa_count[2][28] , \sa_count[2][27] , 
	\sa_count[2][26] , \sa_count[2][25] , \sa_count[2][24] , 
	\sa_count[2][23] , \sa_count[2][22] , \sa_count[2][21] , 
	\sa_count[2][20] , \sa_count[2][19] , \sa_count[2][18] , 
	\sa_count[2][17] , \sa_count[2][16] , \sa_count[2][15] , 
	\sa_count[2][14] , \sa_count[2][13] , \sa_count[2][12] , 
	\sa_count[2][11] , \sa_count[2][10] , \sa_count[2][9] , 
	\sa_count[2][8] , \sa_count[2][7] , \sa_count[2][6] , 
	\sa_count[2][5] , \sa_count[2][4] , \sa_count[2][3] , 
	\sa_count[2][2] , \sa_count[2][1] , \sa_count[2][0] , 
	\sa_count[1][63] , \sa_count[1][62] , \sa_count[1][61] , 
	\sa_count[1][60] , \sa_count[1][59] , \sa_count[1][58] , 
	\sa_count[1][57] , \sa_count[1][56] , \sa_count[1][55] , 
	\sa_count[1][54] , \sa_count[1][53] , \sa_count[1][52] , 
	\sa_count[1][51] , \sa_count[1][50] , \sa_count[1][49] , 
	\sa_count[1][48] , \sa_count[1][47] , \sa_count[1][46] , 
	\sa_count[1][45] , \sa_count[1][44] , \sa_count[1][43] , 
	\sa_count[1][42] , \sa_count[1][41] , \sa_count[1][40] , 
	\sa_count[1][39] , \sa_count[1][38] , \sa_count[1][37] , 
	\sa_count[1][36] , \sa_count[1][35] , \sa_count[1][34] , 
	\sa_count[1][33] , \sa_count[1][32] , \sa_count[1][31] , 
	\sa_count[1][30] , \sa_count[1][29] , \sa_count[1][28] , 
	\sa_count[1][27] , \sa_count[1][26] , \sa_count[1][25] , 
	\sa_count[1][24] , \sa_count[1][23] , \sa_count[1][22] , 
	\sa_count[1][21] , \sa_count[1][20] , \sa_count[1][19] , 
	\sa_count[1][18] , \sa_count[1][17] , \sa_count[1][16] , 
	\sa_count[1][15] , \sa_count[1][14] , \sa_count[1][13] , 
	\sa_count[1][12] , \sa_count[1][11] , \sa_count[1][10] , 
	\sa_count[1][9] , \sa_count[1][8] , \sa_count[1][7] , 
	\sa_count[1][6] , \sa_count[1][5] , \sa_count[1][4] , 
	\sa_count[1][3] , \sa_count[1][2] , \sa_count[1][1] , 
	\sa_count[1][0] , \sa_count[0][63] , \sa_count[0][62] , 
	\sa_count[0][61] , \sa_count[0][60] , \sa_count[0][59] , 
	\sa_count[0][58] , \sa_count[0][57] , \sa_count[0][56] , 
	\sa_count[0][55] , \sa_count[0][54] , \sa_count[0][53] , 
	\sa_count[0][52] , \sa_count[0][51] , \sa_count[0][50] , 
	\sa_count[0][49] , \sa_count[0][48] , \sa_count[0][47] , 
	\sa_count[0][46] , \sa_count[0][45] , \sa_count[0][44] , 
	\sa_count[0][43] , \sa_count[0][42] , \sa_count[0][41] , 
	\sa_count[0][40] , \sa_count[0][39] , \sa_count[0][38] , 
	\sa_count[0][37] , \sa_count[0][36] , \sa_count[0][35] , 
	\sa_count[0][34] , \sa_count[0][33] , \sa_count[0][32] , 
	\sa_count[0][31] , \sa_count[0][30] , \sa_count[0][29] , 
	\sa_count[0][28] , \sa_count[0][27] , \sa_count[0][26] , 
	\sa_count[0][25] , \sa_count[0][24] , \sa_count[0][23] , 
	\sa_count[0][22] , \sa_count[0][21] , \sa_count[0][20] , 
	\sa_count[0][19] , \sa_count[0][18] , \sa_count[0][17] , 
	\sa_count[0][16] , \sa_count[0][15] , \sa_count[0][14] , 
	\sa_count[0][13] , \sa_count[0][12] , \sa_count[0][11] , 
	\sa_count[0][10] , \sa_count[0][9] , \sa_count[0][8] , 
	\sa_count[0][7] , \sa_count[0][6] , \sa_count[0][5] , 
	\sa_count[0][4] , \sa_count[0][3] , \sa_count[0][2] , 
	\sa_count[0][1] , \sa_count[0][0] }));
nx_roreg_indirect_access_xcm130 u_SA_SNAPSHOT ( .stat_code( 
	_zy_simnet_sa_snapshot_ia_status_772_w$[0:2]), .stat_datawords( 
	_zy_simnet_sa_snapshot_ia_status_773_w$[0:4]), .stat_addr( 
	_zy_simnet_sa_snapshot_ia_status_774_w$[0:4]), .capability_lst( 
	_zy_simnet_sa_snapshot_ia_capability_775_w$[0:15]), .capability_type( 
	_zy_simnet_sa_snapshot_ia_capability_776_w$[0:3]), .rd_dat( 
	_zy_simnet_sa_snapshot_ia_rdata_777_w$[0:63]), .clk( clk), .rst_n( 
	rst_n), .addr( _zy_simnet_reg_addr_778_w$[0:10]), .cmnd_op( 
	_zy_simnet_sa_snapshot_ia_config_779_w$[0:3]), .cmnd_addr( 
	_zy_simnet_sa_snapshot_ia_config_780_w$[0:4]), .wr_stb( 
	_zy_simnet_wr_stb_781_w$), .wr_dat( 
	_zy_simnet_sa_snapshot_ia_wdata_782_w$[0:63]), .mem_a( { 
	\sa_snapshot[31][63] , \sa_snapshot[31][62] , \sa_snapshot[31][61] , 
	\sa_snapshot[31][60] , \sa_snapshot[31][59] , \sa_snapshot[31][58] , 
	\sa_snapshot[31][57] , \sa_snapshot[31][56] , \sa_snapshot[31][55] , 
	\sa_snapshot[31][54] , \sa_snapshot[31][53] , \sa_snapshot[31][52] , 
	\sa_snapshot[31][51] , \sa_snapshot[31][50] , \sa_snapshot[31][49] , 
	\sa_snapshot[31][48] , \sa_snapshot[31][47] , \sa_snapshot[31][46] , 
	\sa_snapshot[31][45] , \sa_snapshot[31][44] , \sa_snapshot[31][43] , 
	\sa_snapshot[31][42] , \sa_snapshot[31][41] , \sa_snapshot[31][40] , 
	\sa_snapshot[31][39] , \sa_snapshot[31][38] , \sa_snapshot[31][37] , 
	\sa_snapshot[31][36] , \sa_snapshot[31][35] , \sa_snapshot[31][34] , 
	\sa_snapshot[31][33] , \sa_snapshot[31][32] , \sa_snapshot[31][31] , 
	\sa_snapshot[31][30] , \sa_snapshot[31][29] , \sa_snapshot[31][28] , 
	\sa_snapshot[31][27] , \sa_snapshot[31][26] , \sa_snapshot[31][25] , 
	\sa_snapshot[31][24] , \sa_snapshot[31][23] , \sa_snapshot[31][22] , 
	\sa_snapshot[31][21] , \sa_snapshot[31][20] , \sa_snapshot[31][19] , 
	\sa_snapshot[31][18] , \sa_snapshot[31][17] , \sa_snapshot[31][16] , 
	\sa_snapshot[31][15] , \sa_snapshot[31][14] , \sa_snapshot[31][13] , 
	\sa_snapshot[31][12] , \sa_snapshot[31][11] , \sa_snapshot[31][10] , 
	\sa_snapshot[31][9] , \sa_snapshot[31][8] , \sa_snapshot[31][7] , 
	\sa_snapshot[31][6] , \sa_snapshot[31][5] , \sa_snapshot[31][4] , 
	\sa_snapshot[31][3] , \sa_snapshot[31][2] , \sa_snapshot[31][1] , 
	\sa_snapshot[31][0] , \sa_snapshot[30][63] , \sa_snapshot[30][62] , 
	\sa_snapshot[30][61] , \sa_snapshot[30][60] , \sa_snapshot[30][59] , 
	\sa_snapshot[30][58] , \sa_snapshot[30][57] , \sa_snapshot[30][56] , 
	\sa_snapshot[30][55] , \sa_snapshot[30][54] , \sa_snapshot[30][53] , 
	\sa_snapshot[30][52] , \sa_snapshot[30][51] , \sa_snapshot[30][50] , 
	\sa_snapshot[30][49] , \sa_snapshot[30][48] , \sa_snapshot[30][47] , 
	\sa_snapshot[30][46] , \sa_snapshot[30][45] , \sa_snapshot[30][44] , 
	\sa_snapshot[30][43] , \sa_snapshot[30][42] , \sa_snapshot[30][41] , 
	\sa_snapshot[30][40] , \sa_snapshot[30][39] , \sa_snapshot[30][38] , 
	\sa_snapshot[30][37] , \sa_snapshot[30][36] , \sa_snapshot[30][35] , 
	\sa_snapshot[30][34] , \sa_snapshot[30][33] , \sa_snapshot[30][32] , 
	\sa_snapshot[30][31] , \sa_snapshot[30][30] , \sa_snapshot[30][29] , 
	\sa_snapshot[30][28] , \sa_snapshot[30][27] , \sa_snapshot[30][26] , 
	\sa_snapshot[30][25] , \sa_snapshot[30][24] , \sa_snapshot[30][23] , 
	\sa_snapshot[30][22] , \sa_snapshot[30][21] , \sa_snapshot[30][20] , 
	\sa_snapshot[30][19] , \sa_snapshot[30][18] , \sa_snapshot[30][17] , 
	\sa_snapshot[30][16] , \sa_snapshot[30][15] , \sa_snapshot[30][14] , 
	\sa_snapshot[30][13] , \sa_snapshot[30][12] , \sa_snapshot[30][11] , 
	\sa_snapshot[30][10] , \sa_snapshot[30][9] , \sa_snapshot[30][8] , 
	\sa_snapshot[30][7] , \sa_snapshot[30][6] , \sa_snapshot[30][5] , 
	\sa_snapshot[30][4] , \sa_snapshot[30][3] , \sa_snapshot[30][2] , 
	\sa_snapshot[30][1] , \sa_snapshot[30][0] , \sa_snapshot[29][63] , 
	\sa_snapshot[29][62] , \sa_snapshot[29][61] , \sa_snapshot[29][60] , 
	\sa_snapshot[29][59] , \sa_snapshot[29][58] , \sa_snapshot[29][57] , 
	\sa_snapshot[29][56] , \sa_snapshot[29][55] , \sa_snapshot[29][54] , 
	\sa_snapshot[29][53] , \sa_snapshot[29][52] , \sa_snapshot[29][51] , 
	\sa_snapshot[29][50] , \sa_snapshot[29][49] , \sa_snapshot[29][48] , 
	\sa_snapshot[29][47] , \sa_snapshot[29][46] , \sa_snapshot[29][45] , 
	\sa_snapshot[29][44] , \sa_snapshot[29][43] , \sa_snapshot[29][42] , 
	\sa_snapshot[29][41] , \sa_snapshot[29][40] , \sa_snapshot[29][39] , 
	\sa_snapshot[29][38] , \sa_snapshot[29][37] , \sa_snapshot[29][36] , 
	\sa_snapshot[29][35] , \sa_snapshot[29][34] , \sa_snapshot[29][33] , 
	\sa_snapshot[29][32] , \sa_snapshot[29][31] , \sa_snapshot[29][30] , 
	\sa_snapshot[29][29] , \sa_snapshot[29][28] , \sa_snapshot[29][27] , 
	\sa_snapshot[29][26] , \sa_snapshot[29][25] , \sa_snapshot[29][24] , 
	\sa_snapshot[29][23] , \sa_snapshot[29][22] , \sa_snapshot[29][21] , 
	\sa_snapshot[29][20] , \sa_snapshot[29][19] , \sa_snapshot[29][18] , 
	\sa_snapshot[29][17] , \sa_snapshot[29][16] , \sa_snapshot[29][15] , 
	\sa_snapshot[29][14] , \sa_snapshot[29][13] , \sa_snapshot[29][12] , 
	\sa_snapshot[29][11] , \sa_snapshot[29][10] , \sa_snapshot[29][9] , 
	\sa_snapshot[29][8] , \sa_snapshot[29][7] , \sa_snapshot[29][6] , 
	\sa_snapshot[29][5] , \sa_snapshot[29][4] , \sa_snapshot[29][3] , 
	\sa_snapshot[29][2] , \sa_snapshot[29][1] , \sa_snapshot[29][0] , 
	\sa_snapshot[28][63] , \sa_snapshot[28][62] , \sa_snapshot[28][61] , 
	\sa_snapshot[28][60] , \sa_snapshot[28][59] , \sa_snapshot[28][58] , 
	\sa_snapshot[28][57] , \sa_snapshot[28][56] , \sa_snapshot[28][55] , 
	\sa_snapshot[28][54] , \sa_snapshot[28][53] , \sa_snapshot[28][52] , 
	\sa_snapshot[28][51] , \sa_snapshot[28][50] , \sa_snapshot[28][49] , 
	\sa_snapshot[28][48] , \sa_snapshot[28][47] , \sa_snapshot[28][46] , 
	\sa_snapshot[28][45] , \sa_snapshot[28][44] , \sa_snapshot[28][43] , 
	\sa_snapshot[28][42] , \sa_snapshot[28][41] , \sa_snapshot[28][40] , 
	\sa_snapshot[28][39] , \sa_snapshot[28][38] , \sa_snapshot[28][37] , 
	\sa_snapshot[28][36] , \sa_snapshot[28][35] , \sa_snapshot[28][34] , 
	\sa_snapshot[28][33] , \sa_snapshot[28][32] , \sa_snapshot[28][31] , 
	\sa_snapshot[28][30] , \sa_snapshot[28][29] , \sa_snapshot[28][28] , 
	\sa_snapshot[28][27] , \sa_snapshot[28][26] , \sa_snapshot[28][25] , 
	\sa_snapshot[28][24] , \sa_snapshot[28][23] , \sa_snapshot[28][22] , 
	\sa_snapshot[28][21] , \sa_snapshot[28][20] , \sa_snapshot[28][19] , 
	\sa_snapshot[28][18] , \sa_snapshot[28][17] , \sa_snapshot[28][16] , 
	\sa_snapshot[28][15] , \sa_snapshot[28][14] , \sa_snapshot[28][13] , 
	\sa_snapshot[28][12] , \sa_snapshot[28][11] , \sa_snapshot[28][10] , 
	\sa_snapshot[28][9] , \sa_snapshot[28][8] , \sa_snapshot[28][7] , 
	\sa_snapshot[28][6] , \sa_snapshot[28][5] , \sa_snapshot[28][4] , 
	\sa_snapshot[28][3] , \sa_snapshot[28][2] , \sa_snapshot[28][1] , 
	\sa_snapshot[28][0] , \sa_snapshot[27][63] , \sa_snapshot[27][62] , 
	\sa_snapshot[27][61] , \sa_snapshot[27][60] , \sa_snapshot[27][59] , 
	\sa_snapshot[27][58] , \sa_snapshot[27][57] , \sa_snapshot[27][56] , 
	\sa_snapshot[27][55] , \sa_snapshot[27][54] , \sa_snapshot[27][53] , 
	\sa_snapshot[27][52] , \sa_snapshot[27][51] , \sa_snapshot[27][50] , 
	\sa_snapshot[27][49] , \sa_snapshot[27][48] , \sa_snapshot[27][47] , 
	\sa_snapshot[27][46] , \sa_snapshot[27][45] , \sa_snapshot[27][44] , 
	\sa_snapshot[27][43] , \sa_snapshot[27][42] , \sa_snapshot[27][41] , 
	\sa_snapshot[27][40] , \sa_snapshot[27][39] , \sa_snapshot[27][38] , 
	\sa_snapshot[27][37] , \sa_snapshot[27][36] , \sa_snapshot[27][35] , 
	\sa_snapshot[27][34] , \sa_snapshot[27][33] , \sa_snapshot[27][32] , 
	\sa_snapshot[27][31] , \sa_snapshot[27][30] , \sa_snapshot[27][29] , 
	\sa_snapshot[27][28] , \sa_snapshot[27][27] , \sa_snapshot[27][26] , 
	\sa_snapshot[27][25] , \sa_snapshot[27][24] , \sa_snapshot[27][23] , 
	\sa_snapshot[27][22] , \sa_snapshot[27][21] , \sa_snapshot[27][20] , 
	\sa_snapshot[27][19] , \sa_snapshot[27][18] , \sa_snapshot[27][17] , 
	\sa_snapshot[27][16] , \sa_snapshot[27][15] , \sa_snapshot[27][14] , 
	\sa_snapshot[27][13] , \sa_snapshot[27][12] , \sa_snapshot[27][11] , 
	\sa_snapshot[27][10] , \sa_snapshot[27][9] , \sa_snapshot[27][8] , 
	\sa_snapshot[27][7] , \sa_snapshot[27][6] , \sa_snapshot[27][5] , 
	\sa_snapshot[27][4] , \sa_snapshot[27][3] , \sa_snapshot[27][2] , 
	\sa_snapshot[27][1] , \sa_snapshot[27][0] , \sa_snapshot[26][63] , 
	\sa_snapshot[26][62] , \sa_snapshot[26][61] , \sa_snapshot[26][60] , 
	\sa_snapshot[26][59] , \sa_snapshot[26][58] , \sa_snapshot[26][57] , 
	\sa_snapshot[26][56] , \sa_snapshot[26][55] , \sa_snapshot[26][54] , 
	\sa_snapshot[26][53] , \sa_snapshot[26][52] , \sa_snapshot[26][51] , 
	\sa_snapshot[26][50] , \sa_snapshot[26][49] , \sa_snapshot[26][48] , 
	\sa_snapshot[26][47] , \sa_snapshot[26][46] , \sa_snapshot[26][45] , 
	\sa_snapshot[26][44] , \sa_snapshot[26][43] , \sa_snapshot[26][42] , 
	\sa_snapshot[26][41] , \sa_snapshot[26][40] , \sa_snapshot[26][39] , 
	\sa_snapshot[26][38] , \sa_snapshot[26][37] , \sa_snapshot[26][36] , 
	\sa_snapshot[26][35] , \sa_snapshot[26][34] , \sa_snapshot[26][33] , 
	\sa_snapshot[26][32] , \sa_snapshot[26][31] , \sa_snapshot[26][30] , 
	\sa_snapshot[26][29] , \sa_snapshot[26][28] , \sa_snapshot[26][27] , 
	\sa_snapshot[26][26] , \sa_snapshot[26][25] , \sa_snapshot[26][24] , 
	\sa_snapshot[26][23] , \sa_snapshot[26][22] , \sa_snapshot[26][21] , 
	\sa_snapshot[26][20] , \sa_snapshot[26][19] , \sa_snapshot[26][18] , 
	\sa_snapshot[26][17] , \sa_snapshot[26][16] , \sa_snapshot[26][15] , 
	\sa_snapshot[26][14] , \sa_snapshot[26][13] , \sa_snapshot[26][12] , 
	\sa_snapshot[26][11] , \sa_snapshot[26][10] , \sa_snapshot[26][9] , 
	\sa_snapshot[26][8] , \sa_snapshot[26][7] , \sa_snapshot[26][6] , 
	\sa_snapshot[26][5] , \sa_snapshot[26][4] , \sa_snapshot[26][3] , 
	\sa_snapshot[26][2] , \sa_snapshot[26][1] , \sa_snapshot[26][0] , 
	\sa_snapshot[25][63] , \sa_snapshot[25][62] , \sa_snapshot[25][61] , 
	\sa_snapshot[25][60] , \sa_snapshot[25][59] , \sa_snapshot[25][58] , 
	\sa_snapshot[25][57] , \sa_snapshot[25][56] , \sa_snapshot[25][55] , 
	\sa_snapshot[25][54] , \sa_snapshot[25][53] , \sa_snapshot[25][52] , 
	\sa_snapshot[25][51] , \sa_snapshot[25][50] , \sa_snapshot[25][49] , 
	\sa_snapshot[25][48] , \sa_snapshot[25][47] , \sa_snapshot[25][46] , 
	\sa_snapshot[25][45] , \sa_snapshot[25][44] , \sa_snapshot[25][43] , 
	\sa_snapshot[25][42] , \sa_snapshot[25][41] , \sa_snapshot[25][40] , 
	\sa_snapshot[25][39] , \sa_snapshot[25][38] , \sa_snapshot[25][37] , 
	\sa_snapshot[25][36] , \sa_snapshot[25][35] , \sa_snapshot[25][34] , 
	\sa_snapshot[25][33] , \sa_snapshot[25][32] , \sa_snapshot[25][31] , 
	\sa_snapshot[25][30] , \sa_snapshot[25][29] , \sa_snapshot[25][28] , 
	\sa_snapshot[25][27] , \sa_snapshot[25][26] , \sa_snapshot[25][25] , 
	\sa_snapshot[25][24] , \sa_snapshot[25][23] , \sa_snapshot[25][22] , 
	\sa_snapshot[25][21] , \sa_snapshot[25][20] , \sa_snapshot[25][19] , 
	\sa_snapshot[25][18] , \sa_snapshot[25][17] , \sa_snapshot[25][16] , 
	\sa_snapshot[25][15] , \sa_snapshot[25][14] , \sa_snapshot[25][13] , 
	\sa_snapshot[25][12] , \sa_snapshot[25][11] , \sa_snapshot[25][10] , 
	\sa_snapshot[25][9] , \sa_snapshot[25][8] , \sa_snapshot[25][7] , 
	\sa_snapshot[25][6] , \sa_snapshot[25][5] , \sa_snapshot[25][4] , 
	\sa_snapshot[25][3] , \sa_snapshot[25][2] , \sa_snapshot[25][1] , 
	\sa_snapshot[25][0] , \sa_snapshot[24][63] , \sa_snapshot[24][62] , 
	\sa_snapshot[24][61] , \sa_snapshot[24][60] , \sa_snapshot[24][59] , 
	\sa_snapshot[24][58] , \sa_snapshot[24][57] , \sa_snapshot[24][56] , 
	\sa_snapshot[24][55] , \sa_snapshot[24][54] , \sa_snapshot[24][53] , 
	\sa_snapshot[24][52] , \sa_snapshot[24][51] , \sa_snapshot[24][50] , 
	\sa_snapshot[24][49] , \sa_snapshot[24][48] , \sa_snapshot[24][47] , 
	\sa_snapshot[24][46] , \sa_snapshot[24][45] , \sa_snapshot[24][44] , 
	\sa_snapshot[24][43] , \sa_snapshot[24][42] , \sa_snapshot[24][41] , 
	\sa_snapshot[24][40] , \sa_snapshot[24][39] , \sa_snapshot[24][38] , 
	\sa_snapshot[24][37] , \sa_snapshot[24][36] , \sa_snapshot[24][35] , 
	\sa_snapshot[24][34] , \sa_snapshot[24][33] , \sa_snapshot[24][32] , 
	\sa_snapshot[24][31] , \sa_snapshot[24][30] , \sa_snapshot[24][29] , 
	\sa_snapshot[24][28] , \sa_snapshot[24][27] , \sa_snapshot[24][26] , 
	\sa_snapshot[24][25] , \sa_snapshot[24][24] , \sa_snapshot[24][23] , 
	\sa_snapshot[24][22] , \sa_snapshot[24][21] , \sa_snapshot[24][20] , 
	\sa_snapshot[24][19] , \sa_snapshot[24][18] , \sa_snapshot[24][17] , 
	\sa_snapshot[24][16] , \sa_snapshot[24][15] , \sa_snapshot[24][14] , 
	\sa_snapshot[24][13] , \sa_snapshot[24][12] , \sa_snapshot[24][11] , 
	\sa_snapshot[24][10] , \sa_snapshot[24][9] , \sa_snapshot[24][8] , 
	\sa_snapshot[24][7] , \sa_snapshot[24][6] , \sa_snapshot[24][5] , 
	\sa_snapshot[24][4] , \sa_snapshot[24][3] , \sa_snapshot[24][2] , 
	\sa_snapshot[24][1] , \sa_snapshot[24][0] , \sa_snapshot[23][63] , 
	\sa_snapshot[23][62] , \sa_snapshot[23][61] , \sa_snapshot[23][60] , 
	\sa_snapshot[23][59] , \sa_snapshot[23][58] , \sa_snapshot[23][57] , 
	\sa_snapshot[23][56] , \sa_snapshot[23][55] , \sa_snapshot[23][54] , 
	\sa_snapshot[23][53] , \sa_snapshot[23][52] , \sa_snapshot[23][51] , 
	\sa_snapshot[23][50] , \sa_snapshot[23][49] , \sa_snapshot[23][48] , 
	\sa_snapshot[23][47] , \sa_snapshot[23][46] , \sa_snapshot[23][45] , 
	\sa_snapshot[23][44] , \sa_snapshot[23][43] , \sa_snapshot[23][42] , 
	\sa_snapshot[23][41] , \sa_snapshot[23][40] , \sa_snapshot[23][39] , 
	\sa_snapshot[23][38] , \sa_snapshot[23][37] , \sa_snapshot[23][36] , 
	\sa_snapshot[23][35] , \sa_snapshot[23][34] , \sa_snapshot[23][33] , 
	\sa_snapshot[23][32] , \sa_snapshot[23][31] , \sa_snapshot[23][30] , 
	\sa_snapshot[23][29] , \sa_snapshot[23][28] , \sa_snapshot[23][27] , 
	\sa_snapshot[23][26] , \sa_snapshot[23][25] , \sa_snapshot[23][24] , 
	\sa_snapshot[23][23] , \sa_snapshot[23][22] , \sa_snapshot[23][21] , 
	\sa_snapshot[23][20] , \sa_snapshot[23][19] , \sa_snapshot[23][18] , 
	\sa_snapshot[23][17] , \sa_snapshot[23][16] , \sa_snapshot[23][15] , 
	\sa_snapshot[23][14] , \sa_snapshot[23][13] , \sa_snapshot[23][12] , 
	\sa_snapshot[23][11] , \sa_snapshot[23][10] , \sa_snapshot[23][9] , 
	\sa_snapshot[23][8] , \sa_snapshot[23][7] , \sa_snapshot[23][6] , 
	\sa_snapshot[23][5] , \sa_snapshot[23][4] , \sa_snapshot[23][3] , 
	\sa_snapshot[23][2] , \sa_snapshot[23][1] , \sa_snapshot[23][0] , 
	\sa_snapshot[22][63] , \sa_snapshot[22][62] , \sa_snapshot[22][61] , 
	\sa_snapshot[22][60] , \sa_snapshot[22][59] , \sa_snapshot[22][58] , 
	\sa_snapshot[22][57] , \sa_snapshot[22][56] , \sa_snapshot[22][55] , 
	\sa_snapshot[22][54] , \sa_snapshot[22][53] , \sa_snapshot[22][52] , 
	\sa_snapshot[22][51] , \sa_snapshot[22][50] , \sa_snapshot[22][49] , 
	\sa_snapshot[22][48] , \sa_snapshot[22][47] , \sa_snapshot[22][46] , 
	\sa_snapshot[22][45] , \sa_snapshot[22][44] , \sa_snapshot[22][43] , 
	\sa_snapshot[22][42] , \sa_snapshot[22][41] , \sa_snapshot[22][40] , 
	\sa_snapshot[22][39] , \sa_snapshot[22][38] , \sa_snapshot[22][37] , 
	\sa_snapshot[22][36] , \sa_snapshot[22][35] , \sa_snapshot[22][34] , 
	\sa_snapshot[22][33] , \sa_snapshot[22][32] , \sa_snapshot[22][31] , 
	\sa_snapshot[22][30] , \sa_snapshot[22][29] , \sa_snapshot[22][28] , 
	\sa_snapshot[22][27] , \sa_snapshot[22][26] , \sa_snapshot[22][25] , 
	\sa_snapshot[22][24] , \sa_snapshot[22][23] , \sa_snapshot[22][22] , 
	\sa_snapshot[22][21] , \sa_snapshot[22][20] , \sa_snapshot[22][19] , 
	\sa_snapshot[22][18] , \sa_snapshot[22][17] , \sa_snapshot[22][16] , 
	\sa_snapshot[22][15] , \sa_snapshot[22][14] , \sa_snapshot[22][13] , 
	\sa_snapshot[22][12] , \sa_snapshot[22][11] , \sa_snapshot[22][10] , 
	\sa_snapshot[22][9] , \sa_snapshot[22][8] , \sa_snapshot[22][7] , 
	\sa_snapshot[22][6] , \sa_snapshot[22][5] , \sa_snapshot[22][4] , 
	\sa_snapshot[22][3] , \sa_snapshot[22][2] , \sa_snapshot[22][1] , 
	\sa_snapshot[22][0] , \sa_snapshot[21][63] , \sa_snapshot[21][62] , 
	\sa_snapshot[21][61] , \sa_snapshot[21][60] , \sa_snapshot[21][59] , 
	\sa_snapshot[21][58] , \sa_snapshot[21][57] , \sa_snapshot[21][56] , 
	\sa_snapshot[21][55] , \sa_snapshot[21][54] , \sa_snapshot[21][53] , 
	\sa_snapshot[21][52] , \sa_snapshot[21][51] , \sa_snapshot[21][50] , 
	\sa_snapshot[21][49] , \sa_snapshot[21][48] , \sa_snapshot[21][47] , 
	\sa_snapshot[21][46] , \sa_snapshot[21][45] , \sa_snapshot[21][44] , 
	\sa_snapshot[21][43] , \sa_snapshot[21][42] , \sa_snapshot[21][41] , 
	\sa_snapshot[21][40] , \sa_snapshot[21][39] , \sa_snapshot[21][38] , 
	\sa_snapshot[21][37] , \sa_snapshot[21][36] , \sa_snapshot[21][35] , 
	\sa_snapshot[21][34] , \sa_snapshot[21][33] , \sa_snapshot[21][32] , 
	\sa_snapshot[21][31] , \sa_snapshot[21][30] , \sa_snapshot[21][29] , 
	\sa_snapshot[21][28] , \sa_snapshot[21][27] , \sa_snapshot[21][26] , 
	\sa_snapshot[21][25] , \sa_snapshot[21][24] , \sa_snapshot[21][23] , 
	\sa_snapshot[21][22] , \sa_snapshot[21][21] , \sa_snapshot[21][20] , 
	\sa_snapshot[21][19] , \sa_snapshot[21][18] , \sa_snapshot[21][17] , 
	\sa_snapshot[21][16] , \sa_snapshot[21][15] , \sa_snapshot[21][14] , 
	\sa_snapshot[21][13] , \sa_snapshot[21][12] , \sa_snapshot[21][11] , 
	\sa_snapshot[21][10] , \sa_snapshot[21][9] , \sa_snapshot[21][8] , 
	\sa_snapshot[21][7] , \sa_snapshot[21][6] , \sa_snapshot[21][5] , 
	\sa_snapshot[21][4] , \sa_snapshot[21][3] , \sa_snapshot[21][2] , 
	\sa_snapshot[21][1] , \sa_snapshot[21][0] , \sa_snapshot[20][63] , 
	\sa_snapshot[20][62] , \sa_snapshot[20][61] , \sa_snapshot[20][60] , 
	\sa_snapshot[20][59] , \sa_snapshot[20][58] , \sa_snapshot[20][57] , 
	\sa_snapshot[20][56] , \sa_snapshot[20][55] , \sa_snapshot[20][54] , 
	\sa_snapshot[20][53] , \sa_snapshot[20][52] , \sa_snapshot[20][51] , 
	\sa_snapshot[20][50] , \sa_snapshot[20][49] , \sa_snapshot[20][48] , 
	\sa_snapshot[20][47] , \sa_snapshot[20][46] , \sa_snapshot[20][45] , 
	\sa_snapshot[20][44] , \sa_snapshot[20][43] , \sa_snapshot[20][42] , 
	\sa_snapshot[20][41] , \sa_snapshot[20][40] , \sa_snapshot[20][39] , 
	\sa_snapshot[20][38] , \sa_snapshot[20][37] , \sa_snapshot[20][36] , 
	\sa_snapshot[20][35] , \sa_snapshot[20][34] , \sa_snapshot[20][33] , 
	\sa_snapshot[20][32] , \sa_snapshot[20][31] , \sa_snapshot[20][30] , 
	\sa_snapshot[20][29] , \sa_snapshot[20][28] , \sa_snapshot[20][27] , 
	\sa_snapshot[20][26] , \sa_snapshot[20][25] , \sa_snapshot[20][24] , 
	\sa_snapshot[20][23] , \sa_snapshot[20][22] , \sa_snapshot[20][21] , 
	\sa_snapshot[20][20] , \sa_snapshot[20][19] , \sa_snapshot[20][18] , 
	\sa_snapshot[20][17] , \sa_snapshot[20][16] , \sa_snapshot[20][15] , 
	\sa_snapshot[20][14] , \sa_snapshot[20][13] , \sa_snapshot[20][12] , 
	\sa_snapshot[20][11] , \sa_snapshot[20][10] , \sa_snapshot[20][9] , 
	\sa_snapshot[20][8] , \sa_snapshot[20][7] , \sa_snapshot[20][6] , 
	\sa_snapshot[20][5] , \sa_snapshot[20][4] , \sa_snapshot[20][3] , 
	\sa_snapshot[20][2] , \sa_snapshot[20][1] , \sa_snapshot[20][0] , 
	\sa_snapshot[19][63] , \sa_snapshot[19][62] , \sa_snapshot[19][61] , 
	\sa_snapshot[19][60] , \sa_snapshot[19][59] , \sa_snapshot[19][58] , 
	\sa_snapshot[19][57] , \sa_snapshot[19][56] , \sa_snapshot[19][55] , 
	\sa_snapshot[19][54] , \sa_snapshot[19][53] , \sa_snapshot[19][52] , 
	\sa_snapshot[19][51] , \sa_snapshot[19][50] , \sa_snapshot[19][49] , 
	\sa_snapshot[19][48] , \sa_snapshot[19][47] , \sa_snapshot[19][46] , 
	\sa_snapshot[19][45] , \sa_snapshot[19][44] , \sa_snapshot[19][43] , 
	\sa_snapshot[19][42] , \sa_snapshot[19][41] , \sa_snapshot[19][40] , 
	\sa_snapshot[19][39] , \sa_snapshot[19][38] , \sa_snapshot[19][37] , 
	\sa_snapshot[19][36] , \sa_snapshot[19][35] , \sa_snapshot[19][34] , 
	\sa_snapshot[19][33] , \sa_snapshot[19][32] , \sa_snapshot[19][31] , 
	\sa_snapshot[19][30] , \sa_snapshot[19][29] , \sa_snapshot[19][28] , 
	\sa_snapshot[19][27] , \sa_snapshot[19][26] , \sa_snapshot[19][25] , 
	\sa_snapshot[19][24] , \sa_snapshot[19][23] , \sa_snapshot[19][22] , 
	\sa_snapshot[19][21] , \sa_snapshot[19][20] , \sa_snapshot[19][19] , 
	\sa_snapshot[19][18] , \sa_snapshot[19][17] , \sa_snapshot[19][16] , 
	\sa_snapshot[19][15] , \sa_snapshot[19][14] , \sa_snapshot[19][13] , 
	\sa_snapshot[19][12] , \sa_snapshot[19][11] , \sa_snapshot[19][10] , 
	\sa_snapshot[19][9] , \sa_snapshot[19][8] , \sa_snapshot[19][7] , 
	\sa_snapshot[19][6] , \sa_snapshot[19][5] , \sa_snapshot[19][4] , 
	\sa_snapshot[19][3] , \sa_snapshot[19][2] , \sa_snapshot[19][1] , 
	\sa_snapshot[19][0] , \sa_snapshot[18][63] , \sa_snapshot[18][62] , 
	\sa_snapshot[18][61] , \sa_snapshot[18][60] , \sa_snapshot[18][59] , 
	\sa_snapshot[18][58] , \sa_snapshot[18][57] , \sa_snapshot[18][56] , 
	\sa_snapshot[18][55] , \sa_snapshot[18][54] , \sa_snapshot[18][53] , 
	\sa_snapshot[18][52] , \sa_snapshot[18][51] , \sa_snapshot[18][50] , 
	\sa_snapshot[18][49] , \sa_snapshot[18][48] , \sa_snapshot[18][47] , 
	\sa_snapshot[18][46] , \sa_snapshot[18][45] , \sa_snapshot[18][44] , 
	\sa_snapshot[18][43] , \sa_snapshot[18][42] , \sa_snapshot[18][41] , 
	\sa_snapshot[18][40] , \sa_snapshot[18][39] , \sa_snapshot[18][38] , 
	\sa_snapshot[18][37] , \sa_snapshot[18][36] , \sa_snapshot[18][35] , 
	\sa_snapshot[18][34] , \sa_snapshot[18][33] , \sa_snapshot[18][32] , 
	\sa_snapshot[18][31] , \sa_snapshot[18][30] , \sa_snapshot[18][29] , 
	\sa_snapshot[18][28] , \sa_snapshot[18][27] , \sa_snapshot[18][26] , 
	\sa_snapshot[18][25] , \sa_snapshot[18][24] , \sa_snapshot[18][23] , 
	\sa_snapshot[18][22] , \sa_snapshot[18][21] , \sa_snapshot[18][20] , 
	\sa_snapshot[18][19] , \sa_snapshot[18][18] , \sa_snapshot[18][17] , 
	\sa_snapshot[18][16] , \sa_snapshot[18][15] , \sa_snapshot[18][14] , 
	\sa_snapshot[18][13] , \sa_snapshot[18][12] , \sa_snapshot[18][11] , 
	\sa_snapshot[18][10] , \sa_snapshot[18][9] , \sa_snapshot[18][8] , 
	\sa_snapshot[18][7] , \sa_snapshot[18][6] , \sa_snapshot[18][5] , 
	\sa_snapshot[18][4] , \sa_snapshot[18][3] , \sa_snapshot[18][2] , 
	\sa_snapshot[18][1] , \sa_snapshot[18][0] , \sa_snapshot[17][63] , 
	\sa_snapshot[17][62] , \sa_snapshot[17][61] , \sa_snapshot[17][60] , 
	\sa_snapshot[17][59] , \sa_snapshot[17][58] , \sa_snapshot[17][57] , 
	\sa_snapshot[17][56] , \sa_snapshot[17][55] , \sa_snapshot[17][54] , 
	\sa_snapshot[17][53] , \sa_snapshot[17][52] , \sa_snapshot[17][51] , 
	\sa_snapshot[17][50] , \sa_snapshot[17][49] , \sa_snapshot[17][48] , 
	\sa_snapshot[17][47] , \sa_snapshot[17][46] , \sa_snapshot[17][45] , 
	\sa_snapshot[17][44] , \sa_snapshot[17][43] , \sa_snapshot[17][42] , 
	\sa_snapshot[17][41] , \sa_snapshot[17][40] , \sa_snapshot[17][39] , 
	\sa_snapshot[17][38] , \sa_snapshot[17][37] , \sa_snapshot[17][36] , 
	\sa_snapshot[17][35] , \sa_snapshot[17][34] , \sa_snapshot[17][33] , 
	\sa_snapshot[17][32] , \sa_snapshot[17][31] , \sa_snapshot[17][30] , 
	\sa_snapshot[17][29] , \sa_snapshot[17][28] , \sa_snapshot[17][27] , 
	\sa_snapshot[17][26] , \sa_snapshot[17][25] , \sa_snapshot[17][24] , 
	\sa_snapshot[17][23] , \sa_snapshot[17][22] , \sa_snapshot[17][21] , 
	\sa_snapshot[17][20] , \sa_snapshot[17][19] , \sa_snapshot[17][18] , 
	\sa_snapshot[17][17] , \sa_snapshot[17][16] , \sa_snapshot[17][15] , 
	\sa_snapshot[17][14] , \sa_snapshot[17][13] , \sa_snapshot[17][12] , 
	\sa_snapshot[17][11] , \sa_snapshot[17][10] , \sa_snapshot[17][9] , 
	\sa_snapshot[17][8] , \sa_snapshot[17][7] , \sa_snapshot[17][6] , 
	\sa_snapshot[17][5] , \sa_snapshot[17][4] , \sa_snapshot[17][3] , 
	\sa_snapshot[17][2] , \sa_snapshot[17][1] , \sa_snapshot[17][0] , 
	\sa_snapshot[16][63] , \sa_snapshot[16][62] , \sa_snapshot[16][61] , 
	\sa_snapshot[16][60] , \sa_snapshot[16][59] , \sa_snapshot[16][58] , 
	\sa_snapshot[16][57] , \sa_snapshot[16][56] , \sa_snapshot[16][55] , 
	\sa_snapshot[16][54] , \sa_snapshot[16][53] , \sa_snapshot[16][52] , 
	\sa_snapshot[16][51] , \sa_snapshot[16][50] , \sa_snapshot[16][49] , 
	\sa_snapshot[16][48] , \sa_snapshot[16][47] , \sa_snapshot[16][46] , 
	\sa_snapshot[16][45] , \sa_snapshot[16][44] , \sa_snapshot[16][43] , 
	\sa_snapshot[16][42] , \sa_snapshot[16][41] , \sa_snapshot[16][40] , 
	\sa_snapshot[16][39] , \sa_snapshot[16][38] , \sa_snapshot[16][37] , 
	\sa_snapshot[16][36] , \sa_snapshot[16][35] , \sa_snapshot[16][34] , 
	\sa_snapshot[16][33] , \sa_snapshot[16][32] , \sa_snapshot[16][31] , 
	\sa_snapshot[16][30] , \sa_snapshot[16][29] , \sa_snapshot[16][28] , 
	\sa_snapshot[16][27] , \sa_snapshot[16][26] , \sa_snapshot[16][25] , 
	\sa_snapshot[16][24] , \sa_snapshot[16][23] , \sa_snapshot[16][22] , 
	\sa_snapshot[16][21] , \sa_snapshot[16][20] , \sa_snapshot[16][19] , 
	\sa_snapshot[16][18] , \sa_snapshot[16][17] , \sa_snapshot[16][16] , 
	\sa_snapshot[16][15] , \sa_snapshot[16][14] , \sa_snapshot[16][13] , 
	\sa_snapshot[16][12] , \sa_snapshot[16][11] , \sa_snapshot[16][10] , 
	\sa_snapshot[16][9] , \sa_snapshot[16][8] , \sa_snapshot[16][7] , 
	\sa_snapshot[16][6] , \sa_snapshot[16][5] , \sa_snapshot[16][4] , 
	\sa_snapshot[16][3] , \sa_snapshot[16][2] , \sa_snapshot[16][1] , 
	\sa_snapshot[16][0] , \sa_snapshot[15][63] , \sa_snapshot[15][62] , 
	\sa_snapshot[15][61] , \sa_snapshot[15][60] , \sa_snapshot[15][59] , 
	\sa_snapshot[15][58] , \sa_snapshot[15][57] , \sa_snapshot[15][56] , 
	\sa_snapshot[15][55] , \sa_snapshot[15][54] , \sa_snapshot[15][53] , 
	\sa_snapshot[15][52] , \sa_snapshot[15][51] , \sa_snapshot[15][50] , 
	\sa_snapshot[15][49] , \sa_snapshot[15][48] , \sa_snapshot[15][47] , 
	\sa_snapshot[15][46] , \sa_snapshot[15][45] , \sa_snapshot[15][44] , 
	\sa_snapshot[15][43] , \sa_snapshot[15][42] , \sa_snapshot[15][41] , 
	\sa_snapshot[15][40] , \sa_snapshot[15][39] , \sa_snapshot[15][38] , 
	\sa_snapshot[15][37] , \sa_snapshot[15][36] , \sa_snapshot[15][35] , 
	\sa_snapshot[15][34] , \sa_snapshot[15][33] , \sa_snapshot[15][32] , 
	\sa_snapshot[15][31] , \sa_snapshot[15][30] , \sa_snapshot[15][29] , 
	\sa_snapshot[15][28] , \sa_snapshot[15][27] , \sa_snapshot[15][26] , 
	\sa_snapshot[15][25] , \sa_snapshot[15][24] , \sa_snapshot[15][23] , 
	\sa_snapshot[15][22] , \sa_snapshot[15][21] , \sa_snapshot[15][20] , 
	\sa_snapshot[15][19] , \sa_snapshot[15][18] , \sa_snapshot[15][17] , 
	\sa_snapshot[15][16] , \sa_snapshot[15][15] , \sa_snapshot[15][14] , 
	\sa_snapshot[15][13] , \sa_snapshot[15][12] , \sa_snapshot[15][11] , 
	\sa_snapshot[15][10] , \sa_snapshot[15][9] , \sa_snapshot[15][8] , 
	\sa_snapshot[15][7] , \sa_snapshot[15][6] , \sa_snapshot[15][5] , 
	\sa_snapshot[15][4] , \sa_snapshot[15][3] , \sa_snapshot[15][2] , 
	\sa_snapshot[15][1] , \sa_snapshot[15][0] , \sa_snapshot[14][63] , 
	\sa_snapshot[14][62] , \sa_snapshot[14][61] , \sa_snapshot[14][60] , 
	\sa_snapshot[14][59] , \sa_snapshot[14][58] , \sa_snapshot[14][57] , 
	\sa_snapshot[14][56] , \sa_snapshot[14][55] , \sa_snapshot[14][54] , 
	\sa_snapshot[14][53] , \sa_snapshot[14][52] , \sa_snapshot[14][51] , 
	\sa_snapshot[14][50] , \sa_snapshot[14][49] , \sa_snapshot[14][48] , 
	\sa_snapshot[14][47] , \sa_snapshot[14][46] , \sa_snapshot[14][45] , 
	\sa_snapshot[14][44] , \sa_snapshot[14][43] , \sa_snapshot[14][42] , 
	\sa_snapshot[14][41] , \sa_snapshot[14][40] , \sa_snapshot[14][39] , 
	\sa_snapshot[14][38] , \sa_snapshot[14][37] , \sa_snapshot[14][36] , 
	\sa_snapshot[14][35] , \sa_snapshot[14][34] , \sa_snapshot[14][33] , 
	\sa_snapshot[14][32] , \sa_snapshot[14][31] , \sa_snapshot[14][30] , 
	\sa_snapshot[14][29] , \sa_snapshot[14][28] , \sa_snapshot[14][27] , 
	\sa_snapshot[14][26] , \sa_snapshot[14][25] , \sa_snapshot[14][24] , 
	\sa_snapshot[14][23] , \sa_snapshot[14][22] , \sa_snapshot[14][21] , 
	\sa_snapshot[14][20] , \sa_snapshot[14][19] , \sa_snapshot[14][18] , 
	\sa_snapshot[14][17] , \sa_snapshot[14][16] , \sa_snapshot[14][15] , 
	\sa_snapshot[14][14] , \sa_snapshot[14][13] , \sa_snapshot[14][12] , 
	\sa_snapshot[14][11] , \sa_snapshot[14][10] , \sa_snapshot[14][9] , 
	\sa_snapshot[14][8] , \sa_snapshot[14][7] , \sa_snapshot[14][6] , 
	\sa_snapshot[14][5] , \sa_snapshot[14][4] , \sa_snapshot[14][3] , 
	\sa_snapshot[14][2] , \sa_snapshot[14][1] , \sa_snapshot[14][0] , 
	\sa_snapshot[13][63] , \sa_snapshot[13][62] , \sa_snapshot[13][61] , 
	\sa_snapshot[13][60] , \sa_snapshot[13][59] , \sa_snapshot[13][58] , 
	\sa_snapshot[13][57] , \sa_snapshot[13][56] , \sa_snapshot[13][55] , 
	\sa_snapshot[13][54] , \sa_snapshot[13][53] , \sa_snapshot[13][52] , 
	\sa_snapshot[13][51] , \sa_snapshot[13][50] , \sa_snapshot[13][49] , 
	\sa_snapshot[13][48] , \sa_snapshot[13][47] , \sa_snapshot[13][46] , 
	\sa_snapshot[13][45] , \sa_snapshot[13][44] , \sa_snapshot[13][43] , 
	\sa_snapshot[13][42] , \sa_snapshot[13][41] , \sa_snapshot[13][40] , 
	\sa_snapshot[13][39] , \sa_snapshot[13][38] , \sa_snapshot[13][37] , 
	\sa_snapshot[13][36] , \sa_snapshot[13][35] , \sa_snapshot[13][34] , 
	\sa_snapshot[13][33] , \sa_snapshot[13][32] , \sa_snapshot[13][31] , 
	\sa_snapshot[13][30] , \sa_snapshot[13][29] , \sa_snapshot[13][28] , 
	\sa_snapshot[13][27] , \sa_snapshot[13][26] , \sa_snapshot[13][25] , 
	\sa_snapshot[13][24] , \sa_snapshot[13][23] , \sa_snapshot[13][22] , 
	\sa_snapshot[13][21] , \sa_snapshot[13][20] , \sa_snapshot[13][19] , 
	\sa_snapshot[13][18] , \sa_snapshot[13][17] , \sa_snapshot[13][16] , 
	\sa_snapshot[13][15] , \sa_snapshot[13][14] , \sa_snapshot[13][13] , 
	\sa_snapshot[13][12] , \sa_snapshot[13][11] , \sa_snapshot[13][10] , 
	\sa_snapshot[13][9] , \sa_snapshot[13][8] , \sa_snapshot[13][7] , 
	\sa_snapshot[13][6] , \sa_snapshot[13][5] , \sa_snapshot[13][4] , 
	\sa_snapshot[13][3] , \sa_snapshot[13][2] , \sa_snapshot[13][1] , 
	\sa_snapshot[13][0] , \sa_snapshot[12][63] , \sa_snapshot[12][62] , 
	\sa_snapshot[12][61] , \sa_snapshot[12][60] , \sa_snapshot[12][59] , 
	\sa_snapshot[12][58] , \sa_snapshot[12][57] , \sa_snapshot[12][56] , 
	\sa_snapshot[12][55] , \sa_snapshot[12][54] , \sa_snapshot[12][53] , 
	\sa_snapshot[12][52] , \sa_snapshot[12][51] , \sa_snapshot[12][50] , 
	\sa_snapshot[12][49] , \sa_snapshot[12][48] , \sa_snapshot[12][47] , 
	\sa_snapshot[12][46] , \sa_snapshot[12][45] , \sa_snapshot[12][44] , 
	\sa_snapshot[12][43] , \sa_snapshot[12][42] , \sa_snapshot[12][41] , 
	\sa_snapshot[12][40] , \sa_snapshot[12][39] , \sa_snapshot[12][38] , 
	\sa_snapshot[12][37] , \sa_snapshot[12][36] , \sa_snapshot[12][35] , 
	\sa_snapshot[12][34] , \sa_snapshot[12][33] , \sa_snapshot[12][32] , 
	\sa_snapshot[12][31] , \sa_snapshot[12][30] , \sa_snapshot[12][29] , 
	\sa_snapshot[12][28] , \sa_snapshot[12][27] , \sa_snapshot[12][26] , 
	\sa_snapshot[12][25] , \sa_snapshot[12][24] , \sa_snapshot[12][23] , 
	\sa_snapshot[12][22] , \sa_snapshot[12][21] , \sa_snapshot[12][20] , 
	\sa_snapshot[12][19] , \sa_snapshot[12][18] , \sa_snapshot[12][17] , 
	\sa_snapshot[12][16] , \sa_snapshot[12][15] , \sa_snapshot[12][14] , 
	\sa_snapshot[12][13] , \sa_snapshot[12][12] , \sa_snapshot[12][11] , 
	\sa_snapshot[12][10] , \sa_snapshot[12][9] , \sa_snapshot[12][8] , 
	\sa_snapshot[12][7] , \sa_snapshot[12][6] , \sa_snapshot[12][5] , 
	\sa_snapshot[12][4] , \sa_snapshot[12][3] , \sa_snapshot[12][2] , 
	\sa_snapshot[12][1] , \sa_snapshot[12][0] , \sa_snapshot[11][63] , 
	\sa_snapshot[11][62] , \sa_snapshot[11][61] , \sa_snapshot[11][60] , 
	\sa_snapshot[11][59] , \sa_snapshot[11][58] , \sa_snapshot[11][57] , 
	\sa_snapshot[11][56] , \sa_snapshot[11][55] , \sa_snapshot[11][54] , 
	\sa_snapshot[11][53] , \sa_snapshot[11][52] , \sa_snapshot[11][51] , 
	\sa_snapshot[11][50] , \sa_snapshot[11][49] , \sa_snapshot[11][48] , 
	\sa_snapshot[11][47] , \sa_snapshot[11][46] , \sa_snapshot[11][45] , 
	\sa_snapshot[11][44] , \sa_snapshot[11][43] , \sa_snapshot[11][42] , 
	\sa_snapshot[11][41] , \sa_snapshot[11][40] , \sa_snapshot[11][39] , 
	\sa_snapshot[11][38] , \sa_snapshot[11][37] , \sa_snapshot[11][36] , 
	\sa_snapshot[11][35] , \sa_snapshot[11][34] , \sa_snapshot[11][33] , 
	\sa_snapshot[11][32] , \sa_snapshot[11][31] , \sa_snapshot[11][30] , 
	\sa_snapshot[11][29] , \sa_snapshot[11][28] , \sa_snapshot[11][27] , 
	\sa_snapshot[11][26] , \sa_snapshot[11][25] , \sa_snapshot[11][24] , 
	\sa_snapshot[11][23] , \sa_snapshot[11][22] , \sa_snapshot[11][21] , 
	\sa_snapshot[11][20] , \sa_snapshot[11][19] , \sa_snapshot[11][18] , 
	\sa_snapshot[11][17] , \sa_snapshot[11][16] , \sa_snapshot[11][15] , 
	\sa_snapshot[11][14] , \sa_snapshot[11][13] , \sa_snapshot[11][12] , 
	\sa_snapshot[11][11] , \sa_snapshot[11][10] , \sa_snapshot[11][9] , 
	\sa_snapshot[11][8] , \sa_snapshot[11][7] , \sa_snapshot[11][6] , 
	\sa_snapshot[11][5] , \sa_snapshot[11][4] , \sa_snapshot[11][3] , 
	\sa_snapshot[11][2] , \sa_snapshot[11][1] , \sa_snapshot[11][0] , 
	\sa_snapshot[10][63] , \sa_snapshot[10][62] , \sa_snapshot[10][61] , 
	\sa_snapshot[10][60] , \sa_snapshot[10][59] , \sa_snapshot[10][58] , 
	\sa_snapshot[10][57] , \sa_snapshot[10][56] , \sa_snapshot[10][55] , 
	\sa_snapshot[10][54] , \sa_snapshot[10][53] , \sa_snapshot[10][52] , 
	\sa_snapshot[10][51] , \sa_snapshot[10][50] , \sa_snapshot[10][49] , 
	\sa_snapshot[10][48] , \sa_snapshot[10][47] , \sa_snapshot[10][46] , 
	\sa_snapshot[10][45] , \sa_snapshot[10][44] , \sa_snapshot[10][43] , 
	\sa_snapshot[10][42] , \sa_snapshot[10][41] , \sa_snapshot[10][40] , 
	\sa_snapshot[10][39] , \sa_snapshot[10][38] , \sa_snapshot[10][37] , 
	\sa_snapshot[10][36] , \sa_snapshot[10][35] , \sa_snapshot[10][34] , 
	\sa_snapshot[10][33] , \sa_snapshot[10][32] , \sa_snapshot[10][31] , 
	\sa_snapshot[10][30] , \sa_snapshot[10][29] , \sa_snapshot[10][28] , 
	\sa_snapshot[10][27] , \sa_snapshot[10][26] , \sa_snapshot[10][25] , 
	\sa_snapshot[10][24] , \sa_snapshot[10][23] , \sa_snapshot[10][22] , 
	\sa_snapshot[10][21] , \sa_snapshot[10][20] , \sa_snapshot[10][19] , 
	\sa_snapshot[10][18] , \sa_snapshot[10][17] , \sa_snapshot[10][16] , 
	\sa_snapshot[10][15] , \sa_snapshot[10][14] , \sa_snapshot[10][13] , 
	\sa_snapshot[10][12] , \sa_snapshot[10][11] , \sa_snapshot[10][10] , 
	\sa_snapshot[10][9] , \sa_snapshot[10][8] , \sa_snapshot[10][7] , 
	\sa_snapshot[10][6] , \sa_snapshot[10][5] , \sa_snapshot[10][4] , 
	\sa_snapshot[10][3] , \sa_snapshot[10][2] , \sa_snapshot[10][1] , 
	\sa_snapshot[10][0] , \sa_snapshot[9][63] , \sa_snapshot[9][62] , 
	\sa_snapshot[9][61] , \sa_snapshot[9][60] , \sa_snapshot[9][59] , 
	\sa_snapshot[9][58] , \sa_snapshot[9][57] , \sa_snapshot[9][56] , 
	\sa_snapshot[9][55] , \sa_snapshot[9][54] , \sa_snapshot[9][53] , 
	\sa_snapshot[9][52] , \sa_snapshot[9][51] , \sa_snapshot[9][50] , 
	\sa_snapshot[9][49] , \sa_snapshot[9][48] , \sa_snapshot[9][47] , 
	\sa_snapshot[9][46] , \sa_snapshot[9][45] , \sa_snapshot[9][44] , 
	\sa_snapshot[9][43] , \sa_snapshot[9][42] , \sa_snapshot[9][41] , 
	\sa_snapshot[9][40] , \sa_snapshot[9][39] , \sa_snapshot[9][38] , 
	\sa_snapshot[9][37] , \sa_snapshot[9][36] , \sa_snapshot[9][35] , 
	\sa_snapshot[9][34] , \sa_snapshot[9][33] , \sa_snapshot[9][32] , 
	\sa_snapshot[9][31] , \sa_snapshot[9][30] , \sa_snapshot[9][29] , 
	\sa_snapshot[9][28] , \sa_snapshot[9][27] , \sa_snapshot[9][26] , 
	\sa_snapshot[9][25] , \sa_snapshot[9][24] , \sa_snapshot[9][23] , 
	\sa_snapshot[9][22] , \sa_snapshot[9][21] , \sa_snapshot[9][20] , 
	\sa_snapshot[9][19] , \sa_snapshot[9][18] , \sa_snapshot[9][17] , 
	\sa_snapshot[9][16] , \sa_snapshot[9][15] , \sa_snapshot[9][14] , 
	\sa_snapshot[9][13] , \sa_snapshot[9][12] , \sa_snapshot[9][11] , 
	\sa_snapshot[9][10] , \sa_snapshot[9][9] , \sa_snapshot[9][8] , 
	\sa_snapshot[9][7] , \sa_snapshot[9][6] , \sa_snapshot[9][5] , 
	\sa_snapshot[9][4] , \sa_snapshot[9][3] , \sa_snapshot[9][2] , 
	\sa_snapshot[9][1] , \sa_snapshot[9][0] , \sa_snapshot[8][63] , 
	\sa_snapshot[8][62] , \sa_snapshot[8][61] , \sa_snapshot[8][60] , 
	\sa_snapshot[8][59] , \sa_snapshot[8][58] , \sa_snapshot[8][57] , 
	\sa_snapshot[8][56] , \sa_snapshot[8][55] , \sa_snapshot[8][54] , 
	\sa_snapshot[8][53] , \sa_snapshot[8][52] , \sa_snapshot[8][51] , 
	\sa_snapshot[8][50] , \sa_snapshot[8][49] , \sa_snapshot[8][48] , 
	\sa_snapshot[8][47] , \sa_snapshot[8][46] , \sa_snapshot[8][45] , 
	\sa_snapshot[8][44] , \sa_snapshot[8][43] , \sa_snapshot[8][42] , 
	\sa_snapshot[8][41] , \sa_snapshot[8][40] , \sa_snapshot[8][39] , 
	\sa_snapshot[8][38] , \sa_snapshot[8][37] , \sa_snapshot[8][36] , 
	\sa_snapshot[8][35] , \sa_snapshot[8][34] , \sa_snapshot[8][33] , 
	\sa_snapshot[8][32] , \sa_snapshot[8][31] , \sa_snapshot[8][30] , 
	\sa_snapshot[8][29] , \sa_snapshot[8][28] , \sa_snapshot[8][27] , 
	\sa_snapshot[8][26] , \sa_snapshot[8][25] , \sa_snapshot[8][24] , 
	\sa_snapshot[8][23] , \sa_snapshot[8][22] , \sa_snapshot[8][21] , 
	\sa_snapshot[8][20] , \sa_snapshot[8][19] , \sa_snapshot[8][18] , 
	\sa_snapshot[8][17] , \sa_snapshot[8][16] , \sa_snapshot[8][15] , 
	\sa_snapshot[8][14] , \sa_snapshot[8][13] , \sa_snapshot[8][12] , 
	\sa_snapshot[8][11] , \sa_snapshot[8][10] , \sa_snapshot[8][9] , 
	\sa_snapshot[8][8] , \sa_snapshot[8][7] , \sa_snapshot[8][6] , 
	\sa_snapshot[8][5] , \sa_snapshot[8][4] , \sa_snapshot[8][3] , 
	\sa_snapshot[8][2] , \sa_snapshot[8][1] , \sa_snapshot[8][0] , 
	\sa_snapshot[7][63] , \sa_snapshot[7][62] , \sa_snapshot[7][61] , 
	\sa_snapshot[7][60] , \sa_snapshot[7][59] , \sa_snapshot[7][58] , 
	\sa_snapshot[7][57] , \sa_snapshot[7][56] , \sa_snapshot[7][55] , 
	\sa_snapshot[7][54] , \sa_snapshot[7][53] , \sa_snapshot[7][52] , 
	\sa_snapshot[7][51] , \sa_snapshot[7][50] , \sa_snapshot[7][49] , 
	\sa_snapshot[7][48] , \sa_snapshot[7][47] , \sa_snapshot[7][46] , 
	\sa_snapshot[7][45] , \sa_snapshot[7][44] , \sa_snapshot[7][43] , 
	\sa_snapshot[7][42] , \sa_snapshot[7][41] , \sa_snapshot[7][40] , 
	\sa_snapshot[7][39] , \sa_snapshot[7][38] , \sa_snapshot[7][37] , 
	\sa_snapshot[7][36] , \sa_snapshot[7][35] , \sa_snapshot[7][34] , 
	\sa_snapshot[7][33] , \sa_snapshot[7][32] , \sa_snapshot[7][31] , 
	\sa_snapshot[7][30] , \sa_snapshot[7][29] , \sa_snapshot[7][28] , 
	\sa_snapshot[7][27] , \sa_snapshot[7][26] , \sa_snapshot[7][25] , 
	\sa_snapshot[7][24] , \sa_snapshot[7][23] , \sa_snapshot[7][22] , 
	\sa_snapshot[7][21] , \sa_snapshot[7][20] , \sa_snapshot[7][19] , 
	\sa_snapshot[7][18] , \sa_snapshot[7][17] , \sa_snapshot[7][16] , 
	\sa_snapshot[7][15] , \sa_snapshot[7][14] , \sa_snapshot[7][13] , 
	\sa_snapshot[7][12] , \sa_snapshot[7][11] , \sa_snapshot[7][10] , 
	\sa_snapshot[7][9] , \sa_snapshot[7][8] , \sa_snapshot[7][7] , 
	\sa_snapshot[7][6] , \sa_snapshot[7][5] , \sa_snapshot[7][4] , 
	\sa_snapshot[7][3] , \sa_snapshot[7][2] , \sa_snapshot[7][1] , 
	\sa_snapshot[7][0] , \sa_snapshot[6][63] , \sa_snapshot[6][62] , 
	\sa_snapshot[6][61] , \sa_snapshot[6][60] , \sa_snapshot[6][59] , 
	\sa_snapshot[6][58] , \sa_snapshot[6][57] , \sa_snapshot[6][56] , 
	\sa_snapshot[6][55] , \sa_snapshot[6][54] , \sa_snapshot[6][53] , 
	\sa_snapshot[6][52] , \sa_snapshot[6][51] , \sa_snapshot[6][50] , 
	\sa_snapshot[6][49] , \sa_snapshot[6][48] , \sa_snapshot[6][47] , 
	\sa_snapshot[6][46] , \sa_snapshot[6][45] , \sa_snapshot[6][44] , 
	\sa_snapshot[6][43] , \sa_snapshot[6][42] , \sa_snapshot[6][41] , 
	\sa_snapshot[6][40] , \sa_snapshot[6][39] , \sa_snapshot[6][38] , 
	\sa_snapshot[6][37] , \sa_snapshot[6][36] , \sa_snapshot[6][35] , 
	\sa_snapshot[6][34] , \sa_snapshot[6][33] , \sa_snapshot[6][32] , 
	\sa_snapshot[6][31] , \sa_snapshot[6][30] , \sa_snapshot[6][29] , 
	\sa_snapshot[6][28] , \sa_snapshot[6][27] , \sa_snapshot[6][26] , 
	\sa_snapshot[6][25] , \sa_snapshot[6][24] , \sa_snapshot[6][23] , 
	\sa_snapshot[6][22] , \sa_snapshot[6][21] , \sa_snapshot[6][20] , 
	\sa_snapshot[6][19] , \sa_snapshot[6][18] , \sa_snapshot[6][17] , 
	\sa_snapshot[6][16] , \sa_snapshot[6][15] , \sa_snapshot[6][14] , 
	\sa_snapshot[6][13] , \sa_snapshot[6][12] , \sa_snapshot[6][11] , 
	\sa_snapshot[6][10] , \sa_snapshot[6][9] , \sa_snapshot[6][8] , 
	\sa_snapshot[6][7] , \sa_snapshot[6][6] , \sa_snapshot[6][5] , 
	\sa_snapshot[6][4] , \sa_snapshot[6][3] , \sa_snapshot[6][2] , 
	\sa_snapshot[6][1] , \sa_snapshot[6][0] , \sa_snapshot[5][63] , 
	\sa_snapshot[5][62] , \sa_snapshot[5][61] , \sa_snapshot[5][60] , 
	\sa_snapshot[5][59] , \sa_snapshot[5][58] , \sa_snapshot[5][57] , 
	\sa_snapshot[5][56] , \sa_snapshot[5][55] , \sa_snapshot[5][54] , 
	\sa_snapshot[5][53] , \sa_snapshot[5][52] , \sa_snapshot[5][51] , 
	\sa_snapshot[5][50] , \sa_snapshot[5][49] , \sa_snapshot[5][48] , 
	\sa_snapshot[5][47] , \sa_snapshot[5][46] , \sa_snapshot[5][45] , 
	\sa_snapshot[5][44] , \sa_snapshot[5][43] , \sa_snapshot[5][42] , 
	\sa_snapshot[5][41] , \sa_snapshot[5][40] , \sa_snapshot[5][39] , 
	\sa_snapshot[5][38] , \sa_snapshot[5][37] , \sa_snapshot[5][36] , 
	\sa_snapshot[5][35] , \sa_snapshot[5][34] , \sa_snapshot[5][33] , 
	\sa_snapshot[5][32] , \sa_snapshot[5][31] , \sa_snapshot[5][30] , 
	\sa_snapshot[5][29] , \sa_snapshot[5][28] , \sa_snapshot[5][27] , 
	\sa_snapshot[5][26] , \sa_snapshot[5][25] , \sa_snapshot[5][24] , 
	\sa_snapshot[5][23] , \sa_snapshot[5][22] , \sa_snapshot[5][21] , 
	\sa_snapshot[5][20] , \sa_snapshot[5][19] , \sa_snapshot[5][18] , 
	\sa_snapshot[5][17] , \sa_snapshot[5][16] , \sa_snapshot[5][15] , 
	\sa_snapshot[5][14] , \sa_snapshot[5][13] , \sa_snapshot[5][12] , 
	\sa_snapshot[5][11] , \sa_snapshot[5][10] , \sa_snapshot[5][9] , 
	\sa_snapshot[5][8] , \sa_snapshot[5][7] , \sa_snapshot[5][6] , 
	\sa_snapshot[5][5] , \sa_snapshot[5][4] , \sa_snapshot[5][3] , 
	\sa_snapshot[5][2] , \sa_snapshot[5][1] , \sa_snapshot[5][0] , 
	\sa_snapshot[4][63] , \sa_snapshot[4][62] , \sa_snapshot[4][61] , 
	\sa_snapshot[4][60] , \sa_snapshot[4][59] , \sa_snapshot[4][58] , 
	\sa_snapshot[4][57] , \sa_snapshot[4][56] , \sa_snapshot[4][55] , 
	\sa_snapshot[4][54] , \sa_snapshot[4][53] , \sa_snapshot[4][52] , 
	\sa_snapshot[4][51] , \sa_snapshot[4][50] , \sa_snapshot[4][49] , 
	\sa_snapshot[4][48] , \sa_snapshot[4][47] , \sa_snapshot[4][46] , 
	\sa_snapshot[4][45] , \sa_snapshot[4][44] , \sa_snapshot[4][43] , 
	\sa_snapshot[4][42] , \sa_snapshot[4][41] , \sa_snapshot[4][40] , 
	\sa_snapshot[4][39] , \sa_snapshot[4][38] , \sa_snapshot[4][37] , 
	\sa_snapshot[4][36] , \sa_snapshot[4][35] , \sa_snapshot[4][34] , 
	\sa_snapshot[4][33] , \sa_snapshot[4][32] , \sa_snapshot[4][31] , 
	\sa_snapshot[4][30] , \sa_snapshot[4][29] , \sa_snapshot[4][28] , 
	\sa_snapshot[4][27] , \sa_snapshot[4][26] , \sa_snapshot[4][25] , 
	\sa_snapshot[4][24] , \sa_snapshot[4][23] , \sa_snapshot[4][22] , 
	\sa_snapshot[4][21] , \sa_snapshot[4][20] , \sa_snapshot[4][19] , 
	\sa_snapshot[4][18] , \sa_snapshot[4][17] , \sa_snapshot[4][16] , 
	\sa_snapshot[4][15] , \sa_snapshot[4][14] , \sa_snapshot[4][13] , 
	\sa_snapshot[4][12] , \sa_snapshot[4][11] , \sa_snapshot[4][10] , 
	\sa_snapshot[4][9] , \sa_snapshot[4][8] , \sa_snapshot[4][7] , 
	\sa_snapshot[4][6] , \sa_snapshot[4][5] , \sa_snapshot[4][4] , 
	\sa_snapshot[4][3] , \sa_snapshot[4][2] , \sa_snapshot[4][1] , 
	\sa_snapshot[4][0] , \sa_snapshot[3][63] , \sa_snapshot[3][62] , 
	\sa_snapshot[3][61] , \sa_snapshot[3][60] , \sa_snapshot[3][59] , 
	\sa_snapshot[3][58] , \sa_snapshot[3][57] , \sa_snapshot[3][56] , 
	\sa_snapshot[3][55] , \sa_snapshot[3][54] , \sa_snapshot[3][53] , 
	\sa_snapshot[3][52] , \sa_snapshot[3][51] , \sa_snapshot[3][50] , 
	\sa_snapshot[3][49] , \sa_snapshot[3][48] , \sa_snapshot[3][47] , 
	\sa_snapshot[3][46] , \sa_snapshot[3][45] , \sa_snapshot[3][44] , 
	\sa_snapshot[3][43] , \sa_snapshot[3][42] , \sa_snapshot[3][41] , 
	\sa_snapshot[3][40] , \sa_snapshot[3][39] , \sa_snapshot[3][38] , 
	\sa_snapshot[3][37] , \sa_snapshot[3][36] , \sa_snapshot[3][35] , 
	\sa_snapshot[3][34] , \sa_snapshot[3][33] , \sa_snapshot[3][32] , 
	\sa_snapshot[3][31] , \sa_snapshot[3][30] , \sa_snapshot[3][29] , 
	\sa_snapshot[3][28] , \sa_snapshot[3][27] , \sa_snapshot[3][26] , 
	\sa_snapshot[3][25] , \sa_snapshot[3][24] , \sa_snapshot[3][23] , 
	\sa_snapshot[3][22] , \sa_snapshot[3][21] , \sa_snapshot[3][20] , 
	\sa_snapshot[3][19] , \sa_snapshot[3][18] , \sa_snapshot[3][17] , 
	\sa_snapshot[3][16] , \sa_snapshot[3][15] , \sa_snapshot[3][14] , 
	\sa_snapshot[3][13] , \sa_snapshot[3][12] , \sa_snapshot[3][11] , 
	\sa_snapshot[3][10] , \sa_snapshot[3][9] , \sa_snapshot[3][8] , 
	\sa_snapshot[3][7] , \sa_snapshot[3][6] , \sa_snapshot[3][5] , 
	\sa_snapshot[3][4] , \sa_snapshot[3][3] , \sa_snapshot[3][2] , 
	\sa_snapshot[3][1] , \sa_snapshot[3][0] , \sa_snapshot[2][63] , 
	\sa_snapshot[2][62] , \sa_snapshot[2][61] , \sa_snapshot[2][60] , 
	\sa_snapshot[2][59] , \sa_snapshot[2][58] , \sa_snapshot[2][57] , 
	\sa_snapshot[2][56] , \sa_snapshot[2][55] , \sa_snapshot[2][54] , 
	\sa_snapshot[2][53] , \sa_snapshot[2][52] , \sa_snapshot[2][51] , 
	\sa_snapshot[2][50] , \sa_snapshot[2][49] , \sa_snapshot[2][48] , 
	\sa_snapshot[2][47] , \sa_snapshot[2][46] , \sa_snapshot[2][45] , 
	\sa_snapshot[2][44] , \sa_snapshot[2][43] , \sa_snapshot[2][42] , 
	\sa_snapshot[2][41] , \sa_snapshot[2][40] , \sa_snapshot[2][39] , 
	\sa_snapshot[2][38] , \sa_snapshot[2][37] , \sa_snapshot[2][36] , 
	\sa_snapshot[2][35] , \sa_snapshot[2][34] , \sa_snapshot[2][33] , 
	\sa_snapshot[2][32] , \sa_snapshot[2][31] , \sa_snapshot[2][30] , 
	\sa_snapshot[2][29] , \sa_snapshot[2][28] , \sa_snapshot[2][27] , 
	\sa_snapshot[2][26] , \sa_snapshot[2][25] , \sa_snapshot[2][24] , 
	\sa_snapshot[2][23] , \sa_snapshot[2][22] , \sa_snapshot[2][21] , 
	\sa_snapshot[2][20] , \sa_snapshot[2][19] , \sa_snapshot[2][18] , 
	\sa_snapshot[2][17] , \sa_snapshot[2][16] , \sa_snapshot[2][15] , 
	\sa_snapshot[2][14] , \sa_snapshot[2][13] , \sa_snapshot[2][12] , 
	\sa_snapshot[2][11] , \sa_snapshot[2][10] , \sa_snapshot[2][9] , 
	\sa_snapshot[2][8] , \sa_snapshot[2][7] , \sa_snapshot[2][6] , 
	\sa_snapshot[2][5] , \sa_snapshot[2][4] , \sa_snapshot[2][3] , 
	\sa_snapshot[2][2] , \sa_snapshot[2][1] , \sa_snapshot[2][0] , 
	\sa_snapshot[1][63] , \sa_snapshot[1][62] , \sa_snapshot[1][61] , 
	\sa_snapshot[1][60] , \sa_snapshot[1][59] , \sa_snapshot[1][58] , 
	\sa_snapshot[1][57] , \sa_snapshot[1][56] , \sa_snapshot[1][55] , 
	\sa_snapshot[1][54] , \sa_snapshot[1][53] , \sa_snapshot[1][52] , 
	\sa_snapshot[1][51] , \sa_snapshot[1][50] , \sa_snapshot[1][49] , 
	\sa_snapshot[1][48] , \sa_snapshot[1][47] , \sa_snapshot[1][46] , 
	\sa_snapshot[1][45] , \sa_snapshot[1][44] , \sa_snapshot[1][43] , 
	\sa_snapshot[1][42] , \sa_snapshot[1][41] , \sa_snapshot[1][40] , 
	\sa_snapshot[1][39] , \sa_snapshot[1][38] , \sa_snapshot[1][37] , 
	\sa_snapshot[1][36] , \sa_snapshot[1][35] , \sa_snapshot[1][34] , 
	\sa_snapshot[1][33] , \sa_snapshot[1][32] , \sa_snapshot[1][31] , 
	\sa_snapshot[1][30] , \sa_snapshot[1][29] , \sa_snapshot[1][28] , 
	\sa_snapshot[1][27] , \sa_snapshot[1][26] , \sa_snapshot[1][25] , 
	\sa_snapshot[1][24] , \sa_snapshot[1][23] , \sa_snapshot[1][22] , 
	\sa_snapshot[1][21] , \sa_snapshot[1][20] , \sa_snapshot[1][19] , 
	\sa_snapshot[1][18] , \sa_snapshot[1][17] , \sa_snapshot[1][16] , 
	\sa_snapshot[1][15] , \sa_snapshot[1][14] , \sa_snapshot[1][13] , 
	\sa_snapshot[1][12] , \sa_snapshot[1][11] , \sa_snapshot[1][10] , 
	\sa_snapshot[1][9] , \sa_snapshot[1][8] , \sa_snapshot[1][7] , 
	\sa_snapshot[1][6] , \sa_snapshot[1][5] , \sa_snapshot[1][4] , 
	\sa_snapshot[1][3] , \sa_snapshot[1][2] , \sa_snapshot[1][1] , 
	\sa_snapshot[1][0] , \sa_snapshot[0][63] , \sa_snapshot[0][62] , 
	\sa_snapshot[0][61] , \sa_snapshot[0][60] , \sa_snapshot[0][59] , 
	\sa_snapshot[0][58] , \sa_snapshot[0][57] , \sa_snapshot[0][56] , 
	\sa_snapshot[0][55] , \sa_snapshot[0][54] , \sa_snapshot[0][53] , 
	\sa_snapshot[0][52] , \sa_snapshot[0][51] , \sa_snapshot[0][50] , 
	\sa_snapshot[0][49] , \sa_snapshot[0][48] , \sa_snapshot[0][47] , 
	\sa_snapshot[0][46] , \sa_snapshot[0][45] , \sa_snapshot[0][44] , 
	\sa_snapshot[0][43] , \sa_snapshot[0][42] , \sa_snapshot[0][41] , 
	\sa_snapshot[0][40] , \sa_snapshot[0][39] , \sa_snapshot[0][38] , 
	\sa_snapshot[0][37] , \sa_snapshot[0][36] , \sa_snapshot[0][35] , 
	\sa_snapshot[0][34] , \sa_snapshot[0][33] , \sa_snapshot[0][32] , 
	\sa_snapshot[0][31] , \sa_snapshot[0][30] , \sa_snapshot[0][29] , 
	\sa_snapshot[0][28] , \sa_snapshot[0][27] , \sa_snapshot[0][26] , 
	\sa_snapshot[0][25] , \sa_snapshot[0][24] , \sa_snapshot[0][23] , 
	\sa_snapshot[0][22] , \sa_snapshot[0][21] , \sa_snapshot[0][20] , 
	\sa_snapshot[0][19] , \sa_snapshot[0][18] , \sa_snapshot[0][17] , 
	\sa_snapshot[0][16] , \sa_snapshot[0][15] , \sa_snapshot[0][14] , 
	\sa_snapshot[0][13] , \sa_snapshot[0][12] , \sa_snapshot[0][11] , 
	\sa_snapshot[0][10] , \sa_snapshot[0][9] , \sa_snapshot[0][8] , 
	\sa_snapshot[0][7] , \sa_snapshot[0][6] , \sa_snapshot[0][5] , 
	\sa_snapshot[0][4] , \sa_snapshot[0][3] , \sa_snapshot[0][2] , 
	\sa_snapshot[0][1] , \sa_snapshot[0][0] }));
cr_kme_int_handler int_handler ( .kme_interrupt( kme_interrupt), 
	.interrupt_status( _zy_simnet_interrupt_status_757_w$[0:4]), 
	.suppress_key_tlvs( suppress_key_tlvs), .clk( clk), .rst_n( rst_n), 
	.set_drbg_expired_int( _zy_simnet_set_drbg_expired_int_758_w$), 
	.set_txc_bp_int( set_txc_bp_int), .set_gcm_tag_fail_int( 
	set_gcm_tag_fail_int), .set_key_tlv_miscmp_int( 
	set_key_tlv_miscmp_int), .set_tlv_bip2_error_int( 
	set_tlv_bip2_error_int), .cceip0_ism_mbe( 
	_zy_simnet_cceip0_ism_mbe_759_w$), .cceip1_ism_mbe( 
	_zy_simnet_cceip1_ism_mbe_760_w$), .cceip2_ism_mbe( 
	_zy_simnet_cceip2_ism_mbe_761_w$), .cceip3_ism_mbe( 
	_zy_simnet_cceip3_ism_mbe_762_w$), .cddip0_ism_mbe( 
	_zy_simnet_cddip0_ism_mbe_763_w$), .cddip1_ism_mbe( 
	_zy_simnet_cddip1_ism_mbe_764_w$), .cddip2_ism_mbe( 
	_zy_simnet_cddip2_ism_mbe_765_w$), .cddip3_ism_mbe( 
	_zy_simnet_cddip3_ism_mbe_766_w$), .kim_mbe( kim_mbe), .ckv_mbe( 
	ckv_mbe), .cceip_encrypt_mbe( cceip_encrypt_mbe), 
	.cceip_validate_mbe( cceip_validate_mbe), .cddip_decrypt_mbe( 
	cddip_decrypt_mbe), .axi_mbe( axi_mbe), .bimc_interrupt( 
	_zy_simnet_bimc_interrupt_767_w$), .wr_stb( 
	_zy_simnet_wr_stb_768_w$), .wr_data( _zy_simnet_wr_data_769_w$[0:31]), 
	.reg_addr( _zy_simnet_reg_addr_770_w$[0:10]), .o_interrupt_mask( 
	_zy_simnet_o_interrupt_mask_771_w$[0:4]));
bimc_master bimc_master ( .bimc_ecc_error( _zy_simnet_dio_718), 
	.bimc_interrupt( _zy_simnet_bimc_interrupt_719_w$), .bimc_odat( 
	_zy_simnet_kim_bimc_idat_720_w$), .bimc_osync( 
	_zy_simnet_kim_bimc_isync_721_w$), .bimc_rst_n( bimc_rst_n), .clk( 
	clk), .rst_n( rst_n), .bimc_idat( 
	_zy_simnet_axi_term_bimc_idat_722_w$), .bimc_isync( 
	_zy_simnet_axi_term_bimc_isync_723_w$), .o_bimc_monitor_mask( 
	_zy_simnet_o_bimc_monitor_mask_724_w$[0:6]), 
	.o_bimc_ecc_uncorrectable_error_cnt( 
	_zy_simnet_o_bimc_ecc_uncorrectable_error_cnt_725_w$[0:31]), 
	.o_bimc_ecc_correctable_error_cnt( 
	_zy_simnet_o_bimc_ecc_correctable_error_cnt_726_w$[0:31]), 
	.o_bimc_parity_error_cnt( 
	_zy_simnet_o_bimc_parity_error_cnt_727_w$[0:31]), 
	.o_bimc_global_config( _zy_simnet_o_bimc_global_config_728_w$[0:31]), 
	.o_bimc_eccpar_debug( _zy_simnet_o_bimc_eccpar_debug_729_w$[0:28]), 
	.o_bimc_cmd2( _zy_simnet_o_bimc_cmd2_730_w$[0:10]), .o_bimc_cmd1( 
	_zy_simnet_o_bimc_cmd1_731_w$[0:31]), .o_bimc_cmd0( 
	_zy_simnet_o_bimc_cmd0_732_w$[0:31]), .o_bimc_rxcmd2( 
	_zy_simnet_o_bimc_rxcmd2_733_w$[0:9]), .o_bimc_rxrsp2( 
	_zy_simnet_o_bimc_rxrsp2_734_w$[0:9]), .o_bimc_pollrsp2( 
	_zy_simnet_o_bimc_pollrsp2_735_w$[0:9]), .o_bimc_dbgcmd2( 
	_zy_simnet_o_bimc_dbgcmd2_736_w$[0:9]), .i_bimc_monitor( 
	_zy_simnet_bimc_monitor_737_w$[0:6]), 
	.i_bimc_ecc_uncorrectable_error_cnt( 
	_zy_simnet_bimc_ecc_uncorrectable_error_cnt_738_w$[0:31]), 
	.i_bimc_ecc_correctable_error_cnt( 
	_zy_simnet_bimc_ecc_correctable_error_cnt_739_w$[0:31]), 
	.i_bimc_parity_error_cnt( 
	_zy_simnet_bimc_parity_error_cnt_740_w$[0:31]), .i_bimc_global_config( 
	_zy_simnet_bimc_global_config_741_w$[0:31]), .i_bimc_memid( 
	_zy_simnet_bimc_memid_742_w$[0:11]), .i_bimc_eccpar_debug( 
	_zy_simnet_bimc_eccpar_debug_743_w$[0:28]), .i_bimc_cmd2( 
	_zy_simnet_bimc_cmd2_744_w$[0:10]), .i_bimc_rxcmd2( 
	_zy_simnet_bimc_rxcmd2_745_w$[0:9]), .i_bimc_rxcmd1( 
	_zy_simnet_bimc_rxcmd1_746_w$[0:31]), .i_bimc_rxcmd0( 
	_zy_simnet_bimc_rxcmd0_747_w$[0:31]), .i_bimc_rxrsp2( 
	_zy_simnet_bimc_rxrsp2_748_w$[0:9]), .i_bimc_rxrsp1( 
	_zy_simnet_bimc_rxrsp1_749_w$[0:31]), .i_bimc_rxrsp0( 
	_zy_simnet_bimc_rxrsp0_750_w$[0:31]), .i_bimc_pollrsp2( 
	_zy_simnet_bimc_pollrsp2_751_w$[0:9]), .i_bimc_pollrsp1( 
	_zy_simnet_bimc_pollrsp1_752_w$[0:31]), .i_bimc_pollrsp0( 
	_zy_simnet_bimc_pollrsp0_753_w$[0:31]), .i_bimc_dbgcmd2( 
	_zy_simnet_bimc_dbgcmd2_754_w$[0:9]), .i_bimc_dbgcmd1( 
	_zy_simnet_bimc_dbgcmd1_755_w$[0:31]), .i_bimc_dbgcmd0( 
	_zy_simnet_bimc_dbgcmd0_756_w$[0:31]));
cr_kme_drbg_reggen drbg_register_gen ( .set_drbg_expired_int( 
	_zy_simnet_set_drbg_expired_int_684_w$), .kdf_drbg_ctrl( 
	_zy_simnet_kdf_drbg_ctrl_685_w$[0:1]), .seed0_valid( seed0_valid), 
	.seed0_internal_state_key( seed0_internal_state_key[255:0]), 
	.seed0_internal_state_value( seed0_internal_state_value[127:0]), 
	.seed0_reseed_interval( seed0_reseed_interval[47:0]), 
	.seed1_valid( seed1_valid), .seed1_internal_state_key( 
	seed1_internal_state_key[255:0]), .seed1_internal_state_value( 
	seed1_internal_state_value[127:0]), .seed1_reseed_interval( 
	seed1_reseed_interval[47:0]), .clk( clk), .rst_n( rst_n), .wr_stb( 
	_zy_simnet_wr_stb_686_w$), .wr_data( _zy_simnet_wr_data_687_w$[0:31]), 
	.reg_addr( _zy_simnet_reg_addr_688_w$[0:10]), .o_kdf_drbg_ctrl( 
	_zy_simnet_o_kdf_drbg_ctrl_689_w$[0:1]), 
	.o_kdf_drbg_seed_0_reseed_interval_0( 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_0_690_w$[0:31]), 
	.o_kdf_drbg_seed_0_reseed_interval_1( 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_1_691_w$[0:15]), 
	.o_kdf_drbg_seed_0_state_key_127_96( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_127_96_692_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_159_128( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_159_128_693_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_191_160( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_191_160_694_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_223_192( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_223_192_695_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_255_224( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_255_224_696_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_31_0( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_31_0_697_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_63_32( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_63_32_698_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_95_64( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_95_64_699_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_value_127_96( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_127_96_700_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_value_31_0( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_31_0_701_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_value_63_32( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_63_32_702_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_value_95_64( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_95_64_703_w$[0:31]), 
	.o_kdf_drbg_seed_1_reseed_interval_0( 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_0_704_w$[0:31]), 
	.o_kdf_drbg_seed_1_reseed_interval_1( 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_1_705_w$[0:15]), 
	.o_kdf_drbg_seed_1_state_key_127_96( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_127_96_706_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_159_128( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_159_128_707_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_191_160( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_191_160_708_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_223_192( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_223_192_709_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_255_224( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_255_224_710_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_31_0( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_31_0_711_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_63_32( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_63_32_712_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_95_64( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_95_64_713_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_value_127_96( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_127_96_714_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_value_31_0( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_31_0_715_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_value_63_32( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_63_32_716_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_value_95_64( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_95_64_717_w$[0:31]), 
	.seed0_invalidate( seed0_invalidate), .seed1_invalidate( 
	seed1_invalidate));
nx_ram_1rw_indirect_access_xcm122 kim_indirect_access ( .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_663_w$[0:10]), .cmnd_op( 
	_zy_simnet_kim_cmnd_op_664_w$[0:3]), .cmnd_addr( 
	_zy_simnet_kim_cmnd_addr_665_w$[0:13]), .stat_code( 
	_zy_simnet_kim_stat_code_666_w$[0:2]), .stat_datawords( 
	_zy_simnet_kim_stat_datawords_667_w$[0:4]), .stat_addr( 
	_zy_simnet_kim_stat_addr_668_w$[0:13]), .capability_lst( 
	_zy_simnet_kim_capability_lst_669_w$[0:15]), .capability_type( 
	_zy_simnet_kim_capability_type_670_w$[0:3]), .wr_stb( 
	_zy_simnet_wr_stb_671_w$), .wr_dat( 
	_zy_simnet_kim_wr_dat_672_w$[0:37]), .rd_dat( 
	_zy_simnet_kim_rd_dat_673_w$[0:37]), .ovstb( ovstb), .lvm( lvm), 
	.mlvm( mlvm), .mrdten( _zy_simnet_cio_674), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_kim_bimc_isync_675_w$), 
	.bimc_idat( _zy_simnet_kim_bimc_idat_676_w$), .bimc_odat( 
	_zy_simnet_ckv_bimc_idat_677_w$), .bimc_osync( 
	_zy_simnet_ckv_bimc_isync_678_w$), .ro_uncorrectable_ecc_error( 
	kim_mbe), .hw_add( kim_addr[13:0]), .hw_we( _zy_simnet_cio_679), 
	.hw_bwe( _zy_simnet_cio_680[0:37]), .hw_cs( kim_rd), .hw_din( 
	_zy_simnet_cio_681[0:37]), .hw_dout( _zy_simnet_kim_dout_682_w$[0:37]), 
	.hw_yield( _zy_simnet_dio_683));
nx_ram_1rw_indirect_access_xcm123 ckv_indirect_access ( .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_643_w$[0:10]), .cmnd_op( 
	_zy_simnet_ckv_cmnd_op_644_w$[0:3]), .cmnd_addr( 
	_zy_simnet_ckv_cmnd_addr_645_w$[0:14]), .stat_code( 
	_zy_simnet_ckv_stat_code_646_w$[0:2]), .stat_datawords( 
	_zy_simnet_ckv_stat_datawords_647_w$[0:4]), .stat_addr( 
	_zy_simnet_ckv_stat_addr_648_w$[0:14]), .capability_lst( 
	_zy_simnet_ckv_capability_lst_649_w$[0:15]), .capability_type( 
	_zy_simnet_ckv_capability_type_650_w$[0:3]), .wr_stb( 
	_zy_simnet_wr_stb_651_w$), .wr_dat( 
	_zy_simnet_ckv_wr_dat_652_w$[0:63]), .rd_dat( 
	_zy_simnet_ckv_rd_dat_653_w$[0:63]), .ovstb( ovstb), .lvm( lvm), 
	.mlvm( mlvm), .mrdten( _zy_simnet_cio_654), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_ckv_bimc_isync_655_w$), 
	.bimc_idat( _zy_simnet_ckv_bimc_idat_656_w$), .bimc_odat( 
	_zy_simnet_cceip0_ism_bimc_idat_657_w$), .bimc_osync( 
	_zy_simnet_cceip0_ism_bimc_isync_658_w$), 
	.ro_uncorrectable_ecc_error( ckv_mbe), .hw_add( ckv_addr[14:0]), 
	.hw_we( _zy_simnet_cio_659), .hw_bwe( _zy_simnet_cio_660[0:63]), 
	.hw_cs( ckv_rd), .hw_din( _zy_simnet_cio_661[0:63]), .hw_dout( 
	ckv_dout[63:0]), .hw_yield( _zy_simnet_dio_662));
cr_kme_regfile_glue regfile_glue ( .ckv_cmnd_op( 
	_zy_simnet_ckv_cmnd_op_580_w$[0:3]), .ckv_cmnd_addr( 
	_zy_simnet_ckv_cmnd_addr_581_w$[0:14]), .ckv_wr_dat( 
	_zy_simnet_ckv_wr_dat_582_w$[0:63]), .ckv_ia_capability( 
	_zy_simnet_ckv_ia_capability_583_w$[0:19]), .ckv_ia_rdata_part0( 
	_zy_simnet_ckv_ia_rdata_part0_584_w$[0:31]), .ckv_ia_rdata_part1( 
	_zy_simnet_ckv_ia_rdata_part1_585_w$[0:31]), .ckv_ia_status( 
	_zy_simnet_ckv_ia_status_586_w$[0:22]), .kim_cmnd_op( 
	_zy_simnet_kim_cmnd_op_587_w$[0:3]), .kim_cmnd_addr( 
	_zy_simnet_kim_cmnd_addr_588_w$[0:13]), .kim_wr_dat( 
	_zy_simnet_kim_wr_dat_589_w$[0:37]), .kim_ia_capability( 
	_zy_simnet_kim_ia_capability_590_w$[0:19]), .kim_ia_rdata_part0( 
	_zy_simnet_kim_ia_rdata_part0_591_w$[0:20]), .kim_ia_rdata_part1( 
	_zy_simnet_kim_ia_rdata_part1_592_w$[0:16]), .kim_ia_status( 
	_zy_simnet_kim_ia_status_593_w$[0:21]), .engine_sticky_status( 
	_zy_simnet_engine_sticky_status_594_w$[0:7]), 
	.disable_ckv_kim_ism_reads( 
	_zy_simnet_disable_ckv_kim_ism_reads_595_w$), .send_kme_ib_beat( 
	_zy_simnet_send_kme_ib_beat_596_w$), .debug_kme_ib_tvalid( 
	debug_kme_ib_tvalid), .debug_kme_ib_tlast( debug_kme_ib_tlast), 
	.debug_kme_ib_tid( debug_kme_ib_tid[0]), .debug_kme_ib_tstrb( 
	debug_kme_ib_tstrb[7:0]), .debug_kme_ib_tuser( 
	debug_kme_ib_tuser[7:0]), .debug_kme_ib_tdata( 
	debug_kme_ib_tdata[63:0]), .kme_cceip0_ob_out( 
	_zy_simnet_kme_cceip0_ob_out_597_w$[0:82]), .kme_cceip1_ob_out( 
	_zy_simnet_kme_cceip1_ob_out_598_w$[0:82]), .kme_cceip2_ob_out( 
	_zy_simnet_kme_cceip2_ob_out_599_w$[0:82]), .kme_cceip3_ob_out( 
	_zy_simnet_kme_cceip3_ob_out_600_w$[0:82]), .kme_cddip0_ob_out( 
	_zy_simnet_kme_cddip0_ob_out_601_w$[0:82]), .kme_cddip1_ob_out( 
	_zy_simnet_kme_cddip1_ob_out_602_w$[0:82]), .kme_cddip2_ob_out( 
	_zy_simnet_kme_cddip2_ob_out_603_w$[0:82]), .kme_cddip3_ob_out( 
	_zy_simnet_kme_cddip3_ob_out_604_w$[0:82]), .cceip_encrypt_bimc_isync( 
	cceip_encrypt_bimc_isync), .cceip_encrypt_bimc_idat( 
	cceip_encrypt_bimc_idat), .cceip_validate_bimc_isync( 
	cceip_validate_bimc_isync), .cceip_validate_bimc_idat( 
	cceip_validate_bimc_idat), .cddip_decrypt_bimc_isync( 
	cddip_decrypt_bimc_isync), .cddip_decrypt_bimc_idat( 
	cddip_decrypt_bimc_idat), .axi_bimc_isync( axi_bimc_isync), 
	.axi_bimc_idat( axi_bimc_idat), .axi_term_bimc_isync( 
	_zy_simnet_axi_term_bimc_isync_605_w$), .axi_term_bimc_idat( 
	_zy_simnet_axi_term_bimc_idat_606_w$), .clk( clk), .rst_n( rst_n), 
	.ckv_stat_code( _zy_simnet_ckv_stat_code_607_w$[0:2]), 
	.ckv_stat_datawords( _zy_simnet_ckv_stat_datawords_608_w$[0:4]), 
	.ckv_stat_addr( _zy_simnet_ckv_stat_addr_609_w$[0:14]), 
	.ckv_capability_type( _zy_simnet_ckv_capability_type_610_w$[0:3]), 
	.ckv_capability_lst( _zy_simnet_ckv_capability_lst_611_w$[0:15]), 
	.ckv_rd_dat( _zy_simnet_ckv_rd_dat_612_w$[0:63]), .o_ckv_ia_config( 
	_zy_simnet_o_ckv_ia_config_613_w$[0:18]), .o_ckv_ia_wdata_part0( 
	_zy_simnet_o_ckv_ia_wdata_part0_614_w$[0:31]), .o_ckv_ia_wdata_part1( 
	_zy_simnet_o_ckv_ia_wdata_part1_615_w$[0:31]), .kim_stat_code( 
	_zy_simnet_kim_stat_code_616_w$[0:2]), .kim_stat_datawords( 
	_zy_simnet_kim_stat_datawords_617_w$[0:4]), .kim_stat_addr( 
	_zy_simnet_kim_stat_addr_618_w$[0:13]), .kim_capability_type( 
	_zy_simnet_kim_capability_type_619_w$[0:3]), .kim_capability_lst( 
	_zy_simnet_kim_capability_lst_620_w$[0:15]), .kim_rd_dat( 
	_zy_simnet_kim_rd_dat_621_w$[0:37]), .o_kim_ia_config( 
	_zy_simnet_o_kim_ia_config_622_w$[0:17]), .o_kim_ia_wdata_part0( 
	_zy_simnet_o_kim_ia_wdata_part0_623_w$[0:20]), .o_kim_ia_wdata_part1( 
	_zy_simnet_o_kim_ia_wdata_part1_624_w$[0:16]), 
	.set_rsm_is_backpressuring( set_rsm_is_backpressuring[7:0]), 
	.wr_stb( _zy_simnet_wr_stb_625_w$), .wr_data( 
	_zy_simnet_wr_data_626_w$[0:31]), .reg_addr( 
	_zy_simnet_reg_addr_627_w$[0:10]), .o_engine_sticky_status( 
	_zy_simnet_o_engine_sticky_status_628_w$[0:7]), 
	.o_disable_ckv_kim_ism_reads( 
	_zy_simnet_o_disable_ckv_kim_ism_reads_629_w$), .o_send_kme_ib_beat( 
	_zy_simnet_o_send_kme_ib_beat_630_w$), .cceip0_out_ia_wdata( 
	_zy_simnet_cceip0_out_ia_wdata_631_w$[0:95]), .debug_kme_ib_tready( 
	debug_kme_ib_tready), .tready_override( 
	_zy_simnet_tready_override_632_w$[0:8]), .kme_cceip0_ob_out_post( 
	_zy_simnet_kme_cceip0_ob_out_post_633_w$[0:82]), 
	.kme_cceip1_ob_out_post( 
	_zy_simnet_kme_cceip1_ob_out_post_634_w$[0:82]), 
	.kme_cceip2_ob_out_post( 
	_zy_simnet_kme_cceip2_ob_out_post_635_w$[0:82]), 
	.kme_cceip3_ob_out_post( 
	_zy_simnet_kme_cceip3_ob_out_post_636_w$[0:82]), 
	.kme_cddip0_ob_out_post( 
	_zy_simnet_kme_cddip0_ob_out_post_637_w$[0:82]), 
	.kme_cddip1_ob_out_post( 
	_zy_simnet_kme_cddip1_ob_out_post_638_w$[0:82]), 
	.kme_cddip2_ob_out_post( 
	_zy_simnet_kme_cddip2_ob_out_post_639_w$[0:82]), 
	.kme_cddip3_ob_out_post( 
	_zy_simnet_kme_cddip3_ob_out_post_640_w$[0:82]), .cddip3_ism_osync( 
	_zy_simnet_cddip3_ism_osync_641_w$), .cddip3_ism_odat( 
	_zy_simnet_cddip3_ism_odat_642_w$), .cceip_encrypt_bimc_osync( 
	cceip_encrypt_bimc_osync), .cceip_encrypt_bimc_odat( 
	cceip_encrypt_bimc_odat), .cceip_validate_bimc_osync( 
	cceip_validate_bimc_osync), .cceip_validate_bimc_odat( 
	cceip_validate_bimc_odat), .cddip_decrypt_bimc_osync( 
	cddip_decrypt_bimc_osync), .cddip_decrypt_bimc_odat( 
	cddip_decrypt_bimc_odat), .axi_bimc_osync( axi_bimc_osync), 
	.axi_bimc_odat( axi_bimc_odat));
nx_interface_monitor_xcm97 u_nx_interface_monitor_cddip3 ( .stat_code( 
	_zy_simnet_cddip3_out_ia_status_556_w$[0:2]), .stat_datawords( 
	_zy_simnet_cddip3_out_ia_status_557_w$[0:4]), .stat_addr( 
	_zy_simnet_cddip3_out_ia_status_558_w$[0:8]), .capability_lst( 
	_zy_simnet_cddip3_out_ia_capability_559_w$[0:15]), .capability_type( 
	_zy_simnet_cddip3_out_ia_capability_560_w$[0:3]), .rd_dat( 
	_zy_simnet_cddip3_out_ia_rdata_561_w$[0:95]), .bimc_odat( 
	_zy_simnet_cddip3_ism_odat_562_w$), .bimc_osync( 
	_zy_simnet_cddip3_ism_osync_563_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_cddip3_ism_mbe_564_w$), .im_rdy( 
	_zy_simnet_cddip3_im_rdy_565_w$), .im_available( 
	_zy_simnet_im_available_kme_cddip3_566_w$[0:1]), .im_status( 
	_zy_simnet_cddip3_out_im_status_567_w$[0:11]), .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_568_w$[0:10]), .cmnd_op( 
	_zy_simnet_cddip3_out_ia_config_569_w$[0:3]), .cmnd_addr( 
	_zy_simnet_cddip3_out_ia_config_570_w$[0:8]), .wr_stb( 
	_zy_simnet_wr_stb_571_w$), .wr_dat( 
	_zy_simnet_cddip3_out_ia_wdata_572_w$[0:95]), .ovstb( ovstb), .lvm( 
	lvm), .mlvm( mlvm), .mrdten( _zy_simnet_cio_573), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_cddip3_ism_isync_574_w$), 
	.bimc_idat( _zy_simnet_cddip3_ism_idat_575_w$), .im_din( 
	_zy_simnet_cddip3_im_din_576_w$[0:95]), .im_vld( 
	_zy_simnet_cddip3_im_vld_577_w$), .im_consumed( 
	_zy_simnet_im_consumed_kme_cddip3_578_w$[0:1]), .im_config( 
	_zy_simnet_cddip3_out_im_config_579_w$[0:11]));
nx_interface_monitor_xcm98 u_nx_interface_monitor_cddip2 ( .stat_code( 
	_zy_simnet_cddip2_out_ia_status_532_w$[0:2]), .stat_datawords( 
	_zy_simnet_cddip2_out_ia_status_533_w$[0:4]), .stat_addr( 
	_zy_simnet_cddip2_out_ia_status_534_w$[0:8]), .capability_lst( 
	_zy_simnet_cddip2_out_ia_capability_535_w$[0:15]), .capability_type( 
	_zy_simnet_cddip2_out_ia_capability_536_w$[0:3]), .rd_dat( 
	_zy_simnet_cddip2_out_ia_rdata_537_w$[0:95]), .bimc_odat( 
	_zy_simnet_cddip3_ism_idat_538_w$), .bimc_osync( 
	_zy_simnet_cddip3_ism_isync_539_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_cddip2_ism_mbe_540_w$), .im_rdy( 
	_zy_simnet_cddip2_im_rdy_541_w$), .im_available( 
	_zy_simnet_im_available_kme_cddip2_542_w$[0:1]), .im_status( 
	_zy_simnet_cddip2_out_im_status_543_w$[0:11]), .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_544_w$[0:10]), .cmnd_op( 
	_zy_simnet_cddip2_out_ia_config_545_w$[0:3]), .cmnd_addr( 
	_zy_simnet_cddip2_out_ia_config_546_w$[0:8]), .wr_stb( 
	_zy_simnet_wr_stb_547_w$), .wr_dat( 
	_zy_simnet_cddip2_out_ia_wdata_548_w$[0:95]), .ovstb( ovstb), .lvm( 
	lvm), .mlvm( mlvm), .mrdten( _zy_simnet_cio_549), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_cddip2_ism_isync_550_w$), 
	.bimc_idat( _zy_simnet_cddip2_ism_idat_551_w$), .im_din( 
	_zy_simnet_cddip2_im_din_552_w$[0:95]), .im_vld( 
	_zy_simnet_cddip2_im_vld_553_w$), .im_consumed( 
	_zy_simnet_im_consumed_kme_cddip2_554_w$[0:1]), .im_config( 
	_zy_simnet_cddip2_out_im_config_555_w$[0:11]));
nx_interface_monitor_xcm99 u_nx_interface_monitor_cddip1 ( .stat_code( 
	_zy_simnet_cddip1_out_ia_status_508_w$[0:2]), .stat_datawords( 
	_zy_simnet_cddip1_out_ia_status_509_w$[0:4]), .stat_addr( 
	_zy_simnet_cddip1_out_ia_status_510_w$[0:8]), .capability_lst( 
	_zy_simnet_cddip1_out_ia_capability_511_w$[0:15]), .capability_type( 
	_zy_simnet_cddip1_out_ia_capability_512_w$[0:3]), .rd_dat( 
	_zy_simnet_cddip1_out_ia_rdata_513_w$[0:95]), .bimc_odat( 
	_zy_simnet_cddip2_ism_idat_514_w$), .bimc_osync( 
	_zy_simnet_cddip2_ism_isync_515_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_cddip1_ism_mbe_516_w$), .im_rdy( 
	_zy_simnet_cddip1_im_rdy_517_w$), .im_available( 
	_zy_simnet_im_available_kme_cddip1_518_w$[0:1]), .im_status( 
	_zy_simnet_cddip1_out_im_status_519_w$[0:11]), .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_520_w$[0:10]), .cmnd_op( 
	_zy_simnet_cddip1_out_ia_config_521_w$[0:3]), .cmnd_addr( 
	_zy_simnet_cddip1_out_ia_config_522_w$[0:8]), .wr_stb( 
	_zy_simnet_wr_stb_523_w$), .wr_dat( 
	_zy_simnet_cddip1_out_ia_wdata_524_w$[0:95]), .ovstb( ovstb), .lvm( 
	lvm), .mlvm( mlvm), .mrdten( _zy_simnet_cio_525), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_cddip1_ism_isync_526_w$), 
	.bimc_idat( _zy_simnet_cddip1_ism_idat_527_w$), .im_din( 
	_zy_simnet_cddip1_im_din_528_w$[0:95]), .im_vld( 
	_zy_simnet_cddip1_im_vld_529_w$), .im_consumed( 
	_zy_simnet_im_consumed_kme_cddip1_530_w$[0:1]), .im_config( 
	_zy_simnet_cddip1_out_im_config_531_w$[0:11]));
nx_interface_monitor_xcm100 u_nx_interface_monitor_cddip0 ( .stat_code( 
	_zy_simnet_cddip0_out_ia_status_484_w$[0:2]), .stat_datawords( 
	_zy_simnet_cddip0_out_ia_status_485_w$[0:4]), .stat_addr( 
	_zy_simnet_cddip0_out_ia_status_486_w$[0:8]), .capability_lst( 
	_zy_simnet_cddip0_out_ia_capability_487_w$[0:15]), .capability_type( 
	_zy_simnet_cddip0_out_ia_capability_488_w$[0:3]), .rd_dat( 
	_zy_simnet_cddip0_out_ia_rdata_489_w$[0:95]), .bimc_odat( 
	_zy_simnet_cddip1_ism_idat_490_w$), .bimc_osync( 
	_zy_simnet_cddip1_ism_isync_491_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_cddip0_ism_mbe_492_w$), .im_rdy( 
	_zy_simnet_cddip0_im_rdy_493_w$), .im_available( 
	_zy_simnet_im_available_kme_cddip0_494_w$[0:1]), .im_status( 
	_zy_simnet_cddip0_out_im_status_495_w$[0:11]), .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_496_w$[0:10]), .cmnd_op( 
	_zy_simnet_cddip0_out_ia_config_497_w$[0:3]), .cmnd_addr( 
	_zy_simnet_cddip0_out_ia_config_498_w$[0:8]), .wr_stb( 
	_zy_simnet_wr_stb_499_w$), .wr_dat( 
	_zy_simnet_cddip0_out_ia_wdata_500_w$[0:95]), .ovstb( ovstb), .lvm( 
	lvm), .mlvm( mlvm), .mrdten( _zy_simnet_cio_501), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_cddip0_ism_isync_502_w$), 
	.bimc_idat( _zy_simnet_cddip0_ism_idat_503_w$), .im_din( 
	_zy_simnet_cddip0_im_din_504_w$[0:95]), .im_vld( 
	_zy_simnet_cddip0_im_vld_505_w$), .im_consumed( 
	_zy_simnet_im_consumed_kme_cddip0_506_w$[0:1]), .im_config( 
	_zy_simnet_cddip0_out_im_config_507_w$[0:11]));
nx_interface_monitor_xcm101 u_nx_interface_monitor_cceip3 ( .stat_code( 
	_zy_simnet_cceip3_out_ia_status_460_w$[0:2]), .stat_datawords( 
	_zy_simnet_cceip3_out_ia_status_461_w$[0:4]), .stat_addr( 
	_zy_simnet_cceip3_out_ia_status_462_w$[0:8]), .capability_lst( 
	_zy_simnet_cceip3_out_ia_capability_463_w$[0:15]), .capability_type( 
	_zy_simnet_cceip3_out_ia_capability_464_w$[0:3]), .rd_dat( 
	_zy_simnet_cceip3_out_ia_rdata_465_w$[0:95]), .bimc_odat( 
	_zy_simnet_cddip0_ism_idat_466_w$), .bimc_osync( 
	_zy_simnet_cddip0_ism_isync_467_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_cceip3_ism_mbe_468_w$), .im_rdy( 
	_zy_simnet_cceip3_im_rdy_469_w$), .im_available( 
	_zy_simnet_im_available_kme_cceip3_470_w$[0:1]), .im_status( 
	_zy_simnet_cceip3_out_im_status_471_w$[0:11]), .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_472_w$[0:10]), .cmnd_op( 
	_zy_simnet_cceip3_out_ia_config_473_w$[0:3]), .cmnd_addr( 
	_zy_simnet_cceip3_out_ia_config_474_w$[0:8]), .wr_stb( 
	_zy_simnet_wr_stb_475_w$), .wr_dat( 
	_zy_simnet_cceip3_out_ia_wdata_476_w$[0:95]), .ovstb( ovstb), .lvm( 
	lvm), .mlvm( mlvm), .mrdten( _zy_simnet_cio_477), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_cceip3_ism_isync_478_w$), 
	.bimc_idat( _zy_simnet_cceip3_ism_idat_479_w$), .im_din( 
	_zy_simnet_cceip3_im_din_480_w$[0:95]), .im_vld( 
	_zy_simnet_cceip3_im_vld_481_w$), .im_consumed( 
	_zy_simnet_im_consumed_kme_cceip3_482_w$[0:1]), .im_config( 
	_zy_simnet_cceip3_out_im_config_483_w$[0:11]));
nx_interface_monitor_xcm102 u_nx_interface_monitor_cceip2 ( .stat_code( 
	_zy_simnet_cceip2_out_ia_status_436_w$[0:2]), .stat_datawords( 
	_zy_simnet_cceip2_out_ia_status_437_w$[0:4]), .stat_addr( 
	_zy_simnet_cceip2_out_ia_status_438_w$[0:8]), .capability_lst( 
	_zy_simnet_cceip2_out_ia_capability_439_w$[0:15]), .capability_type( 
	_zy_simnet_cceip2_out_ia_capability_440_w$[0:3]), .rd_dat( 
	_zy_simnet_cceip2_out_ia_rdata_441_w$[0:95]), .bimc_odat( 
	_zy_simnet_cceip3_ism_idat_442_w$), .bimc_osync( 
	_zy_simnet_cceip3_ism_isync_443_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_cceip2_ism_mbe_444_w$), .im_rdy( 
	_zy_simnet_cceip2_im_rdy_445_w$), .im_available( 
	_zy_simnet_im_available_kme_cceip2_446_w$[0:1]), .im_status( 
	_zy_simnet_cceip2_out_im_status_447_w$[0:11]), .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_448_w$[0:10]), .cmnd_op( 
	_zy_simnet_cceip2_out_ia_config_449_w$[0:3]), .cmnd_addr( 
	_zy_simnet_cceip2_out_ia_config_450_w$[0:8]), .wr_stb( 
	_zy_simnet_wr_stb_451_w$), .wr_dat( 
	_zy_simnet_cceip2_out_ia_wdata_452_w$[0:95]), .ovstb( ovstb), .lvm( 
	lvm), .mlvm( mlvm), .mrdten( _zy_simnet_cio_453), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_cceip2_ism_isync_454_w$), 
	.bimc_idat( _zy_simnet_cceip2_ism_idat_455_w$), .im_din( 
	_zy_simnet_cceip2_im_din_456_w$[0:95]), .im_vld( 
	_zy_simnet_cceip2_im_vld_457_w$), .im_consumed( 
	_zy_simnet_im_consumed_kme_cceip2_458_w$[0:1]), .im_config( 
	_zy_simnet_cceip2_out_im_config_459_w$[0:11]));
nx_interface_monitor_xcm103 u_nx_interface_monitor_cceip1 ( .stat_code( 
	_zy_simnet_cceip1_out_ia_status_412_w$[0:2]), .stat_datawords( 
	_zy_simnet_cceip1_out_ia_status_413_w$[0:4]), .stat_addr( 
	_zy_simnet_cceip1_out_ia_status_414_w$[0:8]), .capability_lst( 
	_zy_simnet_cceip1_out_ia_capability_415_w$[0:15]), .capability_type( 
	_zy_simnet_cceip1_out_ia_capability_416_w$[0:3]), .rd_dat( 
	_zy_simnet_cceip1_out_ia_rdata_417_w$[0:95]), .bimc_odat( 
	_zy_simnet_cceip2_ism_idat_418_w$), .bimc_osync( 
	_zy_simnet_cceip2_ism_isync_419_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_cceip1_ism_mbe_420_w$), .im_rdy( 
	_zy_simnet_cceip1_im_rdy_421_w$), .im_available( 
	_zy_simnet_im_available_kme_cceip1_422_w$[0:1]), .im_status( 
	_zy_simnet_cceip1_out_im_status_423_w$[0:11]), .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_424_w$[0:10]), .cmnd_op( 
	_zy_simnet_cceip1_out_ia_config_425_w$[0:3]), .cmnd_addr( 
	_zy_simnet_cceip1_out_ia_config_426_w$[0:8]), .wr_stb( 
	_zy_simnet_wr_stb_427_w$), .wr_dat( 
	_zy_simnet_cceip1_out_ia_wdata_428_w$[0:95]), .ovstb( ovstb), .lvm( 
	lvm), .mlvm( mlvm), .mrdten( _zy_simnet_cio_429), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_cceip1_ism_isync_430_w$), 
	.bimc_idat( _zy_simnet_cceip1_ism_idat_431_w$), .im_din( 
	_zy_simnet_cceip1_im_din_432_w$[0:95]), .im_vld( 
	_zy_simnet_cceip1_im_vld_433_w$), .im_consumed( 
	_zy_simnet_im_consumed_kme_cceip1_434_w$[0:1]), .im_config( 
	_zy_simnet_cceip1_out_im_config_435_w$[0:11]));
nx_interface_monitor_xcm104 u_nx_interface_monitor_cceip0 ( .stat_code( 
	_zy_simnet_cceip0_out_ia_status_388_w$[0:2]), .stat_datawords( 
	_zy_simnet_cceip0_out_ia_status_389_w$[0:4]), .stat_addr( 
	_zy_simnet_cceip0_out_ia_status_390_w$[0:8]), .capability_lst( 
	_zy_simnet_cceip0_out_ia_capability_391_w$[0:15]), .capability_type( 
	_zy_simnet_cceip0_out_ia_capability_392_w$[0:3]), .rd_dat( 
	_zy_simnet_cceip0_out_ia_rdata_393_w$[0:95]), .bimc_odat( 
	_zy_simnet_cceip1_ism_idat_394_w$), .bimc_osync( 
	_zy_simnet_cceip1_ism_isync_395_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_cceip0_ism_mbe_396_w$), .im_rdy( 
	_zy_simnet_cceip0_im_rdy_397_w$), .im_available( 
	_zy_simnet_im_available_kme_cceip0_398_w$[0:1]), .im_status( 
	_zy_simnet_cceip0_out_im_status_399_w$[0:11]), .clk( clk), .rst_n( 
	rst_n), .reg_addr( _zy_simnet_reg_addr_400_w$[0:10]), .cmnd_op( 
	_zy_simnet_cceip0_out_ia_config_401_w$[0:3]), .cmnd_addr( 
	_zy_simnet_cceip0_out_ia_config_402_w$[0:8]), .wr_stb( 
	_zy_simnet_wr_stb_403_w$), .wr_dat( 
	_zy_simnet_cceip0_out_ia_wdata_404_w$[0:95]), .ovstb( ovstb), .lvm( 
	lvm), .mlvm( mlvm), .mrdten( _zy_simnet_cio_405), .bimc_rst_n( 
	bimc_rst_n), .bimc_isync( _zy_simnet_cceip0_ism_bimc_isync_406_w$), 
	.bimc_idat( _zy_simnet_cceip0_ism_bimc_idat_407_w$), .im_din( 
	_zy_simnet_cceip0_im_din_408_w$[0:95]), .im_vld( 
	_zy_simnet_cceip0_im_vld_409_w$), .im_consumed( 
	_zy_simnet_im_consumed_kme_cceip0_410_w$[0:1]), .im_config( 
	_zy_simnet_cceip0_out_im_config_411_w$[0:11]));
nx_interface_monitor_pipe nx_interface_monitor_pipe_cddip3 ( .ob_in_mod( 
	_zy_simnet_kme_cddip3_ob_in_mod_383_w$), .ob_out( 
	_zy_simnet_kme_cddip3_ob_out_post_384_w$[0:82]), .im_vld( 
	_zy_simnet_cddip3_im_vld_385_w$), .clk( clk), .rst_n( rst_n), 
	.ob_out_pre( { kme_cddip3_ob_out_pre[82], kme_cddip3_ob_out_pre[81], 
	cddip3_im_din[14], cddip3_im_din[30], cddip3_im_din[29], 
	cddip3_im_din[28], cddip3_im_din[27], cddip3_im_din[26], 
	cddip3_im_din[25], cddip3_im_din[24], cddip3_im_din[23], 
	cddip3_im_din[13], cddip3_im_din[12], cddip3_im_din[11], 
	cddip3_im_din[10], cddip3_im_din[9], cddip3_im_din[8], 
	kme_cddip3_ob_out_pre[65], cddip3_im_din[6], cddip3_im_din[95], 
	cddip3_im_din[94], cddip3_im_din[93], cddip3_im_din[92], 
	cddip3_im_din[91], cddip3_im_din[90], cddip3_im_din[89], 
	cddip3_im_din[88], cddip3_im_din[87], cddip3_im_din[86], 
	cddip3_im_din[85], cddip3_im_din[84], cddip3_im_din[83], 
	cddip3_im_din[82], cddip3_im_din[81], cddip3_im_din[80], 
	cddip3_im_din[79], cddip3_im_din[78], cddip3_im_din[77], 
	cddip3_im_din[76], cddip3_im_din[75], cddip3_im_din[74], 
	cddip3_im_din[73], cddip3_im_din[72], cddip3_im_din[71], 
	cddip3_im_din[70], cddip3_im_din[69], cddip3_im_din[68], 
	cddip3_im_din[67], cddip3_im_din[66], cddip3_im_din[65], 
	cddip3_im_din[64], cddip3_im_din[63], cddip3_im_din[62], 
	cddip3_im_din[61], cddip3_im_din[60], cddip3_im_din[59], 
	cddip3_im_din[58], cddip3_im_din[57], cddip3_im_din[56], 
	cddip3_im_din[55], cddip3_im_din[54], cddip3_im_din[53], 
	cddip3_im_din[52], cddip3_im_din[51], cddip3_im_din[50], 
	cddip3_im_din[49], cddip3_im_din[48], cddip3_im_din[47], 
	cddip3_im_din[46], cddip3_im_din[45], cddip3_im_din[44], 
	cddip3_im_din[43], cddip3_im_din[42], cddip3_im_din[41], 
	cddip3_im_din[40], cddip3_im_din[39], cddip3_im_din[38], 
	cddip3_im_din[37], cddip3_im_din[36], cddip3_im_din[35], 
	cddip3_im_din[34], cddip3_im_din[33], cddip3_im_din[32]}), .ob_in( 
	_zy_simnet_tvar_386), .im_rdy( _zy_simnet_cddip3_im_rdy_387_w$));
nx_interface_monitor_pipe nx_interface_monitor_pipe_cddip2 ( .ob_in_mod( 
	_zy_simnet_kme_cddip2_ob_in_mod_378_w$), .ob_out( 
	_zy_simnet_kme_cddip2_ob_out_post_379_w$[0:82]), .im_vld( 
	_zy_simnet_cddip2_im_vld_380_w$), .clk( clk), .rst_n( rst_n), 
	.ob_out_pre( { kme_cddip2_ob_out_pre[82], kme_cddip2_ob_out_pre[81], 
	cddip2_im_din[14], cddip2_im_din[30], cddip2_im_din[29], 
	cddip2_im_din[28], cddip2_im_din[27], cddip2_im_din[26], 
	cddip2_im_din[25], cddip2_im_din[24], cddip2_im_din[23], 
	cddip2_im_din[13], cddip2_im_din[12], cddip2_im_din[11], 
	cddip2_im_din[10], cddip2_im_din[9], cddip2_im_din[8], 
	kme_cddip2_ob_out_pre[65], cddip2_im_din[6], cddip2_im_din[95], 
	cddip2_im_din[94], cddip2_im_din[93], cddip2_im_din[92], 
	cddip2_im_din[91], cddip2_im_din[90], cddip2_im_din[89], 
	cddip2_im_din[88], cddip2_im_din[87], cddip2_im_din[86], 
	cddip2_im_din[85], cddip2_im_din[84], cddip2_im_din[83], 
	cddip2_im_din[82], cddip2_im_din[81], cddip2_im_din[80], 
	cddip2_im_din[79], cddip2_im_din[78], cddip2_im_din[77], 
	cddip2_im_din[76], cddip2_im_din[75], cddip2_im_din[74], 
	cddip2_im_din[73], cddip2_im_din[72], cddip2_im_din[71], 
	cddip2_im_din[70], cddip2_im_din[69], cddip2_im_din[68], 
	cddip2_im_din[67], cddip2_im_din[66], cddip2_im_din[65], 
	cddip2_im_din[64], cddip2_im_din[63], cddip2_im_din[62], 
	cddip2_im_din[61], cddip2_im_din[60], cddip2_im_din[59], 
	cddip2_im_din[58], cddip2_im_din[57], cddip2_im_din[56], 
	cddip2_im_din[55], cddip2_im_din[54], cddip2_im_din[53], 
	cddip2_im_din[52], cddip2_im_din[51], cddip2_im_din[50], 
	cddip2_im_din[49], cddip2_im_din[48], cddip2_im_din[47], 
	cddip2_im_din[46], cddip2_im_din[45], cddip2_im_din[44], 
	cddip2_im_din[43], cddip2_im_din[42], cddip2_im_din[41], 
	cddip2_im_din[40], cddip2_im_din[39], cddip2_im_din[38], 
	cddip2_im_din[37], cddip2_im_din[36], cddip2_im_din[35], 
	cddip2_im_din[34], cddip2_im_din[33], cddip2_im_din[32]}), .ob_in( 
	_zy_simnet_tvar_381), .im_rdy( _zy_simnet_cddip2_im_rdy_382_w$));
nx_interface_monitor_pipe nx_interface_monitor_pipe_cddip1 ( .ob_in_mod( 
	_zy_simnet_kme_cddip1_ob_in_mod_373_w$), .ob_out( 
	_zy_simnet_kme_cddip1_ob_out_post_374_w$[0:82]), .im_vld( 
	_zy_simnet_cddip1_im_vld_375_w$), .clk( clk), .rst_n( rst_n), 
	.ob_out_pre( { kme_cddip1_ob_out_pre[82], kme_cddip1_ob_out_pre[81], 
	cddip1_im_din[14], cddip1_im_din[30], cddip1_im_din[29], 
	cddip1_im_din[28], cddip1_im_din[27], cddip1_im_din[26], 
	cddip1_im_din[25], cddip1_im_din[24], cddip1_im_din[23], 
	cddip1_im_din[13], cddip1_im_din[12], cddip1_im_din[11], 
	cddip1_im_din[10], cddip1_im_din[9], cddip1_im_din[8], 
	kme_cddip1_ob_out_pre[65], cddip1_im_din[6], cddip1_im_din[95], 
	cddip1_im_din[94], cddip1_im_din[93], cddip1_im_din[92], 
	cddip1_im_din[91], cddip1_im_din[90], cddip1_im_din[89], 
	cddip1_im_din[88], cddip1_im_din[87], cddip1_im_din[86], 
	cddip1_im_din[85], cddip1_im_din[84], cddip1_im_din[83], 
	cddip1_im_din[82], cddip1_im_din[81], cddip1_im_din[80], 
	cddip1_im_din[79], cddip1_im_din[78], cddip1_im_din[77], 
	cddip1_im_din[76], cddip1_im_din[75], cddip1_im_din[74], 
	cddip1_im_din[73], cddip1_im_din[72], cddip1_im_din[71], 
	cddip1_im_din[70], cddip1_im_din[69], cddip1_im_din[68], 
	cddip1_im_din[67], cddip1_im_din[66], cddip1_im_din[65], 
	cddip1_im_din[64], cddip1_im_din[63], cddip1_im_din[62], 
	cddip1_im_din[61], cddip1_im_din[60], cddip1_im_din[59], 
	cddip1_im_din[58], cddip1_im_din[57], cddip1_im_din[56], 
	cddip1_im_din[55], cddip1_im_din[54], cddip1_im_din[53], 
	cddip1_im_din[52], cddip1_im_din[51], cddip1_im_din[50], 
	cddip1_im_din[49], cddip1_im_din[48], cddip1_im_din[47], 
	cddip1_im_din[46], cddip1_im_din[45], cddip1_im_din[44], 
	cddip1_im_din[43], cddip1_im_din[42], cddip1_im_din[41], 
	cddip1_im_din[40], cddip1_im_din[39], cddip1_im_din[38], 
	cddip1_im_din[37], cddip1_im_din[36], cddip1_im_din[35], 
	cddip1_im_din[34], cddip1_im_din[33], cddip1_im_din[32]}), .ob_in( 
	_zy_simnet_tvar_376), .im_rdy( _zy_simnet_cddip1_im_rdy_377_w$));
nx_interface_monitor_pipe nx_interface_monitor_pipe_cddip0 ( .ob_in_mod( 
	_zy_simnet_kme_cddip0_ob_in_mod_368_w$), .ob_out( 
	_zy_simnet_kme_cddip0_ob_out_post_369_w$[0:82]), .im_vld( 
	_zy_simnet_cddip0_im_vld_370_w$), .clk( clk), .rst_n( rst_n), 
	.ob_out_pre( { kme_cddip0_ob_out_pre[82], kme_cddip0_ob_out_pre[81], 
	cddip0_im_din[14], cddip0_im_din[30], cddip0_im_din[29], 
	cddip0_im_din[28], cddip0_im_din[27], cddip0_im_din[26], 
	cddip0_im_din[25], cddip0_im_din[24], cddip0_im_din[23], 
	cddip0_im_din[13], cddip0_im_din[12], cddip0_im_din[11], 
	cddip0_im_din[10], cddip0_im_din[9], cddip0_im_din[8], 
	kme_cddip0_ob_out_pre[65], cddip0_im_din[6], cddip0_im_din[95], 
	cddip0_im_din[94], cddip0_im_din[93], cddip0_im_din[92], 
	cddip0_im_din[91], cddip0_im_din[90], cddip0_im_din[89], 
	cddip0_im_din[88], cddip0_im_din[87], cddip0_im_din[86], 
	cddip0_im_din[85], cddip0_im_din[84], cddip0_im_din[83], 
	cddip0_im_din[82], cddip0_im_din[81], cddip0_im_din[80], 
	cddip0_im_din[79], cddip0_im_din[78], cddip0_im_din[77], 
	cddip0_im_din[76], cddip0_im_din[75], cddip0_im_din[74], 
	cddip0_im_din[73], cddip0_im_din[72], cddip0_im_din[71], 
	cddip0_im_din[70], cddip0_im_din[69], cddip0_im_din[68], 
	cddip0_im_din[67], cddip0_im_din[66], cddip0_im_din[65], 
	cddip0_im_din[64], cddip0_im_din[63], cddip0_im_din[62], 
	cddip0_im_din[61], cddip0_im_din[60], cddip0_im_din[59], 
	cddip0_im_din[58], cddip0_im_din[57], cddip0_im_din[56], 
	cddip0_im_din[55], cddip0_im_din[54], cddip0_im_din[53], 
	cddip0_im_din[52], cddip0_im_din[51], cddip0_im_din[50], 
	cddip0_im_din[49], cddip0_im_din[48], cddip0_im_din[47], 
	cddip0_im_din[46], cddip0_im_din[45], cddip0_im_din[44], 
	cddip0_im_din[43], cddip0_im_din[42], cddip0_im_din[41], 
	cddip0_im_din[40], cddip0_im_din[39], cddip0_im_din[38], 
	cddip0_im_din[37], cddip0_im_din[36], cddip0_im_din[35], 
	cddip0_im_din[34], cddip0_im_din[33], cddip0_im_din[32]}), .ob_in( 
	_zy_simnet_tvar_371), .im_rdy( _zy_simnet_cddip0_im_rdy_372_w$));
nx_interface_monitor_pipe nx_interface_monitor_pipe_cceip3 ( .ob_in_mod( 
	_zy_simnet_kme_cceip3_ob_in_mod_363_w$), .ob_out( 
	_zy_simnet_kme_cceip3_ob_out_post_364_w$[0:82]), .im_vld( 
	_zy_simnet_cceip3_im_vld_365_w$), .clk( clk), .rst_n( rst_n), 
	.ob_out_pre( { kme_cceip3_ob_out_pre[82], kme_cceip3_ob_out_pre[81], 
	cceip3_im_din[14], cceip3_im_din[30], cceip3_im_din[29], 
	cceip3_im_din[28], cceip3_im_din[27], cceip3_im_din[26], 
	cceip3_im_din[25], cceip3_im_din[24], cceip3_im_din[23], 
	cceip3_im_din[13], cceip3_im_din[12], cceip3_im_din[11], 
	cceip3_im_din[10], cceip3_im_din[9], cceip3_im_din[8], 
	kme_cceip3_ob_out_pre[65], cceip3_im_din[6], cceip3_im_din[95], 
	cceip3_im_din[94], cceip3_im_din[93], cceip3_im_din[92], 
	cceip3_im_din[91], cceip3_im_din[90], cceip3_im_din[89], 
	cceip3_im_din[88], cceip3_im_din[87], cceip3_im_din[86], 
	cceip3_im_din[85], cceip3_im_din[84], cceip3_im_din[83], 
	cceip3_im_din[82], cceip3_im_din[81], cceip3_im_din[80], 
	cceip3_im_din[79], cceip3_im_din[78], cceip3_im_din[77], 
	cceip3_im_din[76], cceip3_im_din[75], cceip3_im_din[74], 
	cceip3_im_din[73], cceip3_im_din[72], cceip3_im_din[71], 
	cceip3_im_din[70], cceip3_im_din[69], cceip3_im_din[68], 
	cceip3_im_din[67], cceip3_im_din[66], cceip3_im_din[65], 
	cceip3_im_din[64], cceip3_im_din[63], cceip3_im_din[62], 
	cceip3_im_din[61], cceip3_im_din[60], cceip3_im_din[59], 
	cceip3_im_din[58], cceip3_im_din[57], cceip3_im_din[56], 
	cceip3_im_din[55], cceip3_im_din[54], cceip3_im_din[53], 
	cceip3_im_din[52], cceip3_im_din[51], cceip3_im_din[50], 
	cceip3_im_din[49], cceip3_im_din[48], cceip3_im_din[47], 
	cceip3_im_din[46], cceip3_im_din[45], cceip3_im_din[44], 
	cceip3_im_din[43], cceip3_im_din[42], cceip3_im_din[41], 
	cceip3_im_din[40], cceip3_im_din[39], cceip3_im_din[38], 
	cceip3_im_din[37], cceip3_im_din[36], cceip3_im_din[35], 
	cceip3_im_din[34], cceip3_im_din[33], cceip3_im_din[32]}), .ob_in( 
	_zy_simnet_tvar_366), .im_rdy( _zy_simnet_cceip3_im_rdy_367_w$));
nx_interface_monitor_pipe nx_interface_monitor_pipe_cceip2 ( .ob_in_mod( 
	_zy_simnet_kme_cceip2_ob_in_mod_358_w$), .ob_out( 
	_zy_simnet_kme_cceip2_ob_out_post_359_w$[0:82]), .im_vld( 
	_zy_simnet_cceip2_im_vld_360_w$), .clk( clk), .rst_n( rst_n), 
	.ob_out_pre( { kme_cceip2_ob_out_pre[82], kme_cceip2_ob_out_pre[81], 
	cceip2_im_din[14], cceip2_im_din[30], cceip2_im_din[29], 
	cceip2_im_din[28], cceip2_im_din[27], cceip2_im_din[26], 
	cceip2_im_din[25], cceip2_im_din[24], cceip2_im_din[23], 
	cceip2_im_din[13], cceip2_im_din[12], cceip2_im_din[11], 
	cceip2_im_din[10], cceip2_im_din[9], cceip2_im_din[8], 
	kme_cceip2_ob_out_pre[65], cceip2_im_din[6], cceip2_im_din[95], 
	cceip2_im_din[94], cceip2_im_din[93], cceip2_im_din[92], 
	cceip2_im_din[91], cceip2_im_din[90], cceip2_im_din[89], 
	cceip2_im_din[88], cceip2_im_din[87], cceip2_im_din[86], 
	cceip2_im_din[85], cceip2_im_din[84], cceip2_im_din[83], 
	cceip2_im_din[82], cceip2_im_din[81], cceip2_im_din[80], 
	cceip2_im_din[79], cceip2_im_din[78], cceip2_im_din[77], 
	cceip2_im_din[76], cceip2_im_din[75], cceip2_im_din[74], 
	cceip2_im_din[73], cceip2_im_din[72], cceip2_im_din[71], 
	cceip2_im_din[70], cceip2_im_din[69], cceip2_im_din[68], 
	cceip2_im_din[67], cceip2_im_din[66], cceip2_im_din[65], 
	cceip2_im_din[64], cceip2_im_din[63], cceip2_im_din[62], 
	cceip2_im_din[61], cceip2_im_din[60], cceip2_im_din[59], 
	cceip2_im_din[58], cceip2_im_din[57], cceip2_im_din[56], 
	cceip2_im_din[55], cceip2_im_din[54], cceip2_im_din[53], 
	cceip2_im_din[52], cceip2_im_din[51], cceip2_im_din[50], 
	cceip2_im_din[49], cceip2_im_din[48], cceip2_im_din[47], 
	cceip2_im_din[46], cceip2_im_din[45], cceip2_im_din[44], 
	cceip2_im_din[43], cceip2_im_din[42], cceip2_im_din[41], 
	cceip2_im_din[40], cceip2_im_din[39], cceip2_im_din[38], 
	cceip2_im_din[37], cceip2_im_din[36], cceip2_im_din[35], 
	cceip2_im_din[34], cceip2_im_din[33], cceip2_im_din[32]}), .ob_in( 
	_zy_simnet_tvar_361), .im_rdy( _zy_simnet_cceip2_im_rdy_362_w$));
nx_interface_monitor_pipe nx_interface_monitor_pipe_cceip1 ( .ob_in_mod( 
	_zy_simnet_kme_cceip1_ob_in_mod_353_w$), .ob_out( 
	_zy_simnet_kme_cceip1_ob_out_post_354_w$[0:82]), .im_vld( 
	_zy_simnet_cceip1_im_vld_355_w$), .clk( clk), .rst_n( rst_n), 
	.ob_out_pre( { kme_cceip1_ob_out_pre[82], kme_cceip1_ob_out_pre[81], 
	cceip1_im_din[14], cceip1_im_din[30], cceip1_im_din[29], 
	cceip1_im_din[28], cceip1_im_din[27], cceip1_im_din[26], 
	cceip1_im_din[25], cceip1_im_din[24], cceip1_im_din[23], 
	cceip1_im_din[13], cceip1_im_din[12], cceip1_im_din[11], 
	cceip1_im_din[10], cceip1_im_din[9], cceip1_im_din[8], 
	kme_cceip1_ob_out_pre[65], cceip1_im_din[6], cceip1_im_din[95], 
	cceip1_im_din[94], cceip1_im_din[93], cceip1_im_din[92], 
	cceip1_im_din[91], cceip1_im_din[90], cceip1_im_din[89], 
	cceip1_im_din[88], cceip1_im_din[87], cceip1_im_din[86], 
	cceip1_im_din[85], cceip1_im_din[84], cceip1_im_din[83], 
	cceip1_im_din[82], cceip1_im_din[81], cceip1_im_din[80], 
	cceip1_im_din[79], cceip1_im_din[78], cceip1_im_din[77], 
	cceip1_im_din[76], cceip1_im_din[75], cceip1_im_din[74], 
	cceip1_im_din[73], cceip1_im_din[72], cceip1_im_din[71], 
	cceip1_im_din[70], cceip1_im_din[69], cceip1_im_din[68], 
	cceip1_im_din[67], cceip1_im_din[66], cceip1_im_din[65], 
	cceip1_im_din[64], cceip1_im_din[63], cceip1_im_din[62], 
	cceip1_im_din[61], cceip1_im_din[60], cceip1_im_din[59], 
	cceip1_im_din[58], cceip1_im_din[57], cceip1_im_din[56], 
	cceip1_im_din[55], cceip1_im_din[54], cceip1_im_din[53], 
	cceip1_im_din[52], cceip1_im_din[51], cceip1_im_din[50], 
	cceip1_im_din[49], cceip1_im_din[48], cceip1_im_din[47], 
	cceip1_im_din[46], cceip1_im_din[45], cceip1_im_din[44], 
	cceip1_im_din[43], cceip1_im_din[42], cceip1_im_din[41], 
	cceip1_im_din[40], cceip1_im_din[39], cceip1_im_din[38], 
	cceip1_im_din[37], cceip1_im_din[36], cceip1_im_din[35], 
	cceip1_im_din[34], cceip1_im_din[33], cceip1_im_din[32]}), .ob_in( 
	_zy_simnet_tvar_356), .im_rdy( _zy_simnet_cceip1_im_rdy_357_w$));
nx_interface_monitor_pipe nx_interface_monitor_pipe_cceip0 ( .ob_in_mod( 
	_zy_simnet_kme_cceip0_ob_in_mod_348_w$), .ob_out( 
	_zy_simnet_kme_cceip0_ob_out_post_349_w$[0:82]), .im_vld( 
	_zy_simnet_cceip0_im_vld_350_w$), .clk( clk), .rst_n( rst_n), 
	.ob_out_pre( { kme_cceip0_ob_out_pre[82], kme_cceip0_ob_out_pre[81], 
	cceip0_im_din[14], cceip0_im_din[30], cceip0_im_din[29], 
	cceip0_im_din[28], cceip0_im_din[27], cceip0_im_din[26], 
	cceip0_im_din[25], cceip0_im_din[24], cceip0_im_din[23], 
	cceip0_im_din[13], cceip0_im_din[12], cceip0_im_din[11], 
	cceip0_im_din[10], cceip0_im_din[9], cceip0_im_din[8], 
	kme_cceip0_ob_out_pre[65], cceip0_im_din[6], cceip0_im_din[95], 
	cceip0_im_din[94], cceip0_im_din[93], cceip0_im_din[92], 
	cceip0_im_din[91], cceip0_im_din[90], cceip0_im_din[89], 
	cceip0_im_din[88], cceip0_im_din[87], cceip0_im_din[86], 
	cceip0_im_din[85], cceip0_im_din[84], cceip0_im_din[83], 
	cceip0_im_din[82], cceip0_im_din[81], cceip0_im_din[80], 
	cceip0_im_din[79], cceip0_im_din[78], cceip0_im_din[77], 
	cceip0_im_din[76], cceip0_im_din[75], cceip0_im_din[74], 
	cceip0_im_din[73], cceip0_im_din[72], cceip0_im_din[71], 
	cceip0_im_din[70], cceip0_im_din[69], cceip0_im_din[68], 
	cceip0_im_din[67], cceip0_im_din[66], cceip0_im_din[65], 
	cceip0_im_din[64], cceip0_im_din[63], cceip0_im_din[62], 
	cceip0_im_din[61], cceip0_im_din[60], cceip0_im_din[59], 
	cceip0_im_din[58], cceip0_im_din[57], cceip0_im_din[56], 
	cceip0_im_din[55], cceip0_im_din[54], cceip0_im_din[53], 
	cceip0_im_din[52], cceip0_im_din[51], cceip0_im_din[50], 
	cceip0_im_din[49], cceip0_im_din[48], cceip0_im_din[47], 
	cceip0_im_din[46], cceip0_im_din[45], cceip0_im_din[44], 
	cceip0_im_din[43], cceip0_im_din[42], cceip0_im_din[41], 
	cceip0_im_din[40], cceip0_im_din[39], cceip0_im_din[38], 
	cceip0_im_din[37], cceip0_im_din[36], cceip0_im_din[35], 
	cceip0_im_din[34], cceip0_im_din[33], cceip0_im_din[32]}), .ob_in( 
	_zy_simnet_tvar_351), .im_rdy( _zy_simnet_cceip0_im_rdy_352_w$));
nx_rbus_ring u_nx_rbus_ring ( .clk( clk), .rst_n( rst_n), .cfg_start_addr( 
	cfg_start_addr[15:0]), .cfg_end_addr( cfg_end_addr[15:0]), 
	.rbus_addr_i( rbus_ring_i[83:68]), .rbus_wr_strb_i( 
	rbus_ring_i[67]), .rbus_wr_data_i( rbus_ring_i[66:35]), 
	.rbus_rd_strb_i( rbus_ring_i[34]), .rbus_addr_o( 
	_zy_simnet_rbus_ring_o_334_w$[0:15]), .rbus_wr_strb_o( 
	_zy_simnet_rbus_ring_o_335_w$), .rbus_wr_data_o( 
	_zy_simnet_rbus_ring_o_336_w$[0:31]), .rbus_rd_strb_o( 
	_zy_simnet_rbus_ring_o_337_w$), .locl_addr_o( 
	_zy_simnet_locl_addr_338_w$[0:10]), .locl_wr_strb_o( 
	_zy_simnet_locl_wr_strb_339_w$), .locl_wr_data_o( 
	_zy_simnet_locl_wr_data_340_w$[0:31]), .locl_rd_strb_o( 
	_zy_simnet_locl_rd_strb_341_w$), .rbus_rd_data_i( 
	rbus_ring_i[33:2]), .rbus_ack_i( rbus_ring_i[1]), .rbus_err_ack_i( 
	rbus_ring_i[0]), .locl_rd_data_i( 
	_zy_simnet_locl_rd_data_342_w$[0:31]), .locl_ack_i( 
	_zy_simnet_locl_ack_343_w$), .locl_err_ack_i( 
	_zy_simnet_locl_err_ack_344_w$), .rbus_rd_data_o( 
	_zy_simnet_rbus_ring_o_345_w$[0:31]), .rbus_ack_o( 
	_zy_simnet_rbus_ring_o_346_w$), .rbus_err_ack_o( 
	_zy_simnet_rbus_ring_o_347_w$));
cr_kme_regs u_cr_kme_regs ( .clk( clk), .i_reset_( rst_n), .i_sw_init( 
	_zy_simnet_cio_24), .i_addr( _zy_simnet_locl_addr_25_w$[0:10]), 
	.i_wr_strb( _zy_simnet_locl_wr_strb_26_w$), .i_wr_data( 
	_zy_simnet_locl_wr_data_27_w$[0:31]), .i_rd_strb( 
	_zy_simnet_locl_rd_strb_28_w$), .o_rd_data( 
	_zy_simnet_locl_rd_data_29_w$[0:31]), .o_ack( 
	_zy_simnet_locl_ack_30_w$), .o_err_ack( 
	_zy_simnet_locl_err_ack_31_w$), .o_spare_config( 
	_zy_simnet_tvar_32[0:31]), .o_cceip0_out_ia_wdata_part0( 
	_zy_simnet_cceip0_out_ia_wdata_38_w$[0:31]), 
	.o_cceip0_out_ia_wdata_part1( 
	_zy_simnet_cceip0_out_ia_wdata_39_w$[0:31]), 
	.o_cceip0_out_ia_wdata_part2( 
	_zy_simnet_cceip0_out_ia_wdata_40_w$[0:31]), .o_cceip0_out_ia_config( 
	_zy_simnet_cceip0_out_ia_config_41_w$[0:12]), .o_cceip0_out_im_config( 
	_zy_simnet_cceip0_out_im_config_42_w$[0:11]), 
	.o_cceip0_out_im_read_done( _zy_simnet_dio_43[0:1]), 
	.o_cceip1_out_ia_wdata_part0( 
	_zy_simnet_cceip1_out_ia_wdata_44_w$[0:31]), 
	.o_cceip1_out_ia_wdata_part1( 
	_zy_simnet_cceip1_out_ia_wdata_45_w$[0:31]), 
	.o_cceip1_out_ia_wdata_part2( 
	_zy_simnet_cceip1_out_ia_wdata_46_w$[0:31]), .o_cceip1_out_ia_config( 
	_zy_simnet_cceip1_out_ia_config_47_w$[0:12]), .o_cceip1_out_im_config( 
	_zy_simnet_cceip1_out_im_config_48_w$[0:11]), 
	.o_cceip1_out_im_read_done( _zy_simnet_dio_49[0:1]), 
	.o_cceip2_out_ia_wdata_part0( 
	_zy_simnet_cceip2_out_ia_wdata_50_w$[0:31]), 
	.o_cceip2_out_ia_wdata_part1( 
	_zy_simnet_cceip2_out_ia_wdata_51_w$[0:31]), 
	.o_cceip2_out_ia_wdata_part2( 
	_zy_simnet_cceip2_out_ia_wdata_52_w$[0:31]), .o_cceip2_out_ia_config( 
	_zy_simnet_cceip2_out_ia_config_53_w$[0:12]), .o_cceip2_out_im_config( 
	_zy_simnet_cceip2_out_im_config_54_w$[0:11]), 
	.o_cceip2_out_im_read_done( _zy_simnet_dio_55[0:1]), 
	.o_cceip3_out_ia_wdata_part0( 
	_zy_simnet_cceip3_out_ia_wdata_56_w$[0:31]), 
	.o_cceip3_out_ia_wdata_part1( 
	_zy_simnet_cceip3_out_ia_wdata_57_w$[0:31]), 
	.o_cceip3_out_ia_wdata_part2( 
	_zy_simnet_cceip3_out_ia_wdata_58_w$[0:31]), .o_cceip3_out_ia_config( 
	_zy_simnet_cceip3_out_ia_config_59_w$[0:12]), .o_cceip3_out_im_config( 
	_zy_simnet_cceip3_out_im_config_60_w$[0:11]), 
	.o_cceip3_out_im_read_done( _zy_simnet_dio_61[0:1]), 
	.o_cddip0_out_ia_wdata_part0( 
	_zy_simnet_cddip0_out_ia_wdata_62_w$[0:31]), 
	.o_cddip0_out_ia_wdata_part1( 
	_zy_simnet_cddip0_out_ia_wdata_63_w$[0:31]), 
	.o_cddip0_out_ia_wdata_part2( 
	_zy_simnet_cddip0_out_ia_wdata_64_w$[0:31]), .o_cddip0_out_ia_config( 
	_zy_simnet_cddip0_out_ia_config_65_w$[0:12]), .o_cddip0_out_im_config( 
	_zy_simnet_cddip0_out_im_config_66_w$[0:11]), 
	.o_cddip0_out_im_read_done( _zy_simnet_dio_67[0:1]), 
	.o_cddip1_out_ia_wdata_part0( 
	_zy_simnet_cddip1_out_ia_wdata_68_w$[0:31]), 
	.o_cddip1_out_ia_wdata_part1( 
	_zy_simnet_cddip1_out_ia_wdata_69_w$[0:31]), 
	.o_cddip1_out_ia_wdata_part2( 
	_zy_simnet_cddip1_out_ia_wdata_70_w$[0:31]), .o_cddip1_out_ia_config( 
	_zy_simnet_cddip1_out_ia_config_71_w$[0:12]), .o_cddip1_out_im_config( 
	_zy_simnet_cddip1_out_im_config_72_w$[0:11]), 
	.o_cddip1_out_im_read_done( _zy_simnet_dio_73[0:1]), 
	.o_cddip2_out_ia_wdata_part0( 
	_zy_simnet_cddip2_out_ia_wdata_74_w$[0:31]), 
	.o_cddip2_out_ia_wdata_part1( 
	_zy_simnet_cddip2_out_ia_wdata_75_w$[0:31]), 
	.o_cddip2_out_ia_wdata_part2( 
	_zy_simnet_cddip2_out_ia_wdata_76_w$[0:31]), .o_cddip2_out_ia_config( 
	_zy_simnet_cddip2_out_ia_config_77_w$[0:12]), .o_cddip2_out_im_config( 
	_zy_simnet_cddip2_out_im_config_78_w$[0:11]), 
	.o_cddip2_out_im_read_done( _zy_simnet_dio_79[0:1]), 
	.o_cddip3_out_ia_wdata_part0( 
	_zy_simnet_cddip3_out_ia_wdata_80_w$[0:31]), 
	.o_cddip3_out_ia_wdata_part1( 
	_zy_simnet_cddip3_out_ia_wdata_81_w$[0:31]), 
	.o_cddip3_out_ia_wdata_part2( 
	_zy_simnet_cddip3_out_ia_wdata_82_w$[0:31]), .o_cddip3_out_ia_config( 
	_zy_simnet_cddip3_out_ia_config_83_w$[0:12]), .o_cddip3_out_im_config( 
	_zy_simnet_cddip3_out_im_config_84_w$[0:11]), 
	.o_cddip3_out_im_read_done( _zy_simnet_dio_85[0:1]), 
	.o_ckv_ia_wdata_part0( _zy_simnet_o_ckv_ia_wdata_part0_86_w$[0:31]), 
	.o_ckv_ia_wdata_part1( _zy_simnet_o_ckv_ia_wdata_part1_87_w$[0:31]), 
	.o_ckv_ia_config( _zy_simnet_o_ckv_ia_config_88_w$[0:18]), 
	.o_kim_ia_wdata_part0( _zy_simnet_o_kim_ia_wdata_part0_89_w$[0:20]), 
	.o_kim_ia_wdata_part1( _zy_simnet_o_kim_ia_wdata_part1_90_w$[0:16]), 
	.o_kim_ia_config( _zy_simnet_o_kim_ia_config_91_w$[0:17]), 
	.o_label0_config( _zy_simnet_tvar_92[0:15]), .o_label0_data7( 
	_zy_simnet_labels_93_w$[0:31]), .o_label0_data6( 
	_zy_simnet_labels_94_w$[0:31]), .o_label0_data5( 
	_zy_simnet_labels_95_w$[0:31]), .o_label0_data4( 
	_zy_simnet_labels_96_w$[0:31]), .o_label0_data3( 
	_zy_simnet_labels_97_w$[0:31]), .o_label0_data2( 
	_zy_simnet_labels_98_w$[0:31]), .o_label0_data1( 
	_zy_simnet_labels_99_w$[0:31]), .o_label0_data0( 
	_zy_simnet_labels_100_w$[0:31]), .o_label1_config( 
	_zy_simnet_tvar_101[0:15]), .o_label1_data7( 
	_zy_simnet_labels_102_w$[0:31]), .o_label1_data6( 
	_zy_simnet_labels_103_w$[0:31]), .o_label1_data5( 
	_zy_simnet_labels_104_w$[0:31]), .o_label1_data4( 
	_zy_simnet_labels_105_w$[0:31]), .o_label1_data3( 
	_zy_simnet_labels_106_w$[0:31]), .o_label1_data2( 
	_zy_simnet_labels_107_w$[0:31]), .o_label1_data1( 
	_zy_simnet_labels_108_w$[0:31]), .o_label1_data0( 
	_zy_simnet_labels_109_w$[0:31]), .o_label2_config( 
	_zy_simnet_tvar_110[0:15]), .o_label2_data7( 
	_zy_simnet_labels_111_w$[0:31]), .o_label2_data6( 
	_zy_simnet_labels_112_w$[0:31]), .o_label2_data5( 
	_zy_simnet_labels_113_w$[0:31]), .o_label2_data4( 
	_zy_simnet_labels_114_w$[0:31]), .o_label2_data3( 
	_zy_simnet_labels_115_w$[0:31]), .o_label2_data2( 
	_zy_simnet_labels_116_w$[0:31]), .o_label2_data1( 
	_zy_simnet_labels_117_w$[0:31]), .o_label2_data0( 
	_zy_simnet_labels_118_w$[0:31]), .o_label3_config( 
	_zy_simnet_tvar_119[0:15]), .o_label3_data7( 
	_zy_simnet_labels_120_w$[0:31]), .o_label3_data6( 
	_zy_simnet_labels_121_w$[0:31]), .o_label3_data5( 
	_zy_simnet_labels_122_w$[0:31]), .o_label3_data4( 
	_zy_simnet_labels_123_w$[0:31]), .o_label3_data3( 
	_zy_simnet_labels_124_w$[0:31]), .o_label3_data2( 
	_zy_simnet_labels_125_w$[0:31]), .o_label3_data1( 
	_zy_simnet_labels_126_w$[0:31]), .o_label3_data0( 
	_zy_simnet_labels_127_w$[0:31]), .o_label4_config( 
	_zy_simnet_tvar_128[0:15]), .o_label4_data7( 
	_zy_simnet_labels_129_w$[0:31]), .o_label4_data6( 
	_zy_simnet_labels_130_w$[0:31]), .o_label4_data5( 
	_zy_simnet_labels_131_w$[0:31]), .o_label4_data4( 
	_zy_simnet_labels_132_w$[0:31]), .o_label4_data3( 
	_zy_simnet_labels_133_w$[0:31]), .o_label4_data2( 
	_zy_simnet_labels_134_w$[0:31]), .o_label4_data1( 
	_zy_simnet_labels_135_w$[0:31]), .o_label4_data0( 
	_zy_simnet_labels_136_w$[0:31]), .o_label5_config( 
	_zy_simnet_tvar_137[0:15]), .o_label5_data7( 
	_zy_simnet_labels_138_w$[0:31]), .o_label5_data6( 
	_zy_simnet_labels_139_w$[0:31]), .o_label5_data5( 
	_zy_simnet_labels_140_w$[0:31]), .o_label5_data4( 
	_zy_simnet_labels_141_w$[0:31]), .o_label5_data3( 
	_zy_simnet_labels_142_w$[0:31]), .o_label5_data2( 
	_zy_simnet_labels_143_w$[0:31]), .o_label5_data1( 
	_zy_simnet_labels_144_w$[0:31]), .o_label5_data0( 
	_zy_simnet_labels_145_w$[0:31]), .o_label6_config( 
	_zy_simnet_tvar_146[0:15]), .o_label6_data7( 
	_zy_simnet_labels_147_w$[0:31]), .o_label6_data6( 
	_zy_simnet_labels_148_w$[0:31]), .o_label6_data5( 
	_zy_simnet_labels_149_w$[0:31]), .o_label6_data4( 
	_zy_simnet_labels_150_w$[0:31]), .o_label6_data3( 
	_zy_simnet_labels_151_w$[0:31]), .o_label6_data2( 
	_zy_simnet_labels_152_w$[0:31]), .o_label6_data1( 
	_zy_simnet_labels_153_w$[0:31]), .o_label6_data0( 
	_zy_simnet_labels_154_w$[0:31]), .o_label7_config( 
	_zy_simnet_tvar_155[0:15]), .o_label7_data7( 
	_zy_simnet_labels_156_w$[0:31]), .o_label7_data6( 
	_zy_simnet_labels_157_w$[0:31]), .o_label7_data5( 
	_zy_simnet_labels_158_w$[0:31]), .o_label7_data4( 
	_zy_simnet_labels_159_w$[0:31]), .o_label7_data3( 
	_zy_simnet_labels_160_w$[0:31]), .o_label7_data2( 
	_zy_simnet_labels_161_w$[0:31]), .o_label7_data1( 
	_zy_simnet_labels_162_w$[0:31]), .o_label7_data0( 
	_zy_simnet_labels_163_w$[0:31]), .o_kdf_drbg_ctrl( 
	_zy_simnet_o_kdf_drbg_ctrl_164_w$[0:1]), 
	.o_kdf_drbg_seed_0_state_key_31_0( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_31_0_165_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_63_32( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_63_32_166_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_95_64( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_95_64_167_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_127_96( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_127_96_168_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_159_128( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_159_128_169_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_191_160( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_191_160_170_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_223_192( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_223_192_171_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_key_255_224( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_255_224_172_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_value_31_0( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_31_0_173_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_value_63_32( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_63_32_174_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_value_95_64( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_95_64_175_w$[0:31]), 
	.o_kdf_drbg_seed_0_state_value_127_96( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_127_96_176_w$[0:31]), 
	.o_kdf_drbg_seed_0_reseed_interval_0( 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_0_177_w$[0:31]), 
	.o_kdf_drbg_seed_0_reseed_interval_1( 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_1_178_w$[0:15]), 
	.o_kdf_drbg_seed_1_state_key_31_0( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_31_0_179_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_63_32( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_63_32_180_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_95_64( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_95_64_181_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_127_96( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_127_96_182_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_159_128( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_159_128_183_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_191_160( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_191_160_184_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_223_192( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_223_192_185_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_key_255_224( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_255_224_186_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_value_31_0( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_31_0_187_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_value_63_32( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_63_32_188_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_value_95_64( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_95_64_189_w$[0:31]), 
	.o_kdf_drbg_seed_1_state_value_127_96( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_127_96_190_w$[0:31]), 
	.o_kdf_drbg_seed_1_reseed_interval_0( 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_0_191_w$[0:31]), 
	.o_kdf_drbg_seed_1_reseed_interval_1( 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_1_192_w$[0:15]), 
	.o_interrupt_status( _zy_simnet_dio_193[0:4]), .o_interrupt_mask( 
	_zy_simnet_o_interrupt_mask_194_w$[0:4]), .o_engine_sticky_status( 
	_zy_simnet_o_engine_sticky_status_195_w$[0:7]), .o_bimc_monitor_mask( 
	_zy_simnet_o_bimc_monitor_mask_196_w$[0:6]), 
	.o_bimc_ecc_uncorrectable_error_cnt( 
	_zy_simnet_o_bimc_ecc_uncorrectable_error_cnt_197_w$[0:31]), 
	.o_bimc_ecc_correctable_error_cnt( 
	_zy_simnet_o_bimc_ecc_correctable_error_cnt_198_w$[0:31]), 
	.o_bimc_parity_error_cnt( 
	_zy_simnet_o_bimc_parity_error_cnt_199_w$[0:31]), 
	.o_bimc_global_config( _zy_simnet_o_bimc_global_config_200_w$[0:31]), 
	.o_bimc_eccpar_debug( _zy_simnet_o_bimc_eccpar_debug_201_w$[0:28]), 
	.o_bimc_cmd2( _zy_simnet_o_bimc_cmd2_202_w$[0:10]), .o_bimc_cmd1( 
	_zy_simnet_o_bimc_cmd1_203_w$[0:31]), .o_bimc_cmd0( 
	_zy_simnet_o_bimc_cmd0_204_w$[0:31]), .o_bimc_rxcmd2( 
	_zy_simnet_o_bimc_rxcmd2_205_w$[0:9]), .o_bimc_rxrsp2( 
	_zy_simnet_o_bimc_rxrsp2_206_w$[0:9]), .o_bimc_pollrsp2( 
	_zy_simnet_o_bimc_pollrsp2_207_w$[0:9]), .o_bimc_dbgcmd2( 
	_zy_simnet_o_bimc_dbgcmd2_208_w$[0:9]), .o_im_consumed( 
	_zy_simnet_dio_209[0:15]), .o_tready_override( 
	_zy_simnet_tready_override_210_w$[0:8]), .o_regs_sa_ctrl( 
	_zy_simnet_regs_sa_ctrl_211_w$[0:31]), .o_sa_snapshot_ia_wdata_part0( 
	_zy_simnet_sa_snapshot_ia_wdata_212_w$[0:31]), 
	.o_sa_snapshot_ia_wdata_part1( 
	_zy_simnet_sa_snapshot_ia_wdata_213_w$[0:31]), 
	.o_sa_snapshot_ia_config( 
	_zy_simnet_sa_snapshot_ia_config_214_w$[0:8]), 
	.o_sa_count_ia_wdata_part0( 
	_zy_simnet_sa_count_ia_wdata_215_w$[0:31]), .o_sa_count_ia_wdata_part1( 
	_zy_simnet_sa_count_ia_wdata_216_w$[0:31]), .o_sa_count_ia_config( 
	_zy_simnet_sa_count_ia_config_217_w$[0:8]), 
	.o_cceip_encrypt_kop_fifo_override( 
	_zy_simnet_cceip_encrypt_kop_fifo_override_218_w$[0:6]), 
	.o_cceip_validate_kop_fifo_override( 
	_zy_simnet_cceip_validate_kop_fifo_override_219_w$[0:6]), 
	.o_cddip_decrypt_kop_fifo_override( 
	_zy_simnet_cddip_decrypt_kop_fifo_override_220_w$[0:6]), 
	.o_sa_global_ctrl( _zy_simnet_sa_global_ctrl_221_w$[0:31]), 
	.o_sa_ctrl_ia_wdata_part0( _zy_simnet_sa_ctrl_ia_wdata_222_w$[0:31]), 
	.o_sa_ctrl_ia_config( _zy_simnet_sa_ctrl_ia_config_223_w$[0:8]), 
	.o_kdf_test_key_size_config( kdf_test_key_size[31:0]), 
	.i_blkid_revid_config( _zy_simnet_blkid_revid_config_224_w$[0:31]), 
	.i_revision_config( _zy_simnet_revid_wire_225_w$[0:7]), 
	.i_spare_config( _zy_simnet_tvar_226[0:31]), 
	.i_cceip0_out_ia_capability( 
	_zy_simnet_cceip0_out_ia_capability_227_w$[0:19]), 
	.i_cceip0_out_ia_status( 
	_zy_simnet_cceip0_out_ia_status_228_w$[0:16]), 
	.i_cceip0_out_ia_rdata_part0( _zy_simnet_tvar_229[0:31]), 
	.i_cceip0_out_ia_rdata_part1( _zy_simnet_tvar_230[0:31]), 
	.i_cceip0_out_ia_rdata_part2( _zy_simnet_tvar_231[0:31]), 
	.i_cceip0_out_im_status( 
	_zy_simnet_cceip0_out_im_status_232_w$[0:11]), 
	.i_cceip0_out_im_read_done( _zy_simnet_cio_233[0:1]), 
	.i_cceip1_out_ia_capability( 
	_zy_simnet_cceip1_out_ia_capability_234_w$[0:19]), 
	.i_cceip1_out_ia_status( 
	_zy_simnet_cceip1_out_ia_status_235_w$[0:16]), 
	.i_cceip1_out_ia_rdata_part0( _zy_simnet_tvar_236[0:31]), 
	.i_cceip1_out_ia_rdata_part1( _zy_simnet_tvar_237[0:31]), 
	.i_cceip1_out_ia_rdata_part2( _zy_simnet_tvar_238[0:31]), 
	.i_cceip1_out_im_status( 
	_zy_simnet_cceip1_out_im_status_239_w$[0:11]), 
	.i_cceip1_out_im_read_done( _zy_simnet_cio_240[0:1]), 
	.i_cceip2_out_ia_capability( 
	_zy_simnet_cceip2_out_ia_capability_241_w$[0:19]), 
	.i_cceip2_out_ia_status( 
	_zy_simnet_cceip2_out_ia_status_242_w$[0:16]), 
	.i_cceip2_out_ia_rdata_part0( _zy_simnet_tvar_243[0:31]), 
	.i_cceip2_out_ia_rdata_part1( _zy_simnet_tvar_244[0:31]), 
	.i_cceip2_out_ia_rdata_part2( _zy_simnet_tvar_245[0:31]), 
	.i_cceip2_out_im_status( 
	_zy_simnet_cceip2_out_im_status_246_w$[0:11]), 
	.i_cceip2_out_im_read_done( _zy_simnet_cio_247[0:1]), 
	.i_cceip3_out_ia_capability( 
	_zy_simnet_cceip3_out_ia_capability_248_w$[0:19]), 
	.i_cceip3_out_ia_status( 
	_zy_simnet_cceip3_out_ia_status_249_w$[0:16]), 
	.i_cceip3_out_ia_rdata_part0( _zy_simnet_tvar_250[0:31]), 
	.i_cceip3_out_ia_rdata_part1( _zy_simnet_tvar_251[0:31]), 
	.i_cceip3_out_ia_rdata_part2( _zy_simnet_tvar_252[0:31]), 
	.i_cceip3_out_im_status( 
	_zy_simnet_cceip3_out_im_status_253_w$[0:11]), 
	.i_cceip3_out_im_read_done( _zy_simnet_cio_254[0:1]), 
	.i_cddip0_out_ia_capability( 
	_zy_simnet_cddip0_out_ia_capability_255_w$[0:19]), 
	.i_cddip0_out_ia_status( 
	_zy_simnet_cddip0_out_ia_status_256_w$[0:16]), 
	.i_cddip0_out_ia_rdata_part0( _zy_simnet_tvar_257[0:31]), 
	.i_cddip0_out_ia_rdata_part1( _zy_simnet_tvar_258[0:31]), 
	.i_cddip0_out_ia_rdata_part2( _zy_simnet_tvar_259[0:31]), 
	.i_cddip0_out_im_status( 
	_zy_simnet_cddip0_out_im_status_260_w$[0:11]), 
	.i_cddip0_out_im_read_done( _zy_simnet_cio_261[0:1]), 
	.i_cddip1_out_ia_capability( 
	_zy_simnet_cddip1_out_ia_capability_262_w$[0:19]), 
	.i_cddip1_out_ia_status( 
	_zy_simnet_cddip1_out_ia_status_263_w$[0:16]), 
	.i_cddip1_out_ia_rdata_part0( _zy_simnet_tvar_264[0:31]), 
	.i_cddip1_out_ia_rdata_part1( _zy_simnet_tvar_265[0:31]), 
	.i_cddip1_out_ia_rdata_part2( _zy_simnet_tvar_266[0:31]), 
	.i_cddip1_out_im_status( 
	_zy_simnet_cddip1_out_im_status_267_w$[0:11]), 
	.i_cddip1_out_im_read_done( _zy_simnet_cio_268[0:1]), 
	.i_cddip2_out_ia_capability( 
	_zy_simnet_cddip2_out_ia_capability_269_w$[0:19]), 
	.i_cddip2_out_ia_status( 
	_zy_simnet_cddip2_out_ia_status_270_w$[0:16]), 
	.i_cddip2_out_ia_rdata_part0( _zy_simnet_tvar_271[0:31]), 
	.i_cddip2_out_ia_rdata_part1( _zy_simnet_tvar_272[0:31]), 
	.i_cddip2_out_ia_rdata_part2( _zy_simnet_tvar_273[0:31]), 
	.i_cddip2_out_im_status( 
	_zy_simnet_cddip2_out_im_status_274_w$[0:11]), 
	.i_cddip2_out_im_read_done( _zy_simnet_cio_275[0:1]), 
	.i_cddip3_out_ia_capability( 
	_zy_simnet_cddip3_out_ia_capability_276_w$[0:19]), 
	.i_cddip3_out_ia_status( 
	_zy_simnet_cddip3_out_ia_status_277_w$[0:16]), 
	.i_cddip3_out_ia_rdata_part0( _zy_simnet_tvar_278[0:31]), 
	.i_cddip3_out_ia_rdata_part1( _zy_simnet_tvar_279[0:31]), 
	.i_cddip3_out_ia_rdata_part2( _zy_simnet_tvar_280[0:31]), 
	.i_cddip3_out_im_status( 
	_zy_simnet_cddip3_out_im_status_281_w$[0:11]), 
	.i_cddip3_out_im_read_done( _zy_simnet_cio_282[0:1]), 
	.i_ckv_ia_capability( _zy_simnet_ckv_ia_capability_283_w$[0:19]), 
	.i_ckv_ia_status( _zy_simnet_ckv_ia_status_284_w$[0:22]), 
	.i_ckv_ia_rdata_part0( _zy_simnet_ckv_ia_rdata_part0_285_w$[0:31]), 
	.i_ckv_ia_rdata_part1( _zy_simnet_ckv_ia_rdata_part1_286_w$[0:31]), 
	.i_kim_ia_capability( _zy_simnet_kim_ia_capability_287_w$[0:19]), 
	.i_kim_ia_status( _zy_simnet_kim_ia_status_288_w$[0:21]), 
	.i_kim_ia_rdata_part0( _zy_simnet_kim_ia_rdata_part0_289_w$[0:20]), 
	.i_kim_ia_rdata_part1( _zy_simnet_kim_ia_rdata_part1_290_w$[0:16]), 
	.i_kdf_drbg_ctrl( _zy_simnet_kdf_drbg_ctrl_291_w$[0:1]), 
	.i_interrupt_status( _zy_simnet_interrupt_status_292_w$[0:4]), 
	.i_engine_sticky_status( 
	_zy_simnet_engine_sticky_status_293_w$[0:7]), .i_bimc_monitor( 
	_zy_simnet_bimc_monitor_294_w$[0:6]), 
	.i_bimc_ecc_uncorrectable_error_cnt( 
	_zy_simnet_bimc_ecc_uncorrectable_error_cnt_295_w$[0:31]), 
	.i_bimc_ecc_correctable_error_cnt( 
	_zy_simnet_bimc_ecc_correctable_error_cnt_296_w$[0:31]), 
	.i_bimc_parity_error_cnt( 
	_zy_simnet_bimc_parity_error_cnt_297_w$[0:31]), .i_bimc_global_config( 
	_zy_simnet_bimc_global_config_298_w$[0:31]), .i_bimc_memid( 
	_zy_simnet_bimc_memid_299_w$[0:11]), .i_bimc_eccpar_debug( 
	_zy_simnet_bimc_eccpar_debug_300_w$[0:28]), .i_bimc_cmd2( 
	_zy_simnet_bimc_cmd2_301_w$[0:10]), .i_bimc_rxcmd2( 
	_zy_simnet_bimc_rxcmd2_302_w$[0:9]), .i_bimc_rxcmd1( 
	_zy_simnet_bimc_rxcmd1_303_w$[0:31]), .i_bimc_rxcmd0( 
	_zy_simnet_bimc_rxcmd0_304_w$[0:31]), .i_bimc_rxrsp2( 
	_zy_simnet_bimc_rxrsp2_305_w$[0:9]), .i_bimc_rxrsp1( 
	_zy_simnet_bimc_rxrsp1_306_w$[0:31]), .i_bimc_rxrsp0( 
	_zy_simnet_bimc_rxrsp0_307_w$[0:31]), .i_bimc_pollrsp2( 
	_zy_simnet_bimc_pollrsp2_308_w$[0:9]), .i_bimc_pollrsp1( 
	_zy_simnet_bimc_pollrsp1_309_w$[0:31]), .i_bimc_pollrsp0( 
	_zy_simnet_bimc_pollrsp0_310_w$[0:31]), .i_bimc_dbgcmd2( 
	_zy_simnet_bimc_dbgcmd2_311_w$[0:9]), .i_bimc_dbgcmd1( 
	_zy_simnet_bimc_dbgcmd1_312_w$[0:31]), .i_bimc_dbgcmd0( 
	_zy_simnet_bimc_dbgcmd0_313_w$[0:31]), .i_im_available( 
	_zy_simnet_im_available_314_w$[0:15]), .i_im_consumed( 
	_zy_simnet_cio_315[0:15]), .i_tready_override( 
	_zy_simnet_tready_override_316_w$[0:8]), .i_regs_sa_ctrl( 
	_zy_simnet_regs_sa_ctrl_317_w$[0:31]), .i_sa_snapshot_ia_capability( 
	_zy_simnet_sa_snapshot_ia_capability_318_w$[0:19]), 
	.i_sa_snapshot_ia_status( 
	_zy_simnet_sa_snapshot_ia_status_319_w$[0:12]), 
	.i_sa_snapshot_ia_rdata_part0( 
	_zy_simnet_sa_snapshot_ia_rdata_320_w$[0:31]), 
	.i_sa_snapshot_ia_rdata_part1( 
	_zy_simnet_sa_snapshot_ia_rdata_321_w$[0:31]), 
	.i_sa_count_ia_capability( 
	_zy_simnet_sa_count_ia_capability_322_w$[0:19]), .i_sa_count_ia_status( 
	_zy_simnet_sa_count_ia_status_323_w$[0:12]), 
	.i_sa_count_ia_rdata_part0( 
	_zy_simnet_sa_count_ia_rdata_324_w$[0:31]), .i_sa_count_ia_rdata_part1( 
	_zy_simnet_sa_count_ia_rdata_325_w$[0:31]), .i_idle_components( 
	idle_components[31:0]), .i_sa_global_ctrl( 
	_zy_simnet_sa_global_ctrl_326_w$[0:31]), .i_sa_ctrl_ia_capability( 
	_zy_simnet_sa_ctrl_ia_capability_327_w$[0:19]), .i_sa_ctrl_ia_status( 
	_zy_simnet_sa_ctrl_ia_status_328_w$[0:12]), .i_sa_ctrl_ia_rdata_part0( 
	_zy_simnet_sa_ctrl_ia_rdata_329_w$[0:31]), .o_reg_written( 
	_zy_simnet_wr_stb_330_w$), .o_reg_read( _zy_simnet_dio_331), 
	.o_reg_wr_data( _zy_simnet_wr_data_332_w$[0:31]), .o_reg_addr( 
	_zy_simnet_reg_addr_333_w$[0:10]));
ixc_assign_32 _zz_strnp_732 ( _zy_simnet_sa_ctrl_ia_wdata_804_w$[0:31], 
	sa_ctrl_ia_wdata[31:0]);
ixc_assign _zz_strnp_731 ( _zy_simnet_wr_stb_803_w$, wr_stb);
ixc_assign_5 _zz_strnp_730 ( _zy_simnet_sa_ctrl_ia_config_802_w$[0:4], 
	sa_ctrl_ia_config[4:0]);
ixc_assign_4 _zz_strnp_729 ( _zy_simnet_sa_ctrl_ia_config_801_w$[0:3], 
	sa_ctrl_ia_config[8:5]);
ixc_assign_11 _zz_strnp_728 ( _zy_simnet_reg_addr_800_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_32 _zz_strnp_727 ( sa_ctrl_ia_rdata[31:0], 
	_zy_simnet_sa_ctrl_ia_rdata_799_w$[0:31]);
ixc_assign_4 _zz_strnp_726 ( sa_ctrl_ia_capability[19:16], 
	_zy_simnet_sa_ctrl_ia_capability_798_w$[0:3]);
ixc_assign_16 _zz_strnp_725 ( sa_ctrl_ia_capability[15:0], 
	_zy_simnet_sa_ctrl_ia_capability_797_w$[0:15]);
ixc_assign_5 _zz_strnp_724 ( sa_ctrl_ia_status[4:0], 
	_zy_simnet_sa_ctrl_ia_status_796_w$[0:4]);
ixc_assign_5 _zz_strnp_723 ( sa_ctrl_ia_status[9:5], 
	_zy_simnet_sa_ctrl_ia_status_795_w$[0:4]);
ixc_assign_3 _zz_strnp_722 ( sa_ctrl_ia_status[12:10], 
	_zy_simnet_sa_ctrl_ia_status_794_w$[0:2]);
ixc_assign_64 _zz_strnp_721 ( _zy_simnet_sa_count_ia_wdata_793_w$[0:63], 
	sa_count_ia_wdata[63:0]);
ixc_assign _zz_strnp_720 ( _zy_simnet_wr_stb_792_w$, wr_stb);
ixc_assign_5 _zz_strnp_719 ( _zy_simnet_sa_count_ia_config_791_w$[0:4], 
	sa_count_ia_config[4:0]);
ixc_assign_4 _zz_strnp_718 ( _zy_simnet_sa_count_ia_config_790_w$[0:3], 
	sa_count_ia_config[8:5]);
ixc_assign_11 _zz_strnp_717 ( _zy_simnet_reg_addr_789_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_64 _zz_strnp_716 ( sa_count_ia_rdata[63:0], 
	_zy_simnet_sa_count_ia_rdata_788_w$[0:63]);
ixc_assign_4 _zz_strnp_715 ( sa_count_ia_capability[19:16], 
	_zy_simnet_sa_count_ia_capability_787_w$[0:3]);
ixc_assign_16 _zz_strnp_714 ( sa_count_ia_capability[15:0], 
	_zy_simnet_sa_count_ia_capability_786_w$[0:15]);
ixc_assign_5 _zz_strnp_713 ( sa_count_ia_status[4:0], 
	_zy_simnet_sa_count_ia_status_785_w$[0:4]);
ixc_assign_5 _zz_strnp_712 ( sa_count_ia_status[9:5], 
	_zy_simnet_sa_count_ia_status_784_w$[0:4]);
ixc_assign_3 _zz_strnp_711 ( sa_count_ia_status[12:10], 
	_zy_simnet_sa_count_ia_status_783_w$[0:2]);
ixc_assign_64 _zz_strnp_710 ( _zy_simnet_sa_snapshot_ia_wdata_782_w$[0:63], 
	sa_snapshot_ia_wdata[63:0]);
ixc_assign _zz_strnp_709 ( _zy_simnet_wr_stb_781_w$, wr_stb);
ixc_assign_5 _zz_strnp_708 ( _zy_simnet_sa_snapshot_ia_config_780_w$[0:4], 
	sa_snapshot_ia_config[4:0]);
ixc_assign_4 _zz_strnp_707 ( _zy_simnet_sa_snapshot_ia_config_779_w$[0:3], 
	sa_snapshot_ia_config[8:5]);
ixc_assign_11 _zz_strnp_706 ( _zy_simnet_reg_addr_778_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_64 _zz_strnp_705 ( sa_snapshot_ia_rdata[63:0], 
	_zy_simnet_sa_snapshot_ia_rdata_777_w$[0:63]);
ixc_assign_4 _zz_strnp_704 ( sa_snapshot_ia_capability[19:16], 
	_zy_simnet_sa_snapshot_ia_capability_776_w$[0:3]);
ixc_assign_16 _zz_strnp_703 ( sa_snapshot_ia_capability[15:0], 
	_zy_simnet_sa_snapshot_ia_capability_775_w$[0:15]);
ixc_assign_5 _zz_strnp_702 ( sa_snapshot_ia_status[4:0], 
	_zy_simnet_sa_snapshot_ia_status_774_w$[0:4]);
ixc_assign_5 _zz_strnp_701 ( sa_snapshot_ia_status[9:5], 
	_zy_simnet_sa_snapshot_ia_status_773_w$[0:4]);
ixc_assign_3 _zz_strnp_700 ( sa_snapshot_ia_status[12:10], 
	_zy_simnet_sa_snapshot_ia_status_772_w$[0:2]);
ixc_assign_5 _zz_strnp_699 ( _zy_simnet_o_interrupt_mask_771_w$[0:4], 
	o_interrupt_mask[4:0]);
ixc_assign_11 _zz_strnp_698 ( _zy_simnet_reg_addr_770_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_32 _zz_strnp_697 ( _zy_simnet_wr_data_769_w$[0:31], wr_data[31:0]);
ixc_assign _zz_strnp_696 ( _zy_simnet_wr_stb_768_w$, wr_stb);
ixc_assign _zz_strnp_695 ( _zy_simnet_bimc_interrupt_767_w$, bimc_interrupt);
ixc_assign _zz_strnp_694 ( _zy_simnet_cddip3_ism_mbe_766_w$, cddip3_ism_mbe);
ixc_assign _zz_strnp_693 ( _zy_simnet_cddip2_ism_mbe_765_w$, cddip2_ism_mbe);
ixc_assign _zz_strnp_692 ( _zy_simnet_cddip1_ism_mbe_764_w$, cddip1_ism_mbe);
ixc_assign _zz_strnp_691 ( _zy_simnet_cddip0_ism_mbe_763_w$, cddip0_ism_mbe);
ixc_assign _zz_strnp_690 ( _zy_simnet_cceip3_ism_mbe_762_w$, cceip3_ism_mbe);
ixc_assign _zz_strnp_689 ( _zy_simnet_cceip2_ism_mbe_761_w$, cceip2_ism_mbe);
ixc_assign _zz_strnp_688 ( _zy_simnet_cceip1_ism_mbe_760_w$, cceip1_ism_mbe);
ixc_assign _zz_strnp_687 ( _zy_simnet_cceip0_ism_mbe_759_w$, cceip0_ism_mbe);
ixc_assign _zz_strnp_686 ( _zy_simnet_set_drbg_expired_int_758_w$, 
	set_drbg_expired_int);
ixc_assign_5 _zz_strnp_685 ( interrupt_status[4:0], 
	_zy_simnet_interrupt_status_757_w$[0:4]);
ixc_assign_32 _zz_strnp_684 ( bimc_dbgcmd0[31:0], 
	_zy_simnet_bimc_dbgcmd0_756_w$[0:31]);
ixc_assign_32 _zz_strnp_683 ( bimc_dbgcmd1[31:0], 
	_zy_simnet_bimc_dbgcmd1_755_w$[0:31]);
ixc_assign_10 _zz_strnp_682 ( bimc_dbgcmd2[9:0], 
	_zy_simnet_bimc_dbgcmd2_754_w$[0:9]);
ixc_assign_32 _zz_strnp_681 ( bimc_pollrsp0[31:0], 
	_zy_simnet_bimc_pollrsp0_753_w$[0:31]);
ixc_assign_32 _zz_strnp_680 ( bimc_pollrsp1[31:0], 
	_zy_simnet_bimc_pollrsp1_752_w$[0:31]);
ixc_assign_10 _zz_strnp_679 ( bimc_pollrsp2[9:0], 
	_zy_simnet_bimc_pollrsp2_751_w$[0:9]);
ixc_assign_32 _zz_strnp_678 ( bimc_rxrsp0[31:0], 
	_zy_simnet_bimc_rxrsp0_750_w$[0:31]);
ixc_assign_32 _zz_strnp_677 ( bimc_rxrsp1[31:0], 
	_zy_simnet_bimc_rxrsp1_749_w$[0:31]);
ixc_assign_10 _zz_strnp_676 ( bimc_rxrsp2[9:0], 
	_zy_simnet_bimc_rxrsp2_748_w$[0:9]);
ixc_assign_32 _zz_strnp_675 ( bimc_rxcmd0[31:0], 
	_zy_simnet_bimc_rxcmd0_747_w$[0:31]);
ixc_assign_32 _zz_strnp_674 ( bimc_rxcmd1[31:0], 
	_zy_simnet_bimc_rxcmd1_746_w$[0:31]);
ixc_assign_10 _zz_strnp_673 ( bimc_rxcmd2[9:0], 
	_zy_simnet_bimc_rxcmd2_745_w$[0:9]);
ixc_assign_11 _zz_strnp_672 ( bimc_cmd2[10:0], 
	_zy_simnet_bimc_cmd2_744_w$[0:10]);
ixc_assign_29 _zz_strnp_671 ( bimc_eccpar_debug[28:0], 
	_zy_simnet_bimc_eccpar_debug_743_w$[0:28]);
ixc_assign_12 _zz_strnp_670 ( bimc_memid[11:0], 
	_zy_simnet_bimc_memid_742_w$[0:11]);
ixc_assign_32 _zz_strnp_669 ( bimc_global_config[31:0], 
	_zy_simnet_bimc_global_config_741_w$[0:31]);
ixc_assign_32 _zz_strnp_668 ( bimc_parity_error_cnt[31:0], 
	_zy_simnet_bimc_parity_error_cnt_740_w$[0:31]);
ixc_assign_32 _zz_strnp_667 ( bimc_ecc_correctable_error_cnt[31:0], 
	_zy_simnet_bimc_ecc_correctable_error_cnt_739_w$[0:31]);
ixc_assign_32 _zz_strnp_666 ( bimc_ecc_uncorrectable_error_cnt[31:0], 
	_zy_simnet_bimc_ecc_uncorrectable_error_cnt_738_w$[0:31]);
ixc_assign_7 _zz_strnp_665 ( bimc_monitor[6:0], 
	_zy_simnet_bimc_monitor_737_w$[0:6]);
ixc_assign_10 _zz_strnp_664 ( _zy_simnet_o_bimc_dbgcmd2_736_w$[0:9], 
	o_bimc_dbgcmd2[9:0]);
ixc_assign_10 _zz_strnp_663 ( _zy_simnet_o_bimc_pollrsp2_735_w$[0:9], 
	o_bimc_pollrsp2[9:0]);
ixc_assign_10 _zz_strnp_662 ( _zy_simnet_o_bimc_rxrsp2_734_w$[0:9], 
	o_bimc_rxrsp2[9:0]);
ixc_assign_10 _zz_strnp_661 ( _zy_simnet_o_bimc_rxcmd2_733_w$[0:9], 
	o_bimc_rxcmd2[9:0]);
ixc_assign_32 _zz_strnp_660 ( _zy_simnet_o_bimc_cmd0_732_w$[0:31], 
	o_bimc_cmd0[31:0]);
ixc_assign_32 _zz_strnp_659 ( _zy_simnet_o_bimc_cmd1_731_w$[0:31], 
	o_bimc_cmd1[31:0]);
ixc_assign_11 _zz_strnp_658 ( _zy_simnet_o_bimc_cmd2_730_w$[0:10], 
	o_bimc_cmd2[10:0]);
ixc_assign_29 _zz_strnp_657 ( _zy_simnet_o_bimc_eccpar_debug_729_w$[0:28], 
	o_bimc_eccpar_debug[28:0]);
ixc_assign_32 _zz_strnp_656 ( _zy_simnet_o_bimc_global_config_728_w$[0:31], 
	o_bimc_global_config[31:0]);
ixc_assign_32 _zz_strnp_655 ( _zy_simnet_o_bimc_parity_error_cnt_727_w$[0:31], 
	o_bimc_parity_error_cnt[31:0]);
ixc_assign_32 _zz_strnp_654 ( 
	_zy_simnet_o_bimc_ecc_correctable_error_cnt_726_w$[0:31], 
	o_bimc_ecc_correctable_error_cnt[31:0]);
ixc_assign_32 _zz_strnp_653 ( 
	_zy_simnet_o_bimc_ecc_uncorrectable_error_cnt_725_w$[0:31], 
	o_bimc_ecc_uncorrectable_error_cnt[31:0]);
ixc_assign_7 _zz_strnp_652 ( _zy_simnet_o_bimc_monitor_mask_724_w$[0:6], 
	o_bimc_monitor_mask[6:0]);
ixc_assign _zz_strnp_651 ( _zy_simnet_axi_term_bimc_isync_723_w$, 
	axi_term_bimc_isync);
ixc_assign _zz_strnp_650 ( _zy_simnet_axi_term_bimc_idat_722_w$, 
	axi_term_bimc_idat);
ixc_assign _zz_strnp_649 ( kim_bimc_isync, _zy_simnet_kim_bimc_isync_721_w$);
ixc_assign _zz_strnp_648 ( kim_bimc_idat, _zy_simnet_kim_bimc_idat_720_w$);
ixc_assign _zz_strnp_647 ( bimc_interrupt, _zy_simnet_bimc_interrupt_719_w$);
ixc_assign_32 _zz_strnp_646 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_95_64_717_w$[0:31], 
	o_kdf_drbg_seed_1_state_value_95_64[31:0]);
ixc_assign_32 _zz_strnp_645 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_63_32_716_w$[0:31], 
	o_kdf_drbg_seed_1_state_value_63_32[31:0]);
ixc_assign_32 _zz_strnp_644 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_31_0_715_w$[0:31], 
	o_kdf_drbg_seed_1_state_value_31_0[31:0]);
ixc_assign_32 _zz_strnp_643 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_127_96_714_w$[0:31], 
	o_kdf_drbg_seed_1_state_value_127_96[31:0]);
ixc_assign_32 _zz_strnp_642 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_95_64_713_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_95_64[31:0]);
ixc_assign_32 _zz_strnp_641 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_63_32_712_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_63_32[31:0]);
ixc_assign_32 _zz_strnp_640 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_31_0_711_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_31_0[31:0]);
ixc_assign_32 _zz_strnp_639 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_255_224_710_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_255_224[31:0]);
ixc_assign_32 _zz_strnp_638 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_223_192_709_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_223_192[31:0]);
ixc_assign_32 _zz_strnp_637 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_191_160_708_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_191_160[31:0]);
ixc_assign_32 _zz_strnp_636 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_159_128_707_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_159_128[31:0]);
ixc_assign_32 _zz_strnp_635 ( 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_127_96_706_w$[0:31], 
	o_kdf_drbg_seed_1_state_key_127_96[31:0]);
ixc_assign_16 _zz_strnp_634 ( 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_1_705_w$[0:15], 
	o_kdf_drbg_seed_1_reseed_interval_1[15:0]);
ixc_assign_32 _zz_strnp_633 ( 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_0_704_w$[0:31], 
	o_kdf_drbg_seed_1_reseed_interval_0[31:0]);
ixc_assign_32 _zz_strnp_632 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_95_64_703_w$[0:31], 
	o_kdf_drbg_seed_0_state_value_95_64[31:0]);
ixc_assign_32 _zz_strnp_631 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_63_32_702_w$[0:31], 
	o_kdf_drbg_seed_0_state_value_63_32[31:0]);
ixc_assign_32 _zz_strnp_630 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_31_0_701_w$[0:31], 
	o_kdf_drbg_seed_0_state_value_31_0[31:0]);
ixc_assign_32 _zz_strnp_629 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_127_96_700_w$[0:31], 
	o_kdf_drbg_seed_0_state_value_127_96[31:0]);
ixc_assign_32 _zz_strnp_628 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_95_64_699_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_95_64[31:0]);
ixc_assign_32 _zz_strnp_627 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_63_32_698_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_63_32[31:0]);
ixc_assign_32 _zz_strnp_626 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_31_0_697_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_31_0[31:0]);
ixc_assign_32 _zz_strnp_625 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_255_224_696_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_255_224[31:0]);
ixc_assign_32 _zz_strnp_624 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_223_192_695_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_223_192[31:0]);
ixc_assign_32 _zz_strnp_623 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_191_160_694_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_191_160[31:0]);
ixc_assign_32 _zz_strnp_622 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_159_128_693_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_159_128[31:0]);
ixc_assign_32 _zz_strnp_621 ( 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_127_96_692_w$[0:31], 
	o_kdf_drbg_seed_0_state_key_127_96[31:0]);
ixc_assign_16 _zz_strnp_620 ( 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_1_691_w$[0:15], 
	o_kdf_drbg_seed_0_reseed_interval_1[15:0]);
ixc_assign_32 _zz_strnp_619 ( 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_0_690_w$[0:31], 
	o_kdf_drbg_seed_0_reseed_interval_0[31:0]);
ixc_assign_2 _zz_strnp_618 ( _zy_simnet_o_kdf_drbg_ctrl_689_w$[0:1], 
	o_kdf_drbg_ctrl[1:0]);
ixc_assign_11 _zz_strnp_617 ( _zy_simnet_reg_addr_688_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_32 _zz_strnp_616 ( _zy_simnet_wr_data_687_w$[0:31], wr_data[31:0]);
ixc_assign _zz_strnp_615 ( _zy_simnet_wr_stb_686_w$, wr_stb);
ixc_assign_2 _zz_strnp_614 ( kdf_drbg_ctrl[1:0], 
	_zy_simnet_kdf_drbg_ctrl_685_w$[0:1]);
ixc_assign _zz_strnp_613 ( set_drbg_expired_int, 
	_zy_simnet_set_drbg_expired_int_684_w$);
ixc_assign_38 _zz_strnp_612 ( kim_dout[37:0], 
	_zy_simnet_kim_dout_682_w$[0:37]);
ixc_assign _zz_strnp_611 ( ckv_bimc_isync, _zy_simnet_ckv_bimc_isync_678_w$);
ixc_assign _zz_strnp_610 ( ckv_bimc_idat, _zy_simnet_ckv_bimc_idat_677_w$);
ixc_assign _zz_strnp_609 ( _zy_simnet_kim_bimc_idat_676_w$, kim_bimc_idat);
ixc_assign _zz_strnp_608 ( _zy_simnet_kim_bimc_isync_675_w$, kim_bimc_isync);
ixc_assign_38 _zz_strnp_607 ( kim_rd_dat[37:0], 
	_zy_simnet_kim_rd_dat_673_w$[0:37]);
ixc_assign_38 _zz_strnp_606 ( _zy_simnet_kim_wr_dat_672_w$[0:37], 
	kim_wr_dat[37:0]);
ixc_assign _zz_strnp_605 ( _zy_simnet_wr_stb_671_w$, wr_stb);
ixc_assign_4 _zz_strnp_604 ( kim_capability_type[3:0], 
	_zy_simnet_kim_capability_type_670_w$[0:3]);
ixc_assign_16 _zz_strnp_603 ( kim_capability_lst[15:0], 
	_zy_simnet_kim_capability_lst_669_w$[0:15]);
ixc_assign_14 _zz_strnp_602 ( kim_stat_addr[13:0], 
	_zy_simnet_kim_stat_addr_668_w$[0:13]);
ixc_assign_5 _zz_strnp_601 ( kim_stat_datawords[4:0], 
	_zy_simnet_kim_stat_datawords_667_w$[0:4]);
ixc_assign_3 _zz_strnp_600 ( kim_stat_code[2:0], 
	_zy_simnet_kim_stat_code_666_w$[0:2]);
ixc_assign_14 _zz_strnp_599 ( _zy_simnet_kim_cmnd_addr_665_w$[0:13], 
	kim_cmnd_addr[13:0]);
ixc_assign_4 _zz_strnp_598 ( _zy_simnet_kim_cmnd_op_664_w$[0:3], 
	kim_cmnd_op[3:0]);
ixc_assign_11 _zz_strnp_597 ( _zy_simnet_reg_addr_663_w$[0:10], 
	reg_addr[10:0]);
ixc_assign _zz_strnp_596 ( cceip0_ism_bimc_isync, 
	_zy_simnet_cceip0_ism_bimc_isync_658_w$);
ixc_assign _zz_strnp_595 ( cceip0_ism_bimc_idat, 
	_zy_simnet_cceip0_ism_bimc_idat_657_w$);
ixc_assign _zz_strnp_594 ( _zy_simnet_ckv_bimc_idat_656_w$, ckv_bimc_idat);
ixc_assign _zz_strnp_593 ( _zy_simnet_ckv_bimc_isync_655_w$, ckv_bimc_isync);
ixc_assign_64 _zz_strnp_592 ( ckv_rd_dat[63:0], 
	_zy_simnet_ckv_rd_dat_653_w$[0:63]);
ixc_assign_64 _zz_strnp_591 ( _zy_simnet_ckv_wr_dat_652_w$[0:63], 
	ckv_wr_dat[63:0]);
ixc_assign _zz_strnp_590 ( _zy_simnet_wr_stb_651_w$, wr_stb);
ixc_assign_4 _zz_strnp_589 ( ckv_capability_type[3:0], 
	_zy_simnet_ckv_capability_type_650_w$[0:3]);
ixc_assign_16 _zz_strnp_588 ( ckv_capability_lst[15:0], 
	_zy_simnet_ckv_capability_lst_649_w$[0:15]);
ixc_assign_15 _zz_strnp_587 ( ckv_stat_addr[14:0], 
	_zy_simnet_ckv_stat_addr_648_w$[0:14]);
ixc_assign_5 _zz_strnp_586 ( ckv_stat_datawords[4:0], 
	_zy_simnet_ckv_stat_datawords_647_w$[0:4]);
ixc_assign_3 _zz_strnp_585 ( ckv_stat_code[2:0], 
	_zy_simnet_ckv_stat_code_646_w$[0:2]);
ixc_assign_15 _zz_strnp_584 ( _zy_simnet_ckv_cmnd_addr_645_w$[0:14], 
	ckv_cmnd_addr[14:0]);
ixc_assign_4 _zz_strnp_583 ( _zy_simnet_ckv_cmnd_op_644_w$[0:3], 
	ckv_cmnd_op[3:0]);
ixc_assign_11 _zz_strnp_582 ( _zy_simnet_reg_addr_643_w$[0:10], 
	reg_addr[10:0]);
ixc_assign _zz_strnp_581 ( _zy_simnet_cddip3_ism_odat_642_w$, cddip3_ism_odat);
ixc_assign _zz_strnp_580 ( _zy_simnet_cddip3_ism_osync_641_w$, 
	cddip3_ism_osync);
ixc_assign_83 _zz_strnp_579 ( _zy_simnet_kme_cddip3_ob_out_post_640_w$[0:82], 
	kme_cddip3_ob_out_post[82:0]);
ixc_assign_83 _zz_strnp_578 ( _zy_simnet_kme_cddip2_ob_out_post_639_w$[0:82], 
	kme_cddip2_ob_out_post[82:0]);
ixc_assign_83 _zz_strnp_577 ( _zy_simnet_kme_cddip1_ob_out_post_638_w$[0:82], 
	kme_cddip1_ob_out_post[82:0]);
ixc_assign_83 _zz_strnp_576 ( _zy_simnet_kme_cddip0_ob_out_post_637_w$[0:82], 
	kme_cddip0_ob_out_post[82:0]);
ixc_assign_83 _zz_strnp_575 ( _zy_simnet_kme_cceip3_ob_out_post_636_w$[0:82], 
	kme_cceip3_ob_out_post[82:0]);
ixc_assign_83 _zz_strnp_574 ( _zy_simnet_kme_cceip2_ob_out_post_635_w$[0:82], 
	kme_cceip2_ob_out_post[82:0]);
ixc_assign_83 _zz_strnp_573 ( _zy_simnet_kme_cceip1_ob_out_post_634_w$[0:82], 
	kme_cceip1_ob_out_post[82:0]);
ixc_assign_83 _zz_strnp_572 ( _zy_simnet_kme_cceip0_ob_out_post_633_w$[0:82], 
	kme_cceip0_ob_out_post[82:0]);
ixc_assign_9 _zz_strnp_571 ( _zy_simnet_tready_override_632_w$[0:8], 
	tready_override[8:0]);
ixc_assign_96 _zz_strnp_570 ( _zy_simnet_cceip0_out_ia_wdata_631_w$[0:95], 
	cceip0_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_569 ( _zy_simnet_o_send_kme_ib_beat_630_w$, 
	o_send_kme_ib_beat);
ixc_assign _zz_strnp_568 ( _zy_simnet_o_disable_ckv_kim_ism_reads_629_w$, 
	o_disable_ckv_kim_ism_reads);
ixc_assign_8 _zz_strnp_567 ( _zy_simnet_o_engine_sticky_status_628_w$[0:7], 
	o_engine_sticky_status[7:0]);
ixc_assign_11 _zz_strnp_566 ( _zy_simnet_reg_addr_627_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_32 _zz_strnp_565 ( _zy_simnet_wr_data_626_w$[0:31], wr_data[31:0]);
ixc_assign _zz_strnp_564 ( _zy_simnet_wr_stb_625_w$, wr_stb);
ixc_assign_17 _zz_strnp_563 ( _zy_simnet_o_kim_ia_wdata_part1_624_w$[0:16], 
	o_kim_ia_wdata_part1[16:0]);
ixc_assign_21 _zz_strnp_562 ( _zy_simnet_o_kim_ia_wdata_part0_623_w$[0:20], 
	o_kim_ia_wdata_part0[20:0]);
ixc_assign_18 _zz_strnp_561 ( _zy_simnet_o_kim_ia_config_622_w$[0:17], 
	o_kim_ia_config[17:0]);
ixc_assign_38 _zz_strnp_560 ( _zy_simnet_kim_rd_dat_621_w$[0:37], 
	kim_rd_dat[37:0]);
ixc_assign_16 _zz_strnp_559 ( _zy_simnet_kim_capability_lst_620_w$[0:15], 
	kim_capability_lst[15:0]);
ixc_assign_4 _zz_strnp_558 ( _zy_simnet_kim_capability_type_619_w$[0:3], 
	kim_capability_type[3:0]);
ixc_assign_14 _zz_strnp_557 ( _zy_simnet_kim_stat_addr_618_w$[0:13], 
	kim_stat_addr[13:0]);
ixc_assign_5 _zz_strnp_556 ( _zy_simnet_kim_stat_datawords_617_w$[0:4], 
	kim_stat_datawords[4:0]);
ixc_assign_3 _zz_strnp_555 ( _zy_simnet_kim_stat_code_616_w$[0:2], 
	kim_stat_code[2:0]);
ixc_assign_32 _zz_strnp_554 ( _zy_simnet_o_ckv_ia_wdata_part1_615_w$[0:31], 
	o_ckv_ia_wdata_part1[31:0]);
ixc_assign_32 _zz_strnp_553 ( _zy_simnet_o_ckv_ia_wdata_part0_614_w$[0:31], 
	o_ckv_ia_wdata_part0[31:0]);
ixc_assign_19 _zz_strnp_552 ( _zy_simnet_o_ckv_ia_config_613_w$[0:18], 
	o_ckv_ia_config[18:0]);
ixc_assign_64 _zz_strnp_551 ( _zy_simnet_ckv_rd_dat_612_w$[0:63], 
	ckv_rd_dat[63:0]);
ixc_assign_16 _zz_strnp_550 ( _zy_simnet_ckv_capability_lst_611_w$[0:15], 
	ckv_capability_lst[15:0]);
ixc_assign_4 _zz_strnp_549 ( _zy_simnet_ckv_capability_type_610_w$[0:3], 
	ckv_capability_type[3:0]);
ixc_assign_15 _zz_strnp_548 ( _zy_simnet_ckv_stat_addr_609_w$[0:14], 
	ckv_stat_addr[14:0]);
ixc_assign_5 _zz_strnp_547 ( _zy_simnet_ckv_stat_datawords_608_w$[0:4], 
	ckv_stat_datawords[4:0]);
ixc_assign_3 _zz_strnp_546 ( _zy_simnet_ckv_stat_code_607_w$[0:2], 
	ckv_stat_code[2:0]);
ixc_assign _zz_strnp_545 ( axi_term_bimc_idat, 
	_zy_simnet_axi_term_bimc_idat_606_w$);
ixc_assign _zz_strnp_544 ( axi_term_bimc_isync, 
	_zy_simnet_axi_term_bimc_isync_605_w$);
ixc_assign_83 _zz_strnp_543 ( kme_cddip3_ob_out[82:0], 
	_zy_simnet_kme_cddip3_ob_out_604_w$[0:82]);
ixc_assign_83 _zz_strnp_542 ( kme_cddip2_ob_out[82:0], 
	_zy_simnet_kme_cddip2_ob_out_603_w$[0:82]);
ixc_assign_83 _zz_strnp_541 ( kme_cddip1_ob_out[82:0], 
	_zy_simnet_kme_cddip1_ob_out_602_w$[0:82]);
ixc_assign_83 _zz_strnp_540 ( kme_cddip0_ob_out[82:0], 
	_zy_simnet_kme_cddip0_ob_out_601_w$[0:82]);
ixc_assign_83 _zz_strnp_539 ( kme_cceip3_ob_out[82:0], 
	_zy_simnet_kme_cceip3_ob_out_600_w$[0:82]);
ixc_assign_83 _zz_strnp_538 ( kme_cceip2_ob_out[82:0], 
	_zy_simnet_kme_cceip2_ob_out_599_w$[0:82]);
ixc_assign_83 _zz_strnp_537 ( kme_cceip1_ob_out[82:0], 
	_zy_simnet_kme_cceip1_ob_out_598_w$[0:82]);
ixc_assign_83 _zz_strnp_536 ( kme_cceip0_ob_out[82:0], 
	_zy_simnet_kme_cceip0_ob_out_597_w$[0:82]);
ixc_assign _zz_strnp_535 ( send_kme_ib_beat, 
	_zy_simnet_send_kme_ib_beat_596_w$);
ixc_assign _zz_strnp_534 ( disable_ckv_kim_ism_reads, 
	_zy_simnet_disable_ckv_kim_ism_reads_595_w$);
ixc_assign_8 _zz_strnp_533 ( engine_sticky_status[7:0], 
	_zy_simnet_engine_sticky_status_594_w$[0:7]);
ixc_assign_22 _zz_strnp_532 ( kim_ia_status[21:0], 
	_zy_simnet_kim_ia_status_593_w$[0:21]);
ixc_assign_17 _zz_strnp_531 ( kim_ia_rdata_part1[16:0], 
	_zy_simnet_kim_ia_rdata_part1_592_w$[0:16]);
ixc_assign_21 _zz_strnp_530 ( kim_ia_rdata_part0[20:0], 
	_zy_simnet_kim_ia_rdata_part0_591_w$[0:20]);
ixc_assign_20 _zz_strnp_529 ( kim_ia_capability[19:0], 
	_zy_simnet_kim_ia_capability_590_w$[0:19]);
ixc_assign_38 _zz_strnp_528 ( kim_wr_dat[37:0], 
	_zy_simnet_kim_wr_dat_589_w$[0:37]);
ixc_assign_14 _zz_strnp_527 ( kim_cmnd_addr[13:0], 
	_zy_simnet_kim_cmnd_addr_588_w$[0:13]);
ixc_assign_4 _zz_strnp_526 ( kim_cmnd_op[3:0], 
	_zy_simnet_kim_cmnd_op_587_w$[0:3]);
ixc_assign_23 _zz_strnp_525 ( ckv_ia_status[22:0], 
	_zy_simnet_ckv_ia_status_586_w$[0:22]);
ixc_assign_32 _zz_strnp_524 ( ckv_ia_rdata_part1[31:0], 
	_zy_simnet_ckv_ia_rdata_part1_585_w$[0:31]);
ixc_assign_32 _zz_strnp_523 ( ckv_ia_rdata_part0[31:0], 
	_zy_simnet_ckv_ia_rdata_part0_584_w$[0:31]);
ixc_assign_20 _zz_strnp_522 ( ckv_ia_capability[19:0], 
	_zy_simnet_ckv_ia_capability_583_w$[0:19]);
ixc_assign_64 _zz_strnp_521 ( ckv_wr_dat[63:0], 
	_zy_simnet_ckv_wr_dat_582_w$[0:63]);
ixc_assign_15 _zz_strnp_520 ( ckv_cmnd_addr[14:0], 
	_zy_simnet_ckv_cmnd_addr_581_w$[0:14]);
ixc_assign_4 _zz_strnp_519 ( ckv_cmnd_op[3:0], 
	_zy_simnet_ckv_cmnd_op_580_w$[0:3]);
ixc_assign_12 _zz_strnp_518 ( _zy_simnet_cddip3_out_im_config_579_w$[0:11], 
	cddip3_out_im_config[11:0]);
ixc_assign_2 _zz_strnp_517 ( _zy_simnet_im_consumed_kme_cddip3_578_w$[0:1], 
	im_consumed_kme_cddip3[1:0]);
ixc_assign _zz_strnp_516 ( _zy_simnet_cddip3_im_vld_577_w$, cddip3_im_vld);
ixc_assign_96 _zz_strnp_515 ( _zy_simnet_cddip3_im_din_576_w$[0:95], { 
	cddip3_im_din[95], cddip3_im_din[94], cddip3_im_din[93], 
	cddip3_im_din[92], cddip3_im_din[91], cddip3_im_din[90], 
	cddip3_im_din[89], cddip3_im_din[88], cddip3_im_din[87], 
	cddip3_im_din[86], cddip3_im_din[85], cddip3_im_din[84], 
	cddip3_im_din[83], cddip3_im_din[82], cddip3_im_din[81], 
	cddip3_im_din[80], cddip3_im_din[79], cddip3_im_din[78], 
	cddip3_im_din[77], cddip3_im_din[76], cddip3_im_din[75], 
	cddip3_im_din[74], cddip3_im_din[73], cddip3_im_din[72], 
	cddip3_im_din[71], cddip3_im_din[70], cddip3_im_din[69], 
	cddip3_im_din[68], cddip3_im_din[67], cddip3_im_din[66], 
	cddip3_im_din[65], cddip3_im_din[64], cddip3_im_din[63], 
	cddip3_im_din[62], cddip3_im_din[61], cddip3_im_din[60], 
	cddip3_im_din[59], cddip3_im_din[58], cddip3_im_din[57], 
	cddip3_im_din[56], cddip3_im_din[55], cddip3_im_din[54], 
	cddip3_im_din[53], cddip3_im_din[52], cddip3_im_din[51], 
	cddip3_im_din[50], cddip3_im_din[49], cddip3_im_din[48], 
	cddip3_im_din[47], cddip3_im_din[46], cddip3_im_din[45], 
	cddip3_im_din[44], cddip3_im_din[43], cddip3_im_din[42], 
	cddip3_im_din[41], cddip3_im_din[40], cddip3_im_din[39], 
	cddip3_im_din[38], cddip3_im_din[37], cddip3_im_din[36], 
	cddip3_im_din[35], cddip3_im_din[34], cddip3_im_din[33], 
	cddip3_im_din[32], kme_cddip3_ob_out_pre[65], cddip3_im_din[30], 
	cddip3_im_din[29], cddip3_im_din[28], cddip3_im_din[27], 
	cddip3_im_din[26], cddip3_im_din[25], cddip3_im_din[24], 
	cddip3_im_din[23], cddip3_im_din[22], cddip3_im_din[21], 
	cddip3_im_din[20], cddip3_im_din[19], cddip3_im_din[18], 
	cddip3_im_din[17], cddip3_im_din[16], cddip3_im_din[15], 
	cddip3_im_din[14], cddip3_im_din[13], cddip3_im_din[12], 
	cddip3_im_din[11], cddip3_im_din[10], cddip3_im_din[9], 
	cddip3_im_din[8], kme_cddip3_ob_out_pre[65], cddip3_im_din[6], 
	cddip3_im_din[5], cddip3_im_din[4], cddip3_im_din[3], 
	cddip3_im_din[2], cddip3_im_din[1], cddip3_im_din[0]});
ixc_assign _zz_strnp_514 ( _zy_simnet_cddip3_ism_idat_575_w$, cddip3_ism_idat);
ixc_assign _zz_strnp_513 ( _zy_simnet_cddip3_ism_isync_574_w$, 
	cddip3_ism_isync);
ixc_assign_96 _zz_strnp_512 ( _zy_simnet_cddip3_out_ia_wdata_572_w$[0:95], 
	cddip3_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_511 ( _zy_simnet_wr_stb_571_w$, wr_stb);
ixc_assign_9 _zz_strnp_510 ( _zy_simnet_cddip3_out_ia_config_570_w$[0:8], 
	cddip3_out_ia_config[8:0]);
ixc_assign_4 _zz_strnp_509 ( _zy_simnet_cddip3_out_ia_config_569_w$[0:3], 
	cddip3_out_ia_config[12:9]);
ixc_assign_11 _zz_strnp_508 ( _zy_simnet_reg_addr_568_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_12 _zz_strnp_507 ( cddip3_out_im_status[11:0], 
	_zy_simnet_cddip3_out_im_status_567_w$[0:11]);
ixc_assign_2 _zz_strnp_506 ( im_available_kme_cddip3[1:0], 
	_zy_simnet_im_available_kme_cddip3_566_w$[0:1]);
ixc_assign _zz_strnp_505 ( cddip3_im_rdy, _zy_simnet_cddip3_im_rdy_565_w$);
ixc_assign _zz_strnp_504 ( cddip3_ism_mbe, _zy_simnet_cddip3_ism_mbe_564_w$);
ixc_assign _zz_strnp_503 ( cddip3_ism_osync, 
	_zy_simnet_cddip3_ism_osync_563_w$);
ixc_assign _zz_strnp_502 ( cddip3_ism_odat, _zy_simnet_cddip3_ism_odat_562_w$);
ixc_assign_96 _zz_strnp_501 ( cddip3_out_ia_rdata[95:0], 
	_zy_simnet_cddip3_out_ia_rdata_561_w$[0:95]);
ixc_assign_4 _zz_strnp_500 ( cddip3_out_ia_capability[19:16], 
	_zy_simnet_cddip3_out_ia_capability_560_w$[0:3]);
ixc_assign_16 _zz_strnp_499 ( cddip3_out_ia_capability[15:0], 
	_zy_simnet_cddip3_out_ia_capability_559_w$[0:15]);
ixc_assign_9 _zz_strnp_498 ( cddip3_out_ia_status[8:0], 
	_zy_simnet_cddip3_out_ia_status_558_w$[0:8]);
ixc_assign_5 _zz_strnp_497 ( cddip3_out_ia_status[13:9], 
	_zy_simnet_cddip3_out_ia_status_557_w$[0:4]);
ixc_assign_3 _zz_strnp_496 ( cddip3_out_ia_status[16:14], 
	_zy_simnet_cddip3_out_ia_status_556_w$[0:2]);
ixc_assign_12 _zz_strnp_495 ( _zy_simnet_cddip2_out_im_config_555_w$[0:11], 
	cddip2_out_im_config[11:0]);
ixc_assign_2 _zz_strnp_494 ( _zy_simnet_im_consumed_kme_cddip2_554_w$[0:1], 
	im_consumed_kme_cddip2[1:0]);
ixc_assign _zz_strnp_493 ( _zy_simnet_cddip2_im_vld_553_w$, cddip2_im_vld);
ixc_assign_96 _zz_strnp_492 ( _zy_simnet_cddip2_im_din_552_w$[0:95], { 
	cddip2_im_din[95], cddip2_im_din[94], cddip2_im_din[93], 
	cddip2_im_din[92], cddip2_im_din[91], cddip2_im_din[90], 
	cddip2_im_din[89], cddip2_im_din[88], cddip2_im_din[87], 
	cddip2_im_din[86], cddip2_im_din[85], cddip2_im_din[84], 
	cddip2_im_din[83], cddip2_im_din[82], cddip2_im_din[81], 
	cddip2_im_din[80], cddip2_im_din[79], cddip2_im_din[78], 
	cddip2_im_din[77], cddip2_im_din[76], cddip2_im_din[75], 
	cddip2_im_din[74], cddip2_im_din[73], cddip2_im_din[72], 
	cddip2_im_din[71], cddip2_im_din[70], cddip2_im_din[69], 
	cddip2_im_din[68], cddip2_im_din[67], cddip2_im_din[66], 
	cddip2_im_din[65], cddip2_im_din[64], cddip2_im_din[63], 
	cddip2_im_din[62], cddip2_im_din[61], cddip2_im_din[60], 
	cddip2_im_din[59], cddip2_im_din[58], cddip2_im_din[57], 
	cddip2_im_din[56], cddip2_im_din[55], cddip2_im_din[54], 
	cddip2_im_din[53], cddip2_im_din[52], cddip2_im_din[51], 
	cddip2_im_din[50], cddip2_im_din[49], cddip2_im_din[48], 
	cddip2_im_din[47], cddip2_im_din[46], cddip2_im_din[45], 
	cddip2_im_din[44], cddip2_im_din[43], cddip2_im_din[42], 
	cddip2_im_din[41], cddip2_im_din[40], cddip2_im_din[39], 
	cddip2_im_din[38], cddip2_im_din[37], cddip2_im_din[36], 
	cddip2_im_din[35], cddip2_im_din[34], cddip2_im_din[33], 
	cddip2_im_din[32], kme_cddip2_ob_out_pre[65], cddip2_im_din[30], 
	cddip2_im_din[29], cddip2_im_din[28], cddip2_im_din[27], 
	cddip2_im_din[26], cddip2_im_din[25], cddip2_im_din[24], 
	cddip2_im_din[23], cddip2_im_din[22], cddip2_im_din[21], 
	cddip2_im_din[20], cddip2_im_din[19], cddip2_im_din[18], 
	cddip2_im_din[17], cddip2_im_din[16], cddip2_im_din[15], 
	cddip2_im_din[14], cddip2_im_din[13], cddip2_im_din[12], 
	cddip2_im_din[11], cddip2_im_din[10], cddip2_im_din[9], 
	cddip2_im_din[8], kme_cddip2_ob_out_pre[65], cddip2_im_din[6], 
	cddip2_im_din[5], cddip2_im_din[4], cddip2_im_din[3], 
	cddip2_im_din[2], cddip2_im_din[1], cddip2_im_din[0]});
ixc_assign _zz_strnp_491 ( _zy_simnet_cddip2_ism_idat_551_w$, cddip2_ism_idat);
ixc_assign _zz_strnp_490 ( _zy_simnet_cddip2_ism_isync_550_w$, 
	cddip2_ism_isync);
ixc_assign_96 _zz_strnp_489 ( _zy_simnet_cddip2_out_ia_wdata_548_w$[0:95], 
	cddip2_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_488 ( _zy_simnet_wr_stb_547_w$, wr_stb);
ixc_assign_9 _zz_strnp_487 ( _zy_simnet_cddip2_out_ia_config_546_w$[0:8], 
	cddip2_out_ia_config[8:0]);
ixc_assign_4 _zz_strnp_486 ( _zy_simnet_cddip2_out_ia_config_545_w$[0:3], 
	cddip2_out_ia_config[12:9]);
ixc_assign_11 _zz_strnp_485 ( _zy_simnet_reg_addr_544_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_12 _zz_strnp_484 ( cddip2_out_im_status[11:0], 
	_zy_simnet_cddip2_out_im_status_543_w$[0:11]);
ixc_assign_2 _zz_strnp_483 ( im_available_kme_cddip2[1:0], 
	_zy_simnet_im_available_kme_cddip2_542_w$[0:1]);
ixc_assign _zz_strnp_482 ( cddip2_im_rdy, _zy_simnet_cddip2_im_rdy_541_w$);
ixc_assign _zz_strnp_481 ( cddip2_ism_mbe, _zy_simnet_cddip2_ism_mbe_540_w$);
ixc_assign _zz_strnp_480 ( cddip3_ism_isync, 
	_zy_simnet_cddip3_ism_isync_539_w$);
ixc_assign _zz_strnp_479 ( cddip3_ism_idat, _zy_simnet_cddip3_ism_idat_538_w$);
ixc_assign_96 _zz_strnp_478 ( cddip2_out_ia_rdata[95:0], 
	_zy_simnet_cddip2_out_ia_rdata_537_w$[0:95]);
ixc_assign_4 _zz_strnp_477 ( cddip2_out_ia_capability[19:16], 
	_zy_simnet_cddip2_out_ia_capability_536_w$[0:3]);
ixc_assign_16 _zz_strnp_476 ( cddip2_out_ia_capability[15:0], 
	_zy_simnet_cddip2_out_ia_capability_535_w$[0:15]);
ixc_assign_9 _zz_strnp_475 ( cddip2_out_ia_status[8:0], 
	_zy_simnet_cddip2_out_ia_status_534_w$[0:8]);
ixc_assign_5 _zz_strnp_474 ( cddip2_out_ia_status[13:9], 
	_zy_simnet_cddip2_out_ia_status_533_w$[0:4]);
ixc_assign_3 _zz_strnp_473 ( cddip2_out_ia_status[16:14], 
	_zy_simnet_cddip2_out_ia_status_532_w$[0:2]);
ixc_assign_12 _zz_strnp_472 ( _zy_simnet_cddip1_out_im_config_531_w$[0:11], 
	cddip1_out_im_config[11:0]);
ixc_assign_2 _zz_strnp_471 ( _zy_simnet_im_consumed_kme_cddip1_530_w$[0:1], 
	im_consumed_kme_cddip1[1:0]);
ixc_assign _zz_strnp_470 ( _zy_simnet_cddip1_im_vld_529_w$, cddip1_im_vld);
ixc_assign_96 _zz_strnp_469 ( _zy_simnet_cddip1_im_din_528_w$[0:95], { 
	cddip1_im_din[95], cddip1_im_din[94], cddip1_im_din[93], 
	cddip1_im_din[92], cddip1_im_din[91], cddip1_im_din[90], 
	cddip1_im_din[89], cddip1_im_din[88], cddip1_im_din[87], 
	cddip1_im_din[86], cddip1_im_din[85], cddip1_im_din[84], 
	cddip1_im_din[83], cddip1_im_din[82], cddip1_im_din[81], 
	cddip1_im_din[80], cddip1_im_din[79], cddip1_im_din[78], 
	cddip1_im_din[77], cddip1_im_din[76], cddip1_im_din[75], 
	cddip1_im_din[74], cddip1_im_din[73], cddip1_im_din[72], 
	cddip1_im_din[71], cddip1_im_din[70], cddip1_im_din[69], 
	cddip1_im_din[68], cddip1_im_din[67], cddip1_im_din[66], 
	cddip1_im_din[65], cddip1_im_din[64], cddip1_im_din[63], 
	cddip1_im_din[62], cddip1_im_din[61], cddip1_im_din[60], 
	cddip1_im_din[59], cddip1_im_din[58], cddip1_im_din[57], 
	cddip1_im_din[56], cddip1_im_din[55], cddip1_im_din[54], 
	cddip1_im_din[53], cddip1_im_din[52], cddip1_im_din[51], 
	cddip1_im_din[50], cddip1_im_din[49], cddip1_im_din[48], 
	cddip1_im_din[47], cddip1_im_din[46], cddip1_im_din[45], 
	cddip1_im_din[44], cddip1_im_din[43], cddip1_im_din[42], 
	cddip1_im_din[41], cddip1_im_din[40], cddip1_im_din[39], 
	cddip1_im_din[38], cddip1_im_din[37], cddip1_im_din[36], 
	cddip1_im_din[35], cddip1_im_din[34], cddip1_im_din[33], 
	cddip1_im_din[32], kme_cddip1_ob_out_pre[65], cddip1_im_din[30], 
	cddip1_im_din[29], cddip1_im_din[28], cddip1_im_din[27], 
	cddip1_im_din[26], cddip1_im_din[25], cddip1_im_din[24], 
	cddip1_im_din[23], cddip1_im_din[22], cddip1_im_din[21], 
	cddip1_im_din[20], cddip1_im_din[19], cddip1_im_din[18], 
	cddip1_im_din[17], cddip1_im_din[16], cddip1_im_din[15], 
	cddip1_im_din[14], cddip1_im_din[13], cddip1_im_din[12], 
	cddip1_im_din[11], cddip1_im_din[10], cddip1_im_din[9], 
	cddip1_im_din[8], kme_cddip1_ob_out_pre[65], cddip1_im_din[6], 
	cddip1_im_din[5], cddip1_im_din[4], cddip1_im_din[3], 
	cddip1_im_din[2], cddip1_im_din[1], cddip1_im_din[0]});
ixc_assign _zz_strnp_468 ( _zy_simnet_cddip1_ism_idat_527_w$, cddip1_ism_idat);
ixc_assign _zz_strnp_467 ( _zy_simnet_cddip1_ism_isync_526_w$, 
	cddip1_ism_isync);
ixc_assign_96 _zz_strnp_466 ( _zy_simnet_cddip1_out_ia_wdata_524_w$[0:95], 
	cddip1_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_465 ( _zy_simnet_wr_stb_523_w$, wr_stb);
ixc_assign_9 _zz_strnp_464 ( _zy_simnet_cddip1_out_ia_config_522_w$[0:8], 
	cddip1_out_ia_config[8:0]);
ixc_assign_4 _zz_strnp_463 ( _zy_simnet_cddip1_out_ia_config_521_w$[0:3], 
	cddip1_out_ia_config[12:9]);
ixc_assign_11 _zz_strnp_462 ( _zy_simnet_reg_addr_520_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_12 _zz_strnp_461 ( cddip1_out_im_status[11:0], 
	_zy_simnet_cddip1_out_im_status_519_w$[0:11]);
ixc_assign_2 _zz_strnp_460 ( im_available_kme_cddip1[1:0], 
	_zy_simnet_im_available_kme_cddip1_518_w$[0:1]);
ixc_assign _zz_strnp_459 ( cddip1_im_rdy, _zy_simnet_cddip1_im_rdy_517_w$);
ixc_assign _zz_strnp_458 ( cddip1_ism_mbe, _zy_simnet_cddip1_ism_mbe_516_w$);
ixc_assign _zz_strnp_457 ( cddip2_ism_isync, 
	_zy_simnet_cddip2_ism_isync_515_w$);
ixc_assign _zz_strnp_456 ( cddip2_ism_idat, _zy_simnet_cddip2_ism_idat_514_w$);
ixc_assign_96 _zz_strnp_455 ( cddip1_out_ia_rdata[95:0], 
	_zy_simnet_cddip1_out_ia_rdata_513_w$[0:95]);
ixc_assign_4 _zz_strnp_454 ( cddip1_out_ia_capability[19:16], 
	_zy_simnet_cddip1_out_ia_capability_512_w$[0:3]);
ixc_assign_16 _zz_strnp_453 ( cddip1_out_ia_capability[15:0], 
	_zy_simnet_cddip1_out_ia_capability_511_w$[0:15]);
ixc_assign_9 _zz_strnp_452 ( cddip1_out_ia_status[8:0], 
	_zy_simnet_cddip1_out_ia_status_510_w$[0:8]);
ixc_assign_5 _zz_strnp_451 ( cddip1_out_ia_status[13:9], 
	_zy_simnet_cddip1_out_ia_status_509_w$[0:4]);
ixc_assign_3 _zz_strnp_450 ( cddip1_out_ia_status[16:14], 
	_zy_simnet_cddip1_out_ia_status_508_w$[0:2]);
ixc_assign_12 _zz_strnp_449 ( _zy_simnet_cddip0_out_im_config_507_w$[0:11], 
	cddip0_out_im_config[11:0]);
ixc_assign_2 _zz_strnp_448 ( _zy_simnet_im_consumed_kme_cddip0_506_w$[0:1], 
	im_consumed_kme_cddip0[1:0]);
ixc_assign _zz_strnp_447 ( _zy_simnet_cddip0_im_vld_505_w$, cddip0_im_vld);
ixc_assign_96 _zz_strnp_446 ( _zy_simnet_cddip0_im_din_504_w$[0:95], { 
	cddip0_im_din[95], cddip0_im_din[94], cddip0_im_din[93], 
	cddip0_im_din[92], cddip0_im_din[91], cddip0_im_din[90], 
	cddip0_im_din[89], cddip0_im_din[88], cddip0_im_din[87], 
	cddip0_im_din[86], cddip0_im_din[85], cddip0_im_din[84], 
	cddip0_im_din[83], cddip0_im_din[82], cddip0_im_din[81], 
	cddip0_im_din[80], cddip0_im_din[79], cddip0_im_din[78], 
	cddip0_im_din[77], cddip0_im_din[76], cddip0_im_din[75], 
	cddip0_im_din[74], cddip0_im_din[73], cddip0_im_din[72], 
	cddip0_im_din[71], cddip0_im_din[70], cddip0_im_din[69], 
	cddip0_im_din[68], cddip0_im_din[67], cddip0_im_din[66], 
	cddip0_im_din[65], cddip0_im_din[64], cddip0_im_din[63], 
	cddip0_im_din[62], cddip0_im_din[61], cddip0_im_din[60], 
	cddip0_im_din[59], cddip0_im_din[58], cddip0_im_din[57], 
	cddip0_im_din[56], cddip0_im_din[55], cddip0_im_din[54], 
	cddip0_im_din[53], cddip0_im_din[52], cddip0_im_din[51], 
	cddip0_im_din[50], cddip0_im_din[49], cddip0_im_din[48], 
	cddip0_im_din[47], cddip0_im_din[46], cddip0_im_din[45], 
	cddip0_im_din[44], cddip0_im_din[43], cddip0_im_din[42], 
	cddip0_im_din[41], cddip0_im_din[40], cddip0_im_din[39], 
	cddip0_im_din[38], cddip0_im_din[37], cddip0_im_din[36], 
	cddip0_im_din[35], cddip0_im_din[34], cddip0_im_din[33], 
	cddip0_im_din[32], kme_cddip0_ob_out_pre[65], cddip0_im_din[30], 
	cddip0_im_din[29], cddip0_im_din[28], cddip0_im_din[27], 
	cddip0_im_din[26], cddip0_im_din[25], cddip0_im_din[24], 
	cddip0_im_din[23], cddip0_im_din[22], cddip0_im_din[21], 
	cddip0_im_din[20], cddip0_im_din[19], cddip0_im_din[18], 
	cddip0_im_din[17], cddip0_im_din[16], cddip0_im_din[15], 
	cddip0_im_din[14], cddip0_im_din[13], cddip0_im_din[12], 
	cddip0_im_din[11], cddip0_im_din[10], cddip0_im_din[9], 
	cddip0_im_din[8], kme_cddip0_ob_out_pre[65], cddip0_im_din[6], 
	cddip0_im_din[5], cddip0_im_din[4], cddip0_im_din[3], 
	cddip0_im_din[2], cddip0_im_din[1], cddip0_im_din[0]});
ixc_assign _zz_strnp_445 ( _zy_simnet_cddip0_ism_idat_503_w$, cddip0_ism_idat);
ixc_assign _zz_strnp_444 ( _zy_simnet_cddip0_ism_isync_502_w$, 
	cddip0_ism_isync);
ixc_assign_96 _zz_strnp_443 ( _zy_simnet_cddip0_out_ia_wdata_500_w$[0:95], 
	cddip0_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_442 ( _zy_simnet_wr_stb_499_w$, wr_stb);
ixc_assign_9 _zz_strnp_441 ( _zy_simnet_cddip0_out_ia_config_498_w$[0:8], 
	cddip0_out_ia_config[8:0]);
ixc_assign_4 _zz_strnp_440 ( _zy_simnet_cddip0_out_ia_config_497_w$[0:3], 
	cddip0_out_ia_config[12:9]);
ixc_assign_11 _zz_strnp_439 ( _zy_simnet_reg_addr_496_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_12 _zz_strnp_438 ( cddip0_out_im_status[11:0], 
	_zy_simnet_cddip0_out_im_status_495_w$[0:11]);
ixc_assign_2 _zz_strnp_437 ( im_available_kme_cddip0[1:0], 
	_zy_simnet_im_available_kme_cddip0_494_w$[0:1]);
ixc_assign _zz_strnp_436 ( cddip0_im_rdy, _zy_simnet_cddip0_im_rdy_493_w$);
ixc_assign _zz_strnp_435 ( cddip0_ism_mbe, _zy_simnet_cddip0_ism_mbe_492_w$);
ixc_assign _zz_strnp_434 ( cddip1_ism_isync, 
	_zy_simnet_cddip1_ism_isync_491_w$);
ixc_assign _zz_strnp_433 ( cddip1_ism_idat, _zy_simnet_cddip1_ism_idat_490_w$);
ixc_assign_96 _zz_strnp_432 ( cddip0_out_ia_rdata[95:0], 
	_zy_simnet_cddip0_out_ia_rdata_489_w$[0:95]);
ixc_assign_4 _zz_strnp_431 ( cddip0_out_ia_capability[19:16], 
	_zy_simnet_cddip0_out_ia_capability_488_w$[0:3]);
ixc_assign_16 _zz_strnp_430 ( cddip0_out_ia_capability[15:0], 
	_zy_simnet_cddip0_out_ia_capability_487_w$[0:15]);
ixc_assign_9 _zz_strnp_429 ( cddip0_out_ia_status[8:0], 
	_zy_simnet_cddip0_out_ia_status_486_w$[0:8]);
ixc_assign_5 _zz_strnp_428 ( cddip0_out_ia_status[13:9], 
	_zy_simnet_cddip0_out_ia_status_485_w$[0:4]);
ixc_assign_3 _zz_strnp_427 ( cddip0_out_ia_status[16:14], 
	_zy_simnet_cddip0_out_ia_status_484_w$[0:2]);
ixc_assign_12 _zz_strnp_426 ( _zy_simnet_cceip3_out_im_config_483_w$[0:11], 
	cceip3_out_im_config[11:0]);
ixc_assign_2 _zz_strnp_425 ( _zy_simnet_im_consumed_kme_cceip3_482_w$[0:1], 
	im_consumed_kme_cceip3[1:0]);
ixc_assign _zz_strnp_424 ( _zy_simnet_cceip3_im_vld_481_w$, cceip3_im_vld);
ixc_assign_96 _zz_strnp_423 ( _zy_simnet_cceip3_im_din_480_w$[0:95], { 
	cceip3_im_din[95], cceip3_im_din[94], cceip3_im_din[93], 
	cceip3_im_din[92], cceip3_im_din[91], cceip3_im_din[90], 
	cceip3_im_din[89], cceip3_im_din[88], cceip3_im_din[87], 
	cceip3_im_din[86], cceip3_im_din[85], cceip3_im_din[84], 
	cceip3_im_din[83], cceip3_im_din[82], cceip3_im_din[81], 
	cceip3_im_din[80], cceip3_im_din[79], cceip3_im_din[78], 
	cceip3_im_din[77], cceip3_im_din[76], cceip3_im_din[75], 
	cceip3_im_din[74], cceip3_im_din[73], cceip3_im_din[72], 
	cceip3_im_din[71], cceip3_im_din[70], cceip3_im_din[69], 
	cceip3_im_din[68], cceip3_im_din[67], cceip3_im_din[66], 
	cceip3_im_din[65], cceip3_im_din[64], cceip3_im_din[63], 
	cceip3_im_din[62], cceip3_im_din[61], cceip3_im_din[60], 
	cceip3_im_din[59], cceip3_im_din[58], cceip3_im_din[57], 
	cceip3_im_din[56], cceip3_im_din[55], cceip3_im_din[54], 
	cceip3_im_din[53], cceip3_im_din[52], cceip3_im_din[51], 
	cceip3_im_din[50], cceip3_im_din[49], cceip3_im_din[48], 
	cceip3_im_din[47], cceip3_im_din[46], cceip3_im_din[45], 
	cceip3_im_din[44], cceip3_im_din[43], cceip3_im_din[42], 
	cceip3_im_din[41], cceip3_im_din[40], cceip3_im_din[39], 
	cceip3_im_din[38], cceip3_im_din[37], cceip3_im_din[36], 
	cceip3_im_din[35], cceip3_im_din[34], cceip3_im_din[33], 
	cceip3_im_din[32], kme_cceip3_ob_out_pre[65], cceip3_im_din[30], 
	cceip3_im_din[29], cceip3_im_din[28], cceip3_im_din[27], 
	cceip3_im_din[26], cceip3_im_din[25], cceip3_im_din[24], 
	cceip3_im_din[23], cceip3_im_din[22], cceip3_im_din[21], 
	cceip3_im_din[20], cceip3_im_din[19], cceip3_im_din[18], 
	cceip3_im_din[17], cceip3_im_din[16], cceip3_im_din[15], 
	cceip3_im_din[14], cceip3_im_din[13], cceip3_im_din[12], 
	cceip3_im_din[11], cceip3_im_din[10], cceip3_im_din[9], 
	cceip3_im_din[8], kme_cceip3_ob_out_pre[65], cceip3_im_din[6], 
	cceip3_im_din[5], cceip3_im_din[4], cceip3_im_din[3], 
	cceip3_im_din[2], cceip3_im_din[1], cceip3_im_din[0]});
ixc_assign _zz_strnp_422 ( _zy_simnet_cceip3_ism_idat_479_w$, cceip3_ism_idat);
ixc_assign _zz_strnp_421 ( _zy_simnet_cceip3_ism_isync_478_w$, 
	cceip3_ism_isync);
ixc_assign_96 _zz_strnp_420 ( _zy_simnet_cceip3_out_ia_wdata_476_w$[0:95], 
	cceip3_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_419 ( _zy_simnet_wr_stb_475_w$, wr_stb);
ixc_assign_9 _zz_strnp_418 ( _zy_simnet_cceip3_out_ia_config_474_w$[0:8], 
	cceip3_out_ia_config[8:0]);
ixc_assign_4 _zz_strnp_417 ( _zy_simnet_cceip3_out_ia_config_473_w$[0:3], 
	cceip3_out_ia_config[12:9]);
ixc_assign_11 _zz_strnp_416 ( _zy_simnet_reg_addr_472_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_12 _zz_strnp_415 ( cceip3_out_im_status[11:0], 
	_zy_simnet_cceip3_out_im_status_471_w$[0:11]);
ixc_assign_2 _zz_strnp_414 ( im_available_kme_cceip3[1:0], 
	_zy_simnet_im_available_kme_cceip3_470_w$[0:1]);
ixc_assign _zz_strnp_413 ( cceip3_im_rdy, _zy_simnet_cceip3_im_rdy_469_w$);
ixc_assign _zz_strnp_412 ( cceip3_ism_mbe, _zy_simnet_cceip3_ism_mbe_468_w$);
ixc_assign _zz_strnp_411 ( cddip0_ism_isync, 
	_zy_simnet_cddip0_ism_isync_467_w$);
ixc_assign _zz_strnp_410 ( cddip0_ism_idat, _zy_simnet_cddip0_ism_idat_466_w$);
ixc_assign_96 _zz_strnp_409 ( cceip3_out_ia_rdata[95:0], 
	_zy_simnet_cceip3_out_ia_rdata_465_w$[0:95]);
ixc_assign_4 _zz_strnp_408 ( cceip3_out_ia_capability[19:16], 
	_zy_simnet_cceip3_out_ia_capability_464_w$[0:3]);
ixc_assign_16 _zz_strnp_407 ( cceip3_out_ia_capability[15:0], 
	_zy_simnet_cceip3_out_ia_capability_463_w$[0:15]);
ixc_assign_9 _zz_strnp_406 ( cceip3_out_ia_status[8:0], 
	_zy_simnet_cceip3_out_ia_status_462_w$[0:8]);
ixc_assign_5 _zz_strnp_405 ( cceip3_out_ia_status[13:9], 
	_zy_simnet_cceip3_out_ia_status_461_w$[0:4]);
ixc_assign_3 _zz_strnp_404 ( cceip3_out_ia_status[16:14], 
	_zy_simnet_cceip3_out_ia_status_460_w$[0:2]);
ixc_assign_12 _zz_strnp_403 ( _zy_simnet_cceip2_out_im_config_459_w$[0:11], 
	cceip2_out_im_config[11:0]);
ixc_assign_2 _zz_strnp_402 ( _zy_simnet_im_consumed_kme_cceip2_458_w$[0:1], 
	im_consumed_kme_cceip2[1:0]);
ixc_assign _zz_strnp_401 ( _zy_simnet_cceip2_im_vld_457_w$, cceip2_im_vld);
ixc_assign_96 _zz_strnp_400 ( _zy_simnet_cceip2_im_din_456_w$[0:95], { 
	cceip2_im_din[95], cceip2_im_din[94], cceip2_im_din[93], 
	cceip2_im_din[92], cceip2_im_din[91], cceip2_im_din[90], 
	cceip2_im_din[89], cceip2_im_din[88], cceip2_im_din[87], 
	cceip2_im_din[86], cceip2_im_din[85], cceip2_im_din[84], 
	cceip2_im_din[83], cceip2_im_din[82], cceip2_im_din[81], 
	cceip2_im_din[80], cceip2_im_din[79], cceip2_im_din[78], 
	cceip2_im_din[77], cceip2_im_din[76], cceip2_im_din[75], 
	cceip2_im_din[74], cceip2_im_din[73], cceip2_im_din[72], 
	cceip2_im_din[71], cceip2_im_din[70], cceip2_im_din[69], 
	cceip2_im_din[68], cceip2_im_din[67], cceip2_im_din[66], 
	cceip2_im_din[65], cceip2_im_din[64], cceip2_im_din[63], 
	cceip2_im_din[62], cceip2_im_din[61], cceip2_im_din[60], 
	cceip2_im_din[59], cceip2_im_din[58], cceip2_im_din[57], 
	cceip2_im_din[56], cceip2_im_din[55], cceip2_im_din[54], 
	cceip2_im_din[53], cceip2_im_din[52], cceip2_im_din[51], 
	cceip2_im_din[50], cceip2_im_din[49], cceip2_im_din[48], 
	cceip2_im_din[47], cceip2_im_din[46], cceip2_im_din[45], 
	cceip2_im_din[44], cceip2_im_din[43], cceip2_im_din[42], 
	cceip2_im_din[41], cceip2_im_din[40], cceip2_im_din[39], 
	cceip2_im_din[38], cceip2_im_din[37], cceip2_im_din[36], 
	cceip2_im_din[35], cceip2_im_din[34], cceip2_im_din[33], 
	cceip2_im_din[32], kme_cceip2_ob_out_pre[65], cceip2_im_din[30], 
	cceip2_im_din[29], cceip2_im_din[28], cceip2_im_din[27], 
	cceip2_im_din[26], cceip2_im_din[25], cceip2_im_din[24], 
	cceip2_im_din[23], cceip2_im_din[22], cceip2_im_din[21], 
	cceip2_im_din[20], cceip2_im_din[19], cceip2_im_din[18], 
	cceip2_im_din[17], cceip2_im_din[16], cceip2_im_din[15], 
	cceip2_im_din[14], cceip2_im_din[13], cceip2_im_din[12], 
	cceip2_im_din[11], cceip2_im_din[10], cceip2_im_din[9], 
	cceip2_im_din[8], kme_cceip2_ob_out_pre[65], cceip2_im_din[6], 
	cceip2_im_din[5], cceip2_im_din[4], cceip2_im_din[3], 
	cceip2_im_din[2], cceip2_im_din[1], cceip2_im_din[0]});
ixc_assign _zz_strnp_399 ( _zy_simnet_cceip2_ism_idat_455_w$, cceip2_ism_idat);
ixc_assign _zz_strnp_398 ( _zy_simnet_cceip2_ism_isync_454_w$, 
	cceip2_ism_isync);
ixc_assign_96 _zz_strnp_397 ( _zy_simnet_cceip2_out_ia_wdata_452_w$[0:95], 
	cceip2_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_396 ( _zy_simnet_wr_stb_451_w$, wr_stb);
ixc_assign_9 _zz_strnp_395 ( _zy_simnet_cceip2_out_ia_config_450_w$[0:8], 
	cceip2_out_ia_config[8:0]);
ixc_assign_4 _zz_strnp_394 ( _zy_simnet_cceip2_out_ia_config_449_w$[0:3], 
	cceip2_out_ia_config[12:9]);
ixc_assign_11 _zz_strnp_393 ( _zy_simnet_reg_addr_448_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_12 _zz_strnp_392 ( cceip2_out_im_status[11:0], 
	_zy_simnet_cceip2_out_im_status_447_w$[0:11]);
ixc_assign_2 _zz_strnp_391 ( im_available_kme_cceip2[1:0], 
	_zy_simnet_im_available_kme_cceip2_446_w$[0:1]);
ixc_assign _zz_strnp_390 ( cceip2_im_rdy, _zy_simnet_cceip2_im_rdy_445_w$);
ixc_assign _zz_strnp_389 ( cceip2_ism_mbe, _zy_simnet_cceip2_ism_mbe_444_w$);
ixc_assign _zz_strnp_388 ( cceip3_ism_isync, 
	_zy_simnet_cceip3_ism_isync_443_w$);
ixc_assign _zz_strnp_387 ( cceip3_ism_idat, _zy_simnet_cceip3_ism_idat_442_w$);
ixc_assign_96 _zz_strnp_386 ( cceip2_out_ia_rdata[95:0], 
	_zy_simnet_cceip2_out_ia_rdata_441_w$[0:95]);
ixc_assign_4 _zz_strnp_385 ( cceip2_out_ia_capability[19:16], 
	_zy_simnet_cceip2_out_ia_capability_440_w$[0:3]);
ixc_assign_16 _zz_strnp_384 ( cceip2_out_ia_capability[15:0], 
	_zy_simnet_cceip2_out_ia_capability_439_w$[0:15]);
ixc_assign_9 _zz_strnp_383 ( cceip2_out_ia_status[8:0], 
	_zy_simnet_cceip2_out_ia_status_438_w$[0:8]);
ixc_assign_5 _zz_strnp_382 ( cceip2_out_ia_status[13:9], 
	_zy_simnet_cceip2_out_ia_status_437_w$[0:4]);
ixc_assign_3 _zz_strnp_381 ( cceip2_out_ia_status[16:14], 
	_zy_simnet_cceip2_out_ia_status_436_w$[0:2]);
ixc_assign_12 _zz_strnp_380 ( _zy_simnet_cceip1_out_im_config_435_w$[0:11], 
	cceip1_out_im_config[11:0]);
ixc_assign_2 _zz_strnp_379 ( _zy_simnet_im_consumed_kme_cceip1_434_w$[0:1], 
	im_consumed_kme_cceip1[1:0]);
ixc_assign _zz_strnp_378 ( _zy_simnet_cceip1_im_vld_433_w$, cceip1_im_vld);
ixc_assign_96 _zz_strnp_377 ( _zy_simnet_cceip1_im_din_432_w$[0:95], { 
	cceip1_im_din[95], cceip1_im_din[94], cceip1_im_din[93], 
	cceip1_im_din[92], cceip1_im_din[91], cceip1_im_din[90], 
	cceip1_im_din[89], cceip1_im_din[88], cceip1_im_din[87], 
	cceip1_im_din[86], cceip1_im_din[85], cceip1_im_din[84], 
	cceip1_im_din[83], cceip1_im_din[82], cceip1_im_din[81], 
	cceip1_im_din[80], cceip1_im_din[79], cceip1_im_din[78], 
	cceip1_im_din[77], cceip1_im_din[76], cceip1_im_din[75], 
	cceip1_im_din[74], cceip1_im_din[73], cceip1_im_din[72], 
	cceip1_im_din[71], cceip1_im_din[70], cceip1_im_din[69], 
	cceip1_im_din[68], cceip1_im_din[67], cceip1_im_din[66], 
	cceip1_im_din[65], cceip1_im_din[64], cceip1_im_din[63], 
	cceip1_im_din[62], cceip1_im_din[61], cceip1_im_din[60], 
	cceip1_im_din[59], cceip1_im_din[58], cceip1_im_din[57], 
	cceip1_im_din[56], cceip1_im_din[55], cceip1_im_din[54], 
	cceip1_im_din[53], cceip1_im_din[52], cceip1_im_din[51], 
	cceip1_im_din[50], cceip1_im_din[49], cceip1_im_din[48], 
	cceip1_im_din[47], cceip1_im_din[46], cceip1_im_din[45], 
	cceip1_im_din[44], cceip1_im_din[43], cceip1_im_din[42], 
	cceip1_im_din[41], cceip1_im_din[40], cceip1_im_din[39], 
	cceip1_im_din[38], cceip1_im_din[37], cceip1_im_din[36], 
	cceip1_im_din[35], cceip1_im_din[34], cceip1_im_din[33], 
	cceip1_im_din[32], kme_cceip1_ob_out_pre[65], cceip1_im_din[30], 
	cceip1_im_din[29], cceip1_im_din[28], cceip1_im_din[27], 
	cceip1_im_din[26], cceip1_im_din[25], cceip1_im_din[24], 
	cceip1_im_din[23], cceip1_im_din[22], cceip1_im_din[21], 
	cceip1_im_din[20], cceip1_im_din[19], cceip1_im_din[18], 
	cceip1_im_din[17], cceip1_im_din[16], cceip1_im_din[15], 
	cceip1_im_din[14], cceip1_im_din[13], cceip1_im_din[12], 
	cceip1_im_din[11], cceip1_im_din[10], cceip1_im_din[9], 
	cceip1_im_din[8], kme_cceip1_ob_out_pre[65], cceip1_im_din[6], 
	cceip1_im_din[5], cceip1_im_din[4], cceip1_im_din[3], 
	cceip1_im_din[2], cceip1_im_din[1], cceip1_im_din[0]});
ixc_assign _zz_strnp_376 ( _zy_simnet_cceip1_ism_idat_431_w$, cceip1_ism_idat);
ixc_assign _zz_strnp_375 ( _zy_simnet_cceip1_ism_isync_430_w$, 
	cceip1_ism_isync);
ixc_assign_96 _zz_strnp_374 ( _zy_simnet_cceip1_out_ia_wdata_428_w$[0:95], 
	cceip1_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_373 ( _zy_simnet_wr_stb_427_w$, wr_stb);
ixc_assign_9 _zz_strnp_372 ( _zy_simnet_cceip1_out_ia_config_426_w$[0:8], 
	cceip1_out_ia_config[8:0]);
ixc_assign_4 _zz_strnp_371 ( _zy_simnet_cceip1_out_ia_config_425_w$[0:3], 
	cceip1_out_ia_config[12:9]);
ixc_assign_11 _zz_strnp_370 ( _zy_simnet_reg_addr_424_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_12 _zz_strnp_369 ( cceip1_out_im_status[11:0], 
	_zy_simnet_cceip1_out_im_status_423_w$[0:11]);
ixc_assign_2 _zz_strnp_368 ( im_available_kme_cceip1[1:0], 
	_zy_simnet_im_available_kme_cceip1_422_w$[0:1]);
ixc_assign _zz_strnp_367 ( cceip1_im_rdy, _zy_simnet_cceip1_im_rdy_421_w$);
ixc_assign _zz_strnp_366 ( cceip1_ism_mbe, _zy_simnet_cceip1_ism_mbe_420_w$);
ixc_assign _zz_strnp_365 ( cceip2_ism_isync, 
	_zy_simnet_cceip2_ism_isync_419_w$);
ixc_assign _zz_strnp_364 ( cceip2_ism_idat, _zy_simnet_cceip2_ism_idat_418_w$);
ixc_assign_96 _zz_strnp_363 ( cceip1_out_ia_rdata[95:0], 
	_zy_simnet_cceip1_out_ia_rdata_417_w$[0:95]);
ixc_assign_4 _zz_strnp_362 ( cceip1_out_ia_capability[19:16], 
	_zy_simnet_cceip1_out_ia_capability_416_w$[0:3]);
ixc_assign_16 _zz_strnp_361 ( cceip1_out_ia_capability[15:0], 
	_zy_simnet_cceip1_out_ia_capability_415_w$[0:15]);
ixc_assign_9 _zz_strnp_360 ( cceip1_out_ia_status[8:0], 
	_zy_simnet_cceip1_out_ia_status_414_w$[0:8]);
ixc_assign_5 _zz_strnp_359 ( cceip1_out_ia_status[13:9], 
	_zy_simnet_cceip1_out_ia_status_413_w$[0:4]);
ixc_assign_3 _zz_strnp_358 ( cceip1_out_ia_status[16:14], 
	_zy_simnet_cceip1_out_ia_status_412_w$[0:2]);
ixc_assign_12 _zz_strnp_357 ( _zy_simnet_cceip0_out_im_config_411_w$[0:11], 
	cceip0_out_im_config[11:0]);
ixc_assign_2 _zz_strnp_356 ( _zy_simnet_im_consumed_kme_cceip0_410_w$[0:1], 
	im_consumed_kme_cceip0[1:0]);
ixc_assign _zz_strnp_355 ( _zy_simnet_cceip0_im_vld_409_w$, cceip0_im_vld);
ixc_assign_96 _zz_strnp_354 ( _zy_simnet_cceip0_im_din_408_w$[0:95], { 
	cceip0_im_din[95], cceip0_im_din[94], cceip0_im_din[93], 
	cceip0_im_din[92], cceip0_im_din[91], cceip0_im_din[90], 
	cceip0_im_din[89], cceip0_im_din[88], cceip0_im_din[87], 
	cceip0_im_din[86], cceip0_im_din[85], cceip0_im_din[84], 
	cceip0_im_din[83], cceip0_im_din[82], cceip0_im_din[81], 
	cceip0_im_din[80], cceip0_im_din[79], cceip0_im_din[78], 
	cceip0_im_din[77], cceip0_im_din[76], cceip0_im_din[75], 
	cceip0_im_din[74], cceip0_im_din[73], cceip0_im_din[72], 
	cceip0_im_din[71], cceip0_im_din[70], cceip0_im_din[69], 
	cceip0_im_din[68], cceip0_im_din[67], cceip0_im_din[66], 
	cceip0_im_din[65], cceip0_im_din[64], cceip0_im_din[63], 
	cceip0_im_din[62], cceip0_im_din[61], cceip0_im_din[60], 
	cceip0_im_din[59], cceip0_im_din[58], cceip0_im_din[57], 
	cceip0_im_din[56], cceip0_im_din[55], cceip0_im_din[54], 
	cceip0_im_din[53], cceip0_im_din[52], cceip0_im_din[51], 
	cceip0_im_din[50], cceip0_im_din[49], cceip0_im_din[48], 
	cceip0_im_din[47], cceip0_im_din[46], cceip0_im_din[45], 
	cceip0_im_din[44], cceip0_im_din[43], cceip0_im_din[42], 
	cceip0_im_din[41], cceip0_im_din[40], cceip0_im_din[39], 
	cceip0_im_din[38], cceip0_im_din[37], cceip0_im_din[36], 
	cceip0_im_din[35], cceip0_im_din[34], cceip0_im_din[33], 
	cceip0_im_din[32], kme_cceip0_ob_out_pre[65], cceip0_im_din[30], 
	cceip0_im_din[29], cceip0_im_din[28], cceip0_im_din[27], 
	cceip0_im_din[26], cceip0_im_din[25], cceip0_im_din[24], 
	cceip0_im_din[23], cceip0_im_din[22], cceip0_im_din[21], 
	cceip0_im_din[20], cceip0_im_din[19], cceip0_im_din[18], 
	cceip0_im_din[17], cceip0_im_din[16], cceip0_im_din[15], 
	cceip0_im_din[14], cceip0_im_din[13], cceip0_im_din[12], 
	cceip0_im_din[11], cceip0_im_din[10], cceip0_im_din[9], 
	cceip0_im_din[8], kme_cceip0_ob_out_pre[65], cceip0_im_din[6], 
	cceip0_im_din[5], cceip0_im_din[4], cceip0_im_din[3], 
	cceip0_im_din[2], cceip0_im_din[1], cceip0_im_din[0]});
ixc_assign _zz_strnp_353 ( _zy_simnet_cceip0_ism_bimc_idat_407_w$, 
	cceip0_ism_bimc_idat);
ixc_assign _zz_strnp_352 ( _zy_simnet_cceip0_ism_bimc_isync_406_w$, 
	cceip0_ism_bimc_isync);
ixc_assign_96 _zz_strnp_351 ( _zy_simnet_cceip0_out_ia_wdata_404_w$[0:95], 
	cceip0_out_ia_wdata[95:0]);
ixc_assign _zz_strnp_350 ( _zy_simnet_wr_stb_403_w$, wr_stb);
ixc_assign_9 _zz_strnp_349 ( _zy_simnet_cceip0_out_ia_config_402_w$[0:8], 
	cceip0_out_ia_config[8:0]);
ixc_assign_4 _zz_strnp_348 ( _zy_simnet_cceip0_out_ia_config_401_w$[0:3], 
	cceip0_out_ia_config[12:9]);
ixc_assign_11 _zz_strnp_347 ( _zy_simnet_reg_addr_400_w$[0:10], 
	reg_addr[10:0]);
ixc_assign_12 _zz_strnp_346 ( cceip0_out_im_status[11:0], 
	_zy_simnet_cceip0_out_im_status_399_w$[0:11]);
ixc_assign_2 _zz_strnp_345 ( im_available_kme_cceip0[1:0], 
	_zy_simnet_im_available_kme_cceip0_398_w$[0:1]);
ixc_assign _zz_strnp_344 ( cceip0_im_rdy, _zy_simnet_cceip0_im_rdy_397_w$);
ixc_assign _zz_strnp_343 ( cceip0_ism_mbe, _zy_simnet_cceip0_ism_mbe_396_w$);
ixc_assign _zz_strnp_342 ( cceip1_ism_isync, 
	_zy_simnet_cceip1_ism_isync_395_w$);
ixc_assign _zz_strnp_341 ( cceip1_ism_idat, _zy_simnet_cceip1_ism_idat_394_w$);
ixc_assign_96 _zz_strnp_340 ( cceip0_out_ia_rdata[95:0], 
	_zy_simnet_cceip0_out_ia_rdata_393_w$[0:95]);
ixc_assign_4 _zz_strnp_339 ( cceip0_out_ia_capability[19:16], 
	_zy_simnet_cceip0_out_ia_capability_392_w$[0:3]);
ixc_assign_16 _zz_strnp_338 ( cceip0_out_ia_capability[15:0], 
	_zy_simnet_cceip0_out_ia_capability_391_w$[0:15]);
ixc_assign_9 _zz_strnp_337 ( cceip0_out_ia_status[8:0], 
	_zy_simnet_cceip0_out_ia_status_390_w$[0:8]);
ixc_assign_5 _zz_strnp_336 ( cceip0_out_ia_status[13:9], 
	_zy_simnet_cceip0_out_ia_status_389_w$[0:4]);
ixc_assign_3 _zz_strnp_335 ( cceip0_out_ia_status[16:14], 
	_zy_simnet_cceip0_out_ia_status_388_w$[0:2]);
ixc_assign _zz_strnp_334 ( _zy_simnet_cddip3_im_rdy_387_w$, cddip3_im_rdy);
ixc_assign _zz_strnp_333 ( cddip3_im_vld, _zy_simnet_cddip3_im_vld_385_w$);
ixc_assign_83 _zz_strnp_332 ( kme_cddip3_ob_out_post[82:0], 
	_zy_simnet_kme_cddip3_ob_out_post_384_w$[0:82]);
ixc_assign _zz_strnp_331 ( kme_cddip3_ob_in_mod[0], 
	_zy_simnet_kme_cddip3_ob_in_mod_383_w$);
ixc_assign _zz_strnp_330 ( _zy_simnet_cddip2_im_rdy_382_w$, cddip2_im_rdy);
ixc_assign _zz_strnp_329 ( cddip2_im_vld, _zy_simnet_cddip2_im_vld_380_w$);
ixc_assign_83 _zz_strnp_328 ( kme_cddip2_ob_out_post[82:0], 
	_zy_simnet_kme_cddip2_ob_out_post_379_w$[0:82]);
ixc_assign _zz_strnp_327 ( kme_cddip2_ob_in_mod[0], 
	_zy_simnet_kme_cddip2_ob_in_mod_378_w$);
ixc_assign _zz_strnp_326 ( _zy_simnet_cddip1_im_rdy_377_w$, cddip1_im_rdy);
ixc_assign _zz_strnp_325 ( cddip1_im_vld, _zy_simnet_cddip1_im_vld_375_w$);
ixc_assign_83 _zz_strnp_324 ( kme_cddip1_ob_out_post[82:0], 
	_zy_simnet_kme_cddip1_ob_out_post_374_w$[0:82]);
ixc_assign _zz_strnp_323 ( kme_cddip1_ob_in_mod[0], 
	_zy_simnet_kme_cddip1_ob_in_mod_373_w$);
ixc_assign _zz_strnp_322 ( _zy_simnet_cddip0_im_rdy_372_w$, cddip0_im_rdy);
ixc_assign _zz_strnp_321 ( cddip0_im_vld, _zy_simnet_cddip0_im_vld_370_w$);
ixc_assign_83 _zz_strnp_320 ( kme_cddip0_ob_out_post[82:0], 
	_zy_simnet_kme_cddip0_ob_out_post_369_w$[0:82]);
ixc_assign _zz_strnp_319 ( kme_cddip0_ob_in_mod[0], 
	_zy_simnet_kme_cddip0_ob_in_mod_368_w$);
ixc_assign _zz_strnp_318 ( _zy_simnet_cceip3_im_rdy_367_w$, cceip3_im_rdy);
ixc_assign _zz_strnp_317 ( cceip3_im_vld, _zy_simnet_cceip3_im_vld_365_w$);
ixc_assign_83 _zz_strnp_316 ( kme_cceip3_ob_out_post[82:0], 
	_zy_simnet_kme_cceip3_ob_out_post_364_w$[0:82]);
ixc_assign _zz_strnp_315 ( kme_cceip3_ob_in_mod[0], 
	_zy_simnet_kme_cceip3_ob_in_mod_363_w$);
ixc_assign _zz_strnp_314 ( _zy_simnet_cceip2_im_rdy_362_w$, cceip2_im_rdy);
ixc_assign _zz_strnp_313 ( cceip2_im_vld, _zy_simnet_cceip2_im_vld_360_w$);
ixc_assign_83 _zz_strnp_312 ( kme_cceip2_ob_out_post[82:0], 
	_zy_simnet_kme_cceip2_ob_out_post_359_w$[0:82]);
ixc_assign _zz_strnp_311 ( kme_cceip2_ob_in_mod[0], 
	_zy_simnet_kme_cceip2_ob_in_mod_358_w$);
ixc_assign _zz_strnp_310 ( _zy_simnet_cceip1_im_rdy_357_w$, cceip1_im_rdy);
ixc_assign _zz_strnp_309 ( cceip1_im_vld, _zy_simnet_cceip1_im_vld_355_w$);
ixc_assign_83 _zz_strnp_308 ( kme_cceip1_ob_out_post[82:0], 
	_zy_simnet_kme_cceip1_ob_out_post_354_w$[0:82]);
ixc_assign _zz_strnp_307 ( kme_cceip1_ob_in_mod[0], 
	_zy_simnet_kme_cceip1_ob_in_mod_353_w$);
ixc_assign _zz_strnp_306 ( _zy_simnet_cceip0_im_rdy_352_w$, cceip0_im_rdy);
ixc_assign _zz_strnp_305 ( cceip0_im_vld, _zy_simnet_cceip0_im_vld_350_w$);
ixc_assign_83 _zz_strnp_304 ( kme_cceip0_ob_out_post[82:0], 
	_zy_simnet_kme_cceip0_ob_out_post_349_w$[0:82]);
ixc_assign _zz_strnp_303 ( kme_cceip0_ob_in_mod[0], 
	_zy_simnet_kme_cceip0_ob_in_mod_348_w$);
ixc_assign _zz_strnp_302 ( rbus_ring_o[0], _zy_simnet_rbus_ring_o_347_w$);
ixc_assign _zz_strnp_301 ( rbus_ring_o[1], _zy_simnet_rbus_ring_o_346_w$);
ixc_assign_32 _zz_strnp_300 ( rbus_ring_o[33:2], 
	_zy_simnet_rbus_ring_o_345_w$[0:31]);
ixc_assign _zz_strnp_299 ( _zy_simnet_locl_err_ack_344_w$, locl_err_ack);
ixc_assign _zz_strnp_298 ( _zy_simnet_locl_ack_343_w$, locl_ack);
ixc_assign_32 _zz_strnp_297 ( _zy_simnet_locl_rd_data_342_w$[0:31], 
	locl_rd_data[31:0]);
ixc_assign _zz_strnp_296 ( locl_rd_strb, _zy_simnet_locl_rd_strb_341_w$);
ixc_assign_32 _zz_strnp_295 ( locl_wr_data[31:0], 
	_zy_simnet_locl_wr_data_340_w$[0:31]);
ixc_assign _zz_strnp_294 ( locl_wr_strb, _zy_simnet_locl_wr_strb_339_w$);
ixc_assign_11 _zz_strnp_293 ( locl_addr[10:0], 
	_zy_simnet_locl_addr_338_w$[0:10]);
ixc_assign _zz_strnp_292 ( rbus_ring_o[34], _zy_simnet_rbus_ring_o_337_w$);
ixc_assign_32 _zz_strnp_291 ( rbus_ring_o[66:35], 
	_zy_simnet_rbus_ring_o_336_w$[0:31]);
ixc_assign _zz_strnp_290 ( rbus_ring_o[67], _zy_simnet_rbus_ring_o_335_w$);
ixc_assign_16 _zz_strnp_289 ( rbus_ring_o[83:68], 
	_zy_simnet_rbus_ring_o_334_w$[0:15]);
ixc_assign_11 _zz_strnp_288 ( reg_addr[10:0], 
	_zy_simnet_reg_addr_333_w$[0:10]);
ixc_assign_32 _zz_strnp_287 ( wr_data[31:0], _zy_simnet_wr_data_332_w$[0:31]);
ixc_assign _zz_strnp_286 ( wr_stb, _zy_simnet_wr_stb_330_w$);
ixc_assign_32 _zz_strnp_285 ( _zy_simnet_sa_ctrl_ia_rdata_329_w$[0:31], 
	sa_ctrl_ia_rdata[31:0]);
ixc_assign_13 _zz_strnp_284 ( _zy_simnet_sa_ctrl_ia_status_328_w$[0:12], 
	sa_ctrl_ia_status[12:0]);
ixc_assign_20 _zz_strnp_283 ( _zy_simnet_sa_ctrl_ia_capability_327_w$[0:19], 
	sa_ctrl_ia_capability[19:0]);
ixc_assign_32 _zz_strnp_282 ( _zy_simnet_sa_global_ctrl_326_w$[0:31], 
	sa_global_ctrl[31:0]);
ixc_assign_32 _zz_strnp_281 ( _zy_simnet_sa_count_ia_rdata_325_w$[0:31], 
	sa_count_ia_rdata[63:32]);
ixc_assign_32 _zz_strnp_280 ( _zy_simnet_sa_count_ia_rdata_324_w$[0:31], 
	sa_count_ia_rdata[31:0]);
ixc_assign_13 _zz_strnp_279 ( _zy_simnet_sa_count_ia_status_323_w$[0:12], 
	sa_count_ia_status[12:0]);
ixc_assign_20 _zz_strnp_278 ( _zy_simnet_sa_count_ia_capability_322_w$[0:19], 
	sa_count_ia_capability[19:0]);
ixc_assign_32 _zz_strnp_277 ( _zy_simnet_sa_snapshot_ia_rdata_321_w$[0:31], 
	sa_snapshot_ia_rdata[63:32]);
ixc_assign_32 _zz_strnp_276 ( _zy_simnet_sa_snapshot_ia_rdata_320_w$[0:31], 
	sa_snapshot_ia_rdata[31:0]);
ixc_assign_13 _zz_strnp_275 ( _zy_simnet_sa_snapshot_ia_status_319_w$[0:12], 
	sa_snapshot_ia_status[12:0]);
ixc_assign_20 _zz_strnp_274 ( 
	_zy_simnet_sa_snapshot_ia_capability_318_w$[0:19], 
	sa_snapshot_ia_capability[19:0]);
ixc_assign_32 _zz_strnp_273 ( _zy_simnet_regs_sa_ctrl_317_w$[0:31], 
	regs_sa_ctrl[31:0]);
ixc_assign_9 _zz_strnp_272 ( _zy_simnet_tready_override_316_w$[0:8], 
	tready_override[8:0]);
ixc_assign_16 _zz_strnp_271 ( _zy_simnet_im_available_314_w$[0:15], { 
	im_available_kme_cddip3[1], im_available_kme_cddip3[0], 
	im_available_kme_cddip2[1], im_available_kme_cddip2[0], 
	im_available_kme_cddip1[1], im_available_kme_cddip1[0], 
	im_available_kme_cddip0[1], im_available_kme_cddip0[0], 
	im_available_kme_cceip3[1], im_available_kme_cceip3[0], 
	im_available_kme_cceip2[1], im_available_kme_cceip2[0], 
	im_available_kme_cceip1[1], im_available_kme_cceip1[0], 
	im_available_kme_cceip0[1], im_available_kme_cceip0[0]});
ixc_assign_32 _zz_strnp_270 ( _zy_simnet_bimc_dbgcmd0_313_w$[0:31], 
	bimc_dbgcmd0[31:0]);
ixc_assign_32 _zz_strnp_269 ( _zy_simnet_bimc_dbgcmd1_312_w$[0:31], 
	bimc_dbgcmd1[31:0]);
ixc_assign_10 _zz_strnp_268 ( _zy_simnet_bimc_dbgcmd2_311_w$[0:9], 
	bimc_dbgcmd2[9:0]);
ixc_assign_32 _zz_strnp_267 ( _zy_simnet_bimc_pollrsp0_310_w$[0:31], 
	bimc_pollrsp0[31:0]);
ixc_assign_32 _zz_strnp_266 ( _zy_simnet_bimc_pollrsp1_309_w$[0:31], 
	bimc_pollrsp1[31:0]);
ixc_assign_10 _zz_strnp_265 ( _zy_simnet_bimc_pollrsp2_308_w$[0:9], 
	bimc_pollrsp2[9:0]);
ixc_assign_32 _zz_strnp_264 ( _zy_simnet_bimc_rxrsp0_307_w$[0:31], 
	bimc_rxrsp0[31:0]);
ixc_assign_32 _zz_strnp_263 ( _zy_simnet_bimc_rxrsp1_306_w$[0:31], 
	bimc_rxrsp1[31:0]);
ixc_assign_10 _zz_strnp_262 ( _zy_simnet_bimc_rxrsp2_305_w$[0:9], 
	bimc_rxrsp2[9:0]);
ixc_assign_32 _zz_strnp_261 ( _zy_simnet_bimc_rxcmd0_304_w$[0:31], 
	bimc_rxcmd0[31:0]);
ixc_assign_32 _zz_strnp_260 ( _zy_simnet_bimc_rxcmd1_303_w$[0:31], 
	bimc_rxcmd1[31:0]);
ixc_assign_10 _zz_strnp_259 ( _zy_simnet_bimc_rxcmd2_302_w$[0:9], 
	bimc_rxcmd2[9:0]);
ixc_assign_11 _zz_strnp_258 ( _zy_simnet_bimc_cmd2_301_w$[0:10], 
	bimc_cmd2[10:0]);
ixc_assign_29 _zz_strnp_257 ( _zy_simnet_bimc_eccpar_debug_300_w$[0:28], 
	bimc_eccpar_debug[28:0]);
ixc_assign_12 _zz_strnp_256 ( _zy_simnet_bimc_memid_299_w$[0:11], 
	bimc_memid[11:0]);
ixc_assign_32 _zz_strnp_255 ( _zy_simnet_bimc_global_config_298_w$[0:31], 
	bimc_global_config[31:0]);
ixc_assign_32 _zz_strnp_254 ( _zy_simnet_bimc_parity_error_cnt_297_w$[0:31], 
	bimc_parity_error_cnt[31:0]);
ixc_assign_32 _zz_strnp_253 ( 
	_zy_simnet_bimc_ecc_correctable_error_cnt_296_w$[0:31], 
	bimc_ecc_correctable_error_cnt[31:0]);
ixc_assign_32 _zz_strnp_252 ( 
	_zy_simnet_bimc_ecc_uncorrectable_error_cnt_295_w$[0:31], 
	bimc_ecc_uncorrectable_error_cnt[31:0]);
ixc_assign_7 _zz_strnp_251 ( _zy_simnet_bimc_monitor_294_w$[0:6], 
	bimc_monitor[6:0]);
ixc_assign_8 _zz_strnp_250 ( _zy_simnet_engine_sticky_status_293_w$[0:7], 
	engine_sticky_status[7:0]);
ixc_assign_5 _zz_strnp_249 ( _zy_simnet_interrupt_status_292_w$[0:4], 
	interrupt_status[4:0]);
ixc_assign_2 _zz_strnp_248 ( _zy_simnet_kdf_drbg_ctrl_291_w$[0:1], 
	kdf_drbg_ctrl[1:0]);
ixc_assign_17 _zz_strnp_247 ( _zy_simnet_kim_ia_rdata_part1_290_w$[0:16], 
	kim_ia_rdata_part1[16:0]);
ixc_assign_21 _zz_strnp_246 ( _zy_simnet_kim_ia_rdata_part0_289_w$[0:20], 
	kim_ia_rdata_part0[20:0]);
ixc_assign_22 _zz_strnp_245 ( _zy_simnet_kim_ia_status_288_w$[0:21], 
	kim_ia_status[21:0]);
ixc_assign_20 _zz_strnp_244 ( _zy_simnet_kim_ia_capability_287_w$[0:19], 
	kim_ia_capability[19:0]);
ixc_assign_32 _zz_strnp_243 ( _zy_simnet_ckv_ia_rdata_part1_286_w$[0:31], 
	ckv_ia_rdata_part1[31:0]);
ixc_assign_32 _zz_strnp_242 ( _zy_simnet_ckv_ia_rdata_part0_285_w$[0:31], 
	ckv_ia_rdata_part0[31:0]);
ixc_assign_23 _zz_strnp_241 ( _zy_simnet_ckv_ia_status_284_w$[0:22], 
	ckv_ia_status[22:0]);
ixc_assign_20 _zz_strnp_240 ( _zy_simnet_ckv_ia_capability_283_w$[0:19], 
	ckv_ia_capability[19:0]);
ixc_assign_12 _zz_strnp_239 ( _zy_simnet_cddip3_out_im_status_281_w$[0:11], 
	cddip3_out_im_status[11:0]);
ixc_assign_17 _zz_strnp_238 ( _zy_simnet_cddip3_out_ia_status_277_w$[0:16], 
	cddip3_out_ia_status[16:0]);
ixc_assign_20 _zz_strnp_237 ( _zy_simnet_cddip3_out_ia_capability_276_w$[0:19], 
	cddip3_out_ia_capability[19:0]);
ixc_assign_12 _zz_strnp_236 ( _zy_simnet_cddip2_out_im_status_274_w$[0:11], 
	cddip2_out_im_status[11:0]);
ixc_assign_17 _zz_strnp_235 ( _zy_simnet_cddip2_out_ia_status_270_w$[0:16], 
	cddip2_out_ia_status[16:0]);
ixc_assign_20 _zz_strnp_234 ( _zy_simnet_cddip2_out_ia_capability_269_w$[0:19], 
	cddip2_out_ia_capability[19:0]);
ixc_assign_12 _zz_strnp_233 ( _zy_simnet_cddip1_out_im_status_267_w$[0:11], 
	cddip1_out_im_status[11:0]);
ixc_assign_17 _zz_strnp_232 ( _zy_simnet_cddip1_out_ia_status_263_w$[0:16], 
	cddip1_out_ia_status[16:0]);
ixc_assign_20 _zz_strnp_231 ( _zy_simnet_cddip1_out_ia_capability_262_w$[0:19], 
	cddip1_out_ia_capability[19:0]);
ixc_assign_12 _zz_strnp_230 ( _zy_simnet_cddip0_out_im_status_260_w$[0:11], 
	cddip0_out_im_status[11:0]);
ixc_assign_17 _zz_strnp_229 ( _zy_simnet_cddip0_out_ia_status_256_w$[0:16], 
	cddip0_out_ia_status[16:0]);
ixc_assign_20 _zz_strnp_228 ( _zy_simnet_cddip0_out_ia_capability_255_w$[0:19], 
	cddip0_out_ia_capability[19:0]);
ixc_assign_12 _zz_strnp_227 ( _zy_simnet_cceip3_out_im_status_253_w$[0:11], 
	cceip3_out_im_status[11:0]);
ixc_assign_17 _zz_strnp_226 ( _zy_simnet_cceip3_out_ia_status_249_w$[0:16], 
	cceip3_out_ia_status[16:0]);
ixc_assign_20 _zz_strnp_225 ( _zy_simnet_cceip3_out_ia_capability_248_w$[0:19], 
	cceip3_out_ia_capability[19:0]);
ixc_assign_12 _zz_strnp_224 ( _zy_simnet_cceip2_out_im_status_246_w$[0:11], 
	cceip2_out_im_status[11:0]);
ixc_assign_17 _zz_strnp_223 ( _zy_simnet_cceip2_out_ia_status_242_w$[0:16], 
	cceip2_out_ia_status[16:0]);
ixc_assign_20 _zz_strnp_222 ( _zy_simnet_cceip2_out_ia_capability_241_w$[0:19], 
	cceip2_out_ia_capability[19:0]);
ixc_assign_12 _zz_strnp_221 ( _zy_simnet_cceip1_out_im_status_239_w$[0:11], 
	cceip1_out_im_status[11:0]);
ixc_assign_17 _zz_strnp_220 ( _zy_simnet_cceip1_out_ia_status_235_w$[0:16], 
	cceip1_out_ia_status[16:0]);
ixc_assign_20 _zz_strnp_219 ( _zy_simnet_cceip1_out_ia_capability_234_w$[0:19], 
	cceip1_out_ia_capability[19:0]);
ixc_assign_12 _zz_strnp_218 ( _zy_simnet_cceip0_out_im_status_232_w$[0:11], 
	cceip0_out_im_status[11:0]);
ixc_assign_17 _zz_strnp_217 ( _zy_simnet_cceip0_out_ia_status_228_w$[0:16], 
	cceip0_out_ia_status[16:0]);
ixc_assign_20 _zz_strnp_216 ( _zy_simnet_cceip0_out_ia_capability_227_w$[0:19], 
	cceip0_out_ia_capability[19:0]);
ixc_assign_32 _zz_strnp_215 ( _zy_simnet_tvar_226[0:31], { spare[31], 
	spare[30], spare[29], spare[28], spare[27], spare[26], spare[25], 
	spare[24], spare[23], spare[22], spare[21], spare[20], spare[19], 
	spare[18], spare[17], spare[16], spare[15], spare[14], spare[13], 
	spare[12], spare[11], spare[10], spare[9], spare[8], spare[7], 
	kdf_test_mode_en, always_validate_kim_ref, manual_txc, spare[3], 
	o_tready_override_val, disable_ckv_kim_ism_reads, send_kme_ib_beat});
ixc_assign_8 _zz_strnp_214 ( _zy_simnet_revid_wire_225_w$[0:7], 
	blkid_revid_config[7:0]);
ixc_assign_32 _zz_strnp_213 ( _zy_simnet_blkid_revid_config_224_w$[0:31], 
	blkid_revid_config[31:0]);
ixc_assign_9 _zz_strnp_212 ( sa_ctrl_ia_config[8:0], 
	_zy_simnet_sa_ctrl_ia_config_223_w$[0:8]);
ixc_assign_32 _zz_strnp_211 ( sa_ctrl_ia_wdata[31:0], 
	_zy_simnet_sa_ctrl_ia_wdata_222_w$[0:31]);
ixc_assign_32 _zz_strnp_210 ( sa_global_ctrl[31:0], 
	_zy_simnet_sa_global_ctrl_221_w$[0:31]);
ixc_assign_7 _zz_strnp_209 ( cddip_decrypt_kop_fifo_override[6:0], 
	_zy_simnet_cddip_decrypt_kop_fifo_override_220_w$[0:6]);
ixc_assign_7 _zz_strnp_208 ( cceip_validate_kop_fifo_override[6:0], 
	_zy_simnet_cceip_validate_kop_fifo_override_219_w$[0:6]);
ixc_assign_7 _zz_strnp_207 ( cceip_encrypt_kop_fifo_override[6:0], 
	_zy_simnet_cceip_encrypt_kop_fifo_override_218_w$[0:6]);
ixc_assign_9 _zz_strnp_206 ( sa_count_ia_config[8:0], 
	_zy_simnet_sa_count_ia_config_217_w$[0:8]);
ixc_assign_32 _zz_strnp_205 ( sa_count_ia_wdata[63:32], 
	_zy_simnet_sa_count_ia_wdata_216_w$[0:31]);
ixc_assign_32 _zz_strnp_204 ( sa_count_ia_wdata[31:0], 
	_zy_simnet_sa_count_ia_wdata_215_w$[0:31]);
ixc_assign_9 _zz_strnp_203 ( sa_snapshot_ia_config[8:0], 
	_zy_simnet_sa_snapshot_ia_config_214_w$[0:8]);
ixc_assign_32 _zz_strnp_202 ( sa_snapshot_ia_wdata[63:32], 
	_zy_simnet_sa_snapshot_ia_wdata_213_w$[0:31]);
ixc_assign_32 _zz_strnp_201 ( sa_snapshot_ia_wdata[31:0], 
	_zy_simnet_sa_snapshot_ia_wdata_212_w$[0:31]);
ixc_assign_32 _zz_strnp_200 ( regs_sa_ctrl[31:0], 
	_zy_simnet_regs_sa_ctrl_211_w$[0:31]);
ixc_assign_9 _zz_strnp_199 ( tready_override[8:0], 
	_zy_simnet_tready_override_210_w$[0:8]);
ixc_assign_10 _zz_strnp_198 ( o_bimc_dbgcmd2[9:0], 
	_zy_simnet_o_bimc_dbgcmd2_208_w$[0:9]);
ixc_assign_10 _zz_strnp_197 ( o_bimc_pollrsp2[9:0], 
	_zy_simnet_o_bimc_pollrsp2_207_w$[0:9]);
ixc_assign_10 _zz_strnp_196 ( o_bimc_rxrsp2[9:0], 
	_zy_simnet_o_bimc_rxrsp2_206_w$[0:9]);
ixc_assign_10 _zz_strnp_195 ( o_bimc_rxcmd2[9:0], 
	_zy_simnet_o_bimc_rxcmd2_205_w$[0:9]);
ixc_assign_32 _zz_strnp_194 ( o_bimc_cmd0[31:0], 
	_zy_simnet_o_bimc_cmd0_204_w$[0:31]);
ixc_assign_32 _zz_strnp_193 ( o_bimc_cmd1[31:0], 
	_zy_simnet_o_bimc_cmd1_203_w$[0:31]);
ixc_assign_11 _zz_strnp_192 ( o_bimc_cmd2[10:0], 
	_zy_simnet_o_bimc_cmd2_202_w$[0:10]);
ixc_assign_29 _zz_strnp_191 ( o_bimc_eccpar_debug[28:0], 
	_zy_simnet_o_bimc_eccpar_debug_201_w$[0:28]);
ixc_assign_32 _zz_strnp_190 ( o_bimc_global_config[31:0], 
	_zy_simnet_o_bimc_global_config_200_w$[0:31]);
ixc_assign_32 _zz_strnp_189 ( o_bimc_parity_error_cnt[31:0], 
	_zy_simnet_o_bimc_parity_error_cnt_199_w$[0:31]);
ixc_assign_32 _zz_strnp_188 ( o_bimc_ecc_correctable_error_cnt[31:0], 
	_zy_simnet_o_bimc_ecc_correctable_error_cnt_198_w$[0:31]);
ixc_assign_32 _zz_strnp_187 ( o_bimc_ecc_uncorrectable_error_cnt[31:0], 
	_zy_simnet_o_bimc_ecc_uncorrectable_error_cnt_197_w$[0:31]);
ixc_assign_7 _zz_strnp_186 ( o_bimc_monitor_mask[6:0], 
	_zy_simnet_o_bimc_monitor_mask_196_w$[0:6]);
ixc_assign_8 _zz_strnp_185 ( o_engine_sticky_status[7:0], 
	_zy_simnet_o_engine_sticky_status_195_w$[0:7]);
ixc_assign_5 _zz_strnp_184 ( o_interrupt_mask[4:0], 
	_zy_simnet_o_interrupt_mask_194_w$[0:4]);
ixc_assign_16 _zz_strnp_183 ( o_kdf_drbg_seed_1_reseed_interval_1[15:0], 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_1_192_w$[0:15]);
ixc_assign_32 _zz_strnp_182 ( o_kdf_drbg_seed_1_reseed_interval_0[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_reseed_interval_0_191_w$[0:31]);
ixc_assign_32 _zz_strnp_181 ( o_kdf_drbg_seed_1_state_value_127_96[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_127_96_190_w$[0:31]);
ixc_assign_32 _zz_strnp_180 ( o_kdf_drbg_seed_1_state_value_95_64[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_95_64_189_w$[0:31]);
ixc_assign_32 _zz_strnp_179 ( o_kdf_drbg_seed_1_state_value_63_32[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_63_32_188_w$[0:31]);
ixc_assign_32 _zz_strnp_178 ( o_kdf_drbg_seed_1_state_value_31_0[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_value_31_0_187_w$[0:31]);
ixc_assign_32 _zz_strnp_177 ( o_kdf_drbg_seed_1_state_key_255_224[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_255_224_186_w$[0:31]);
ixc_assign_32 _zz_strnp_176 ( o_kdf_drbg_seed_1_state_key_223_192[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_223_192_185_w$[0:31]);
ixc_assign_32 _zz_strnp_175 ( o_kdf_drbg_seed_1_state_key_191_160[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_191_160_184_w$[0:31]);
ixc_assign_32 _zz_strnp_174 ( o_kdf_drbg_seed_1_state_key_159_128[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_159_128_183_w$[0:31]);
ixc_assign_32 _zz_strnp_173 ( o_kdf_drbg_seed_1_state_key_127_96[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_127_96_182_w$[0:31]);
ixc_assign_32 _zz_strnp_172 ( o_kdf_drbg_seed_1_state_key_95_64[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_95_64_181_w$[0:31]);
ixc_assign_32 _zz_strnp_171 ( o_kdf_drbg_seed_1_state_key_63_32[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_63_32_180_w$[0:31]);
ixc_assign_32 _zz_strnp_170 ( o_kdf_drbg_seed_1_state_key_31_0[31:0], 
	_zy_simnet_o_kdf_drbg_seed_1_state_key_31_0_179_w$[0:31]);
ixc_assign_16 _zz_strnp_169 ( o_kdf_drbg_seed_0_reseed_interval_1[15:0], 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_1_178_w$[0:15]);
ixc_assign_32 _zz_strnp_168 ( o_kdf_drbg_seed_0_reseed_interval_0[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_reseed_interval_0_177_w$[0:31]);
ixc_assign_32 _zz_strnp_167 ( o_kdf_drbg_seed_0_state_value_127_96[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_127_96_176_w$[0:31]);
ixc_assign_32 _zz_strnp_166 ( o_kdf_drbg_seed_0_state_value_95_64[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_95_64_175_w$[0:31]);
ixc_assign_32 _zz_strnp_165 ( o_kdf_drbg_seed_0_state_value_63_32[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_63_32_174_w$[0:31]);
ixc_assign_32 _zz_strnp_164 ( o_kdf_drbg_seed_0_state_value_31_0[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_value_31_0_173_w$[0:31]);
ixc_assign_32 _zz_strnp_163 ( o_kdf_drbg_seed_0_state_key_255_224[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_255_224_172_w$[0:31]);
ixc_assign_32 _zz_strnp_162 ( o_kdf_drbg_seed_0_state_key_223_192[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_223_192_171_w$[0:31]);
ixc_assign_32 _zz_strnp_161 ( o_kdf_drbg_seed_0_state_key_191_160[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_191_160_170_w$[0:31]);
ixc_assign_32 _zz_strnp_160 ( o_kdf_drbg_seed_0_state_key_159_128[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_159_128_169_w$[0:31]);
ixc_assign_32 _zz_strnp_159 ( o_kdf_drbg_seed_0_state_key_127_96[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_127_96_168_w$[0:31]);
ixc_assign_32 _zz_strnp_158 ( o_kdf_drbg_seed_0_state_key_95_64[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_95_64_167_w$[0:31]);
ixc_assign_32 _zz_strnp_157 ( o_kdf_drbg_seed_0_state_key_63_32[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_63_32_166_w$[0:31]);
ixc_assign_32 _zz_strnp_156 ( o_kdf_drbg_seed_0_state_key_31_0[31:0], 
	_zy_simnet_o_kdf_drbg_seed_0_state_key_31_0_165_w$[0:31]);
ixc_assign_2 _zz_strnp_155 ( o_kdf_drbg_ctrl[1:0], 
	_zy_simnet_o_kdf_drbg_ctrl_164_w$[0:1]);
ixc_assign_32 _zz_strnp_154 ( { \labels[7][40] , \labels[7][39] , 
	\labels[7][38] , \labels[7][37] , \labels[7][36] , \labels[7][35] , 
	\labels[7][34] , \labels[7][33] , \labels[7][32] , \labels[7][31] , 
	\labels[7][30] , \labels[7][29] , \labels[7][28] , \labels[7][27] , 
	\labels[7][26] , \labels[7][25] , \labels[7][24] , \labels[7][23] , 
	\labels[7][22] , \labels[7][21] , \labels[7][20] , \labels[7][19] , 
	\labels[7][18] , \labels[7][17] , \labels[7][16] , \labels[7][15] , 
	\labels[7][14] , \labels[7][13] , \labels[7][12] , \labels[7][11] , 
	\labels[7][10] , \labels[7][9] }, _zy_simnet_labels_163_w$[0:31]);
ixc_assign_32 _zz_strnp_153 ( { \labels[7][72] , \labels[7][71] , 
	\labels[7][70] , \labels[7][69] , \labels[7][68] , \labels[7][67] , 
	\labels[7][66] , \labels[7][65] , \labels[7][64] , \labels[7][63] , 
	\labels[7][62] , \labels[7][61] , \labels[7][60] , \labels[7][59] , 
	\labels[7][58] , \labels[7][57] , \labels[7][56] , \labels[7][55] , 
	\labels[7][54] , \labels[7][53] , \labels[7][52] , \labels[7][51] , 
	\labels[7][50] , \labels[7][49] , \labels[7][48] , \labels[7][47] , 
	\labels[7][46] , \labels[7][45] , \labels[7][44] , \labels[7][43] , 
	\labels[7][42] , \labels[7][41] }, _zy_simnet_labels_162_w$[0:31]);
ixc_assign_32 _zz_strnp_152 ( { \labels[7][104] , \labels[7][103] , 
	\labels[7][102] , \labels[7][101] , \labels[7][100] , 
	\labels[7][99] , \labels[7][98] , \labels[7][97] , \labels[7][96] , 
	\labels[7][95] , \labels[7][94] , \labels[7][93] , \labels[7][92] , 
	\labels[7][91] , \labels[7][90] , \labels[7][89] , \labels[7][88] , 
	\labels[7][87] , \labels[7][86] , \labels[7][85] , \labels[7][84] , 
	\labels[7][83] , \labels[7][82] , \labels[7][81] , \labels[7][80] , 
	\labels[7][79] , \labels[7][78] , \labels[7][77] , \labels[7][76] , 
	\labels[7][75] , \labels[7][74] , \labels[7][73] }, 
	_zy_simnet_labels_161_w$[0:31]);
ixc_assign_32 _zz_strnp_151 ( { \labels[7][136] , \labels[7][135] , 
	\labels[7][134] , \labels[7][133] , \labels[7][132] , 
	\labels[7][131] , \labels[7][130] , \labels[7][129] , 
	\labels[7][128] , \labels[7][127] , \labels[7][126] , 
	\labels[7][125] , \labels[7][124] , \labels[7][123] , 
	\labels[7][122] , \labels[7][121] , \labels[7][120] , 
	\labels[7][119] , \labels[7][118] , \labels[7][117] , 
	\labels[7][116] , \labels[7][115] , \labels[7][114] , 
	\labels[7][113] , \labels[7][112] , \labels[7][111] , 
	\labels[7][110] , \labels[7][109] , \labels[7][108] , 
	\labels[7][107] , \labels[7][106] , \labels[7][105] }, 
	_zy_simnet_labels_160_w$[0:31]);
ixc_assign_32 _zz_strnp_150 ( { \labels[7][168] , \labels[7][167] , 
	\labels[7][166] , \labels[7][165] , \labels[7][164] , 
	\labels[7][163] , \labels[7][162] , \labels[7][161] , 
	\labels[7][160] , \labels[7][159] , \labels[7][158] , 
	\labels[7][157] , \labels[7][156] , \labels[7][155] , 
	\labels[7][154] , \labels[7][153] , \labels[7][152] , 
	\labels[7][151] , \labels[7][150] , \labels[7][149] , 
	\labels[7][148] , \labels[7][147] , \labels[7][146] , 
	\labels[7][145] , \labels[7][144] , \labels[7][143] , 
	\labels[7][142] , \labels[7][141] , \labels[7][140] , 
	\labels[7][139] , \labels[7][138] , \labels[7][137] }, 
	_zy_simnet_labels_159_w$[0:31]);
ixc_assign_32 _zz_strnp_149 ( { \labels[7][200] , \labels[7][199] , 
	\labels[7][198] , \labels[7][197] , \labels[7][196] , 
	\labels[7][195] , \labels[7][194] , \labels[7][193] , 
	\labels[7][192] , \labels[7][191] , \labels[7][190] , 
	\labels[7][189] , \labels[7][188] , \labels[7][187] , 
	\labels[7][186] , \labels[7][185] , \labels[7][184] , 
	\labels[7][183] , \labels[7][182] , \labels[7][181] , 
	\labels[7][180] , \labels[7][179] , \labels[7][178] , 
	\labels[7][177] , \labels[7][176] , \labels[7][175] , 
	\labels[7][174] , \labels[7][173] , \labels[7][172] , 
	\labels[7][171] , \labels[7][170] , \labels[7][169] }, 
	_zy_simnet_labels_158_w$[0:31]);
ixc_assign_32 _zz_strnp_148 ( { \labels[7][232] , \labels[7][231] , 
	\labels[7][230] , \labels[7][229] , \labels[7][228] , 
	\labels[7][227] , \labels[7][226] , \labels[7][225] , 
	\labels[7][224] , \labels[7][223] , \labels[7][222] , 
	\labels[7][221] , \labels[7][220] , \labels[7][219] , 
	\labels[7][218] , \labels[7][217] , \labels[7][216] , 
	\labels[7][215] , \labels[7][214] , \labels[7][213] , 
	\labels[7][212] , \labels[7][211] , \labels[7][210] , 
	\labels[7][209] , \labels[7][208] , \labels[7][207] , 
	\labels[7][206] , \labels[7][205] , \labels[7][204] , 
	\labels[7][203] , \labels[7][202] , \labels[7][201] }, 
	_zy_simnet_labels_157_w$[0:31]);
ixc_assign_32 _zz_strnp_147 ( { \labels[7][264] , \labels[7][263] , 
	\labels[7][262] , \labels[7][261] , \labels[7][260] , 
	\labels[7][259] , \labels[7][258] , \labels[7][257] , 
	\labels[7][256] , \labels[7][255] , \labels[7][254] , 
	\labels[7][253] , \labels[7][252] , \labels[7][251] , 
	\labels[7][250] , \labels[7][249] , \labels[7][248] , 
	\labels[7][247] , \labels[7][246] , \labels[7][245] , 
	\labels[7][244] , \labels[7][243] , \labels[7][242] , 
	\labels[7][241] , \labels[7][240] , \labels[7][239] , 
	\labels[7][238] , \labels[7][237] , \labels[7][236] , 
	\labels[7][235] , \labels[7][234] , \labels[7][233] }, 
	_zy_simnet_labels_156_w$[0:31]);
ixc_assign_16 _zz_strnp_146 ( { \labels[7][271] , \labels[7][270] , 
	\labels[7][269] , \labels[7][268] , \labels[7][267] , 
	\labels[7][266] , \labels[7][265] , \labels[7][8] , \labels[7][7] , 
	\labels[7][6] , \labels[7][5] , \labels[7][4] , \labels[7][3] , 
	\labels[7][2] , \labels[7][1] , \labels[7][0] }, 
	_zy_simnet_tvar_155[0:15]);
ixc_assign_32 _zz_strnp_145 ( { \labels[6][40] , \labels[6][39] , 
	\labels[6][38] , \labels[6][37] , \labels[6][36] , \labels[6][35] , 
	\labels[6][34] , \labels[6][33] , \labels[6][32] , \labels[6][31] , 
	\labels[6][30] , \labels[6][29] , \labels[6][28] , \labels[6][27] , 
	\labels[6][26] , \labels[6][25] , \labels[6][24] , \labels[6][23] , 
	\labels[6][22] , \labels[6][21] , \labels[6][20] , \labels[6][19] , 
	\labels[6][18] , \labels[6][17] , \labels[6][16] , \labels[6][15] , 
	\labels[6][14] , \labels[6][13] , \labels[6][12] , \labels[6][11] , 
	\labels[6][10] , \labels[6][9] }, _zy_simnet_labels_154_w$[0:31]);
ixc_assign_32 _zz_strnp_144 ( { \labels[6][72] , \labels[6][71] , 
	\labels[6][70] , \labels[6][69] , \labels[6][68] , \labels[6][67] , 
	\labels[6][66] , \labels[6][65] , \labels[6][64] , \labels[6][63] , 
	\labels[6][62] , \labels[6][61] , \labels[6][60] , \labels[6][59] , 
	\labels[6][58] , \labels[6][57] , \labels[6][56] , \labels[6][55] , 
	\labels[6][54] , \labels[6][53] , \labels[6][52] , \labels[6][51] , 
	\labels[6][50] , \labels[6][49] , \labels[6][48] , \labels[6][47] , 
	\labels[6][46] , \labels[6][45] , \labels[6][44] , \labels[6][43] , 
	\labels[6][42] , \labels[6][41] }, _zy_simnet_labels_153_w$[0:31]);
ixc_assign_32 _zz_strnp_143 ( { \labels[6][104] , \labels[6][103] , 
	\labels[6][102] , \labels[6][101] , \labels[6][100] , 
	\labels[6][99] , \labels[6][98] , \labels[6][97] , \labels[6][96] , 
	\labels[6][95] , \labels[6][94] , \labels[6][93] , \labels[6][92] , 
	\labels[6][91] , \labels[6][90] , \labels[6][89] , \labels[6][88] , 
	\labels[6][87] , \labels[6][86] , \labels[6][85] , \labels[6][84] , 
	\labels[6][83] , \labels[6][82] , \labels[6][81] , \labels[6][80] , 
	\labels[6][79] , \labels[6][78] , \labels[6][77] , \labels[6][76] , 
	\labels[6][75] , \labels[6][74] , \labels[6][73] }, 
	_zy_simnet_labels_152_w$[0:31]);
ixc_assign_32 _zz_strnp_142 ( { \labels[6][136] , \labels[6][135] , 
	\labels[6][134] , \labels[6][133] , \labels[6][132] , 
	\labels[6][131] , \labels[6][130] , \labels[6][129] , 
	\labels[6][128] , \labels[6][127] , \labels[6][126] , 
	\labels[6][125] , \labels[6][124] , \labels[6][123] , 
	\labels[6][122] , \labels[6][121] , \labels[6][120] , 
	\labels[6][119] , \labels[6][118] , \labels[6][117] , 
	\labels[6][116] , \labels[6][115] , \labels[6][114] , 
	\labels[6][113] , \labels[6][112] , \labels[6][111] , 
	\labels[6][110] , \labels[6][109] , \labels[6][108] , 
	\labels[6][107] , \labels[6][106] , \labels[6][105] }, 
	_zy_simnet_labels_151_w$[0:31]);
ixc_assign_32 _zz_strnp_141 ( { \labels[6][168] , \labels[6][167] , 
	\labels[6][166] , \labels[6][165] , \labels[6][164] , 
	\labels[6][163] , \labels[6][162] , \labels[6][161] , 
	\labels[6][160] , \labels[6][159] , \labels[6][158] , 
	\labels[6][157] , \labels[6][156] , \labels[6][155] , 
	\labels[6][154] , \labels[6][153] , \labels[6][152] , 
	\labels[6][151] , \labels[6][150] , \labels[6][149] , 
	\labels[6][148] , \labels[6][147] , \labels[6][146] , 
	\labels[6][145] , \labels[6][144] , \labels[6][143] , 
	\labels[6][142] , \labels[6][141] , \labels[6][140] , 
	\labels[6][139] , \labels[6][138] , \labels[6][137] }, 
	_zy_simnet_labels_150_w$[0:31]);
ixc_assign_32 _zz_strnp_140 ( { \labels[6][200] , \labels[6][199] , 
	\labels[6][198] , \labels[6][197] , \labels[6][196] , 
	\labels[6][195] , \labels[6][194] , \labels[6][193] , 
	\labels[6][192] , \labels[6][191] , \labels[6][190] , 
	\labels[6][189] , \labels[6][188] , \labels[6][187] , 
	\labels[6][186] , \labels[6][185] , \labels[6][184] , 
	\labels[6][183] , \labels[6][182] , \labels[6][181] , 
	\labels[6][180] , \labels[6][179] , \labels[6][178] , 
	\labels[6][177] , \labels[6][176] , \labels[6][175] , 
	\labels[6][174] , \labels[6][173] , \labels[6][172] , 
	\labels[6][171] , \labels[6][170] , \labels[6][169] }, 
	_zy_simnet_labels_149_w$[0:31]);
ixc_assign_32 _zz_strnp_139 ( { \labels[6][232] , \labels[6][231] , 
	\labels[6][230] , \labels[6][229] , \labels[6][228] , 
	\labels[6][227] , \labels[6][226] , \labels[6][225] , 
	\labels[6][224] , \labels[6][223] , \labels[6][222] , 
	\labels[6][221] , \labels[6][220] , \labels[6][219] , 
	\labels[6][218] , \labels[6][217] , \labels[6][216] , 
	\labels[6][215] , \labels[6][214] , \labels[6][213] , 
	\labels[6][212] , \labels[6][211] , \labels[6][210] , 
	\labels[6][209] , \labels[6][208] , \labels[6][207] , 
	\labels[6][206] , \labels[6][205] , \labels[6][204] , 
	\labels[6][203] , \labels[6][202] , \labels[6][201] }, 
	_zy_simnet_labels_148_w$[0:31]);
ixc_assign_32 _zz_strnp_138 ( { \labels[6][264] , \labels[6][263] , 
	\labels[6][262] , \labels[6][261] , \labels[6][260] , 
	\labels[6][259] , \labels[6][258] , \labels[6][257] , 
	\labels[6][256] , \labels[6][255] , \labels[6][254] , 
	\labels[6][253] , \labels[6][252] , \labels[6][251] , 
	\labels[6][250] , \labels[6][249] , \labels[6][248] , 
	\labels[6][247] , \labels[6][246] , \labels[6][245] , 
	\labels[6][244] , \labels[6][243] , \labels[6][242] , 
	\labels[6][241] , \labels[6][240] , \labels[6][239] , 
	\labels[6][238] , \labels[6][237] , \labels[6][236] , 
	\labels[6][235] , \labels[6][234] , \labels[6][233] }, 
	_zy_simnet_labels_147_w$[0:31]);
ixc_assign_16 _zz_strnp_137 ( { \labels[6][271] , \labels[6][270] , 
	\labels[6][269] , \labels[6][268] , \labels[6][267] , 
	\labels[6][266] , \labels[6][265] , \labels[6][8] , \labels[6][7] , 
	\labels[6][6] , \labels[6][5] , \labels[6][4] , \labels[6][3] , 
	\labels[6][2] , \labels[6][1] , \labels[6][0] }, 
	_zy_simnet_tvar_146[0:15]);
ixc_assign_32 _zz_strnp_136 ( { \labels[5][40] , \labels[5][39] , 
	\labels[5][38] , \labels[5][37] , \labels[5][36] , \labels[5][35] , 
	\labels[5][34] , \labels[5][33] , \labels[5][32] , \labels[5][31] , 
	\labels[5][30] , \labels[5][29] , \labels[5][28] , \labels[5][27] , 
	\labels[5][26] , \labels[5][25] , \labels[5][24] , \labels[5][23] , 
	\labels[5][22] , \labels[5][21] , \labels[5][20] , \labels[5][19] , 
	\labels[5][18] , \labels[5][17] , \labels[5][16] , \labels[5][15] , 
	\labels[5][14] , \labels[5][13] , \labels[5][12] , \labels[5][11] , 
	\labels[5][10] , \labels[5][9] }, _zy_simnet_labels_145_w$[0:31]);
ixc_assign_32 _zz_strnp_135 ( { \labels[5][72] , \labels[5][71] , 
	\labels[5][70] , \labels[5][69] , \labels[5][68] , \labels[5][67] , 
	\labels[5][66] , \labels[5][65] , \labels[5][64] , \labels[5][63] , 
	\labels[5][62] , \labels[5][61] , \labels[5][60] , \labels[5][59] , 
	\labels[5][58] , \labels[5][57] , \labels[5][56] , \labels[5][55] , 
	\labels[5][54] , \labels[5][53] , \labels[5][52] , \labels[5][51] , 
	\labels[5][50] , \labels[5][49] , \labels[5][48] , \labels[5][47] , 
	\labels[5][46] , \labels[5][45] , \labels[5][44] , \labels[5][43] , 
	\labels[5][42] , \labels[5][41] }, _zy_simnet_labels_144_w$[0:31]);
ixc_assign_32 _zz_strnp_134 ( { \labels[5][104] , \labels[5][103] , 
	\labels[5][102] , \labels[5][101] , \labels[5][100] , 
	\labels[5][99] , \labels[5][98] , \labels[5][97] , \labels[5][96] , 
	\labels[5][95] , \labels[5][94] , \labels[5][93] , \labels[5][92] , 
	\labels[5][91] , \labels[5][90] , \labels[5][89] , \labels[5][88] , 
	\labels[5][87] , \labels[5][86] , \labels[5][85] , \labels[5][84] , 
	\labels[5][83] , \labels[5][82] , \labels[5][81] , \labels[5][80] , 
	\labels[5][79] , \labels[5][78] , \labels[5][77] , \labels[5][76] , 
	\labels[5][75] , \labels[5][74] , \labels[5][73] }, 
	_zy_simnet_labels_143_w$[0:31]);
ixc_assign_32 _zz_strnp_133 ( { \labels[5][136] , \labels[5][135] , 
	\labels[5][134] , \labels[5][133] , \labels[5][132] , 
	\labels[5][131] , \labels[5][130] , \labels[5][129] , 
	\labels[5][128] , \labels[5][127] , \labels[5][126] , 
	\labels[5][125] , \labels[5][124] , \labels[5][123] , 
	\labels[5][122] , \labels[5][121] , \labels[5][120] , 
	\labels[5][119] , \labels[5][118] , \labels[5][117] , 
	\labels[5][116] , \labels[5][115] , \labels[5][114] , 
	\labels[5][113] , \labels[5][112] , \labels[5][111] , 
	\labels[5][110] , \labels[5][109] , \labels[5][108] , 
	\labels[5][107] , \labels[5][106] , \labels[5][105] }, 
	_zy_simnet_labels_142_w$[0:31]);
ixc_assign_32 _zz_strnp_132 ( { \labels[5][168] , \labels[5][167] , 
	\labels[5][166] , \labels[5][165] , \labels[5][164] , 
	\labels[5][163] , \labels[5][162] , \labels[5][161] , 
	\labels[5][160] , \labels[5][159] , \labels[5][158] , 
	\labels[5][157] , \labels[5][156] , \labels[5][155] , 
	\labels[5][154] , \labels[5][153] , \labels[5][152] , 
	\labels[5][151] , \labels[5][150] , \labels[5][149] , 
	\labels[5][148] , \labels[5][147] , \labels[5][146] , 
	\labels[5][145] , \labels[5][144] , \labels[5][143] , 
	\labels[5][142] , \labels[5][141] , \labels[5][140] , 
	\labels[5][139] , \labels[5][138] , \labels[5][137] }, 
	_zy_simnet_labels_141_w$[0:31]);
ixc_assign_32 _zz_strnp_131 ( { \labels[5][200] , \labels[5][199] , 
	\labels[5][198] , \labels[5][197] , \labels[5][196] , 
	\labels[5][195] , \labels[5][194] , \labels[5][193] , 
	\labels[5][192] , \labels[5][191] , \labels[5][190] , 
	\labels[5][189] , \labels[5][188] , \labels[5][187] , 
	\labels[5][186] , \labels[5][185] , \labels[5][184] , 
	\labels[5][183] , \labels[5][182] , \labels[5][181] , 
	\labels[5][180] , \labels[5][179] , \labels[5][178] , 
	\labels[5][177] , \labels[5][176] , \labels[5][175] , 
	\labels[5][174] , \labels[5][173] , \labels[5][172] , 
	\labels[5][171] , \labels[5][170] , \labels[5][169] }, 
	_zy_simnet_labels_140_w$[0:31]);
ixc_assign_32 _zz_strnp_130 ( { \labels[5][232] , \labels[5][231] , 
	\labels[5][230] , \labels[5][229] , \labels[5][228] , 
	\labels[5][227] , \labels[5][226] , \labels[5][225] , 
	\labels[5][224] , \labels[5][223] , \labels[5][222] , 
	\labels[5][221] , \labels[5][220] , \labels[5][219] , 
	\labels[5][218] , \labels[5][217] , \labels[5][216] , 
	\labels[5][215] , \labels[5][214] , \labels[5][213] , 
	\labels[5][212] , \labels[5][211] , \labels[5][210] , 
	\labels[5][209] , \labels[5][208] , \labels[5][207] , 
	\labels[5][206] , \labels[5][205] , \labels[5][204] , 
	\labels[5][203] , \labels[5][202] , \labels[5][201] }, 
	_zy_simnet_labels_139_w$[0:31]);
ixc_assign_32 _zz_strnp_129 ( { \labels[5][264] , \labels[5][263] , 
	\labels[5][262] , \labels[5][261] , \labels[5][260] , 
	\labels[5][259] , \labels[5][258] , \labels[5][257] , 
	\labels[5][256] , \labels[5][255] , \labels[5][254] , 
	\labels[5][253] , \labels[5][252] , \labels[5][251] , 
	\labels[5][250] , \labels[5][249] , \labels[5][248] , 
	\labels[5][247] , \labels[5][246] , \labels[5][245] , 
	\labels[5][244] , \labels[5][243] , \labels[5][242] , 
	\labels[5][241] , \labels[5][240] , \labels[5][239] , 
	\labels[5][238] , \labels[5][237] , \labels[5][236] , 
	\labels[5][235] , \labels[5][234] , \labels[5][233] }, 
	_zy_simnet_labels_138_w$[0:31]);
ixc_assign_16 _zz_strnp_128 ( { \labels[5][271] , \labels[5][270] , 
	\labels[5][269] , \labels[5][268] , \labels[5][267] , 
	\labels[5][266] , \labels[5][265] , \labels[5][8] , \labels[5][7] , 
	\labels[5][6] , \labels[5][5] , \labels[5][4] , \labels[5][3] , 
	\labels[5][2] , \labels[5][1] , \labels[5][0] }, 
	_zy_simnet_tvar_137[0:15]);
ixc_assign_32 _zz_strnp_127 ( { \labels[4][40] , \labels[4][39] , 
	\labels[4][38] , \labels[4][37] , \labels[4][36] , \labels[4][35] , 
	\labels[4][34] , \labels[4][33] , \labels[4][32] , \labels[4][31] , 
	\labels[4][30] , \labels[4][29] , \labels[4][28] , \labels[4][27] , 
	\labels[4][26] , \labels[4][25] , \labels[4][24] , \labels[4][23] , 
	\labels[4][22] , \labels[4][21] , \labels[4][20] , \labels[4][19] , 
	\labels[4][18] , \labels[4][17] , \labels[4][16] , \labels[4][15] , 
	\labels[4][14] , \labels[4][13] , \labels[4][12] , \labels[4][11] , 
	\labels[4][10] , \labels[4][9] }, _zy_simnet_labels_136_w$[0:31]);
ixc_assign_32 _zz_strnp_126 ( { \labels[4][72] , \labels[4][71] , 
	\labels[4][70] , \labels[4][69] , \labels[4][68] , \labels[4][67] , 
	\labels[4][66] , \labels[4][65] , \labels[4][64] , \labels[4][63] , 
	\labels[4][62] , \labels[4][61] , \labels[4][60] , \labels[4][59] , 
	\labels[4][58] , \labels[4][57] , \labels[4][56] , \labels[4][55] , 
	\labels[4][54] , \labels[4][53] , \labels[4][52] , \labels[4][51] , 
	\labels[4][50] , \labels[4][49] , \labels[4][48] , \labels[4][47] , 
	\labels[4][46] , \labels[4][45] , \labels[4][44] , \labels[4][43] , 
	\labels[4][42] , \labels[4][41] }, _zy_simnet_labels_135_w$[0:31]);
ixc_assign_32 _zz_strnp_125 ( { \labels[4][104] , \labels[4][103] , 
	\labels[4][102] , \labels[4][101] , \labels[4][100] , 
	\labels[4][99] , \labels[4][98] , \labels[4][97] , \labels[4][96] , 
	\labels[4][95] , \labels[4][94] , \labels[4][93] , \labels[4][92] , 
	\labels[4][91] , \labels[4][90] , \labels[4][89] , \labels[4][88] , 
	\labels[4][87] , \labels[4][86] , \labels[4][85] , \labels[4][84] , 
	\labels[4][83] , \labels[4][82] , \labels[4][81] , \labels[4][80] , 
	\labels[4][79] , \labels[4][78] , \labels[4][77] , \labels[4][76] , 
	\labels[4][75] , \labels[4][74] , \labels[4][73] }, 
	_zy_simnet_labels_134_w$[0:31]);
ixc_assign_32 _zz_strnp_124 ( { \labels[4][136] , \labels[4][135] , 
	\labels[4][134] , \labels[4][133] , \labels[4][132] , 
	\labels[4][131] , \labels[4][130] , \labels[4][129] , 
	\labels[4][128] , \labels[4][127] , \labels[4][126] , 
	\labels[4][125] , \labels[4][124] , \labels[4][123] , 
	\labels[4][122] , \labels[4][121] , \labels[4][120] , 
	\labels[4][119] , \labels[4][118] , \labels[4][117] , 
	\labels[4][116] , \labels[4][115] , \labels[4][114] , 
	\labels[4][113] , \labels[4][112] , \labels[4][111] , 
	\labels[4][110] , \labels[4][109] , \labels[4][108] , 
	\labels[4][107] , \labels[4][106] , \labels[4][105] }, 
	_zy_simnet_labels_133_w$[0:31]);
ixc_assign_32 _zz_strnp_123 ( { \labels[4][168] , \labels[4][167] , 
	\labels[4][166] , \labels[4][165] , \labels[4][164] , 
	\labels[4][163] , \labels[4][162] , \labels[4][161] , 
	\labels[4][160] , \labels[4][159] , \labels[4][158] , 
	\labels[4][157] , \labels[4][156] , \labels[4][155] , 
	\labels[4][154] , \labels[4][153] , \labels[4][152] , 
	\labels[4][151] , \labels[4][150] , \labels[4][149] , 
	\labels[4][148] , \labels[4][147] , \labels[4][146] , 
	\labels[4][145] , \labels[4][144] , \labels[4][143] , 
	\labels[4][142] , \labels[4][141] , \labels[4][140] , 
	\labels[4][139] , \labels[4][138] , \labels[4][137] }, 
	_zy_simnet_labels_132_w$[0:31]);
ixc_assign_32 _zz_strnp_122 ( { \labels[4][200] , \labels[4][199] , 
	\labels[4][198] , \labels[4][197] , \labels[4][196] , 
	\labels[4][195] , \labels[4][194] , \labels[4][193] , 
	\labels[4][192] , \labels[4][191] , \labels[4][190] , 
	\labels[4][189] , \labels[4][188] , \labels[4][187] , 
	\labels[4][186] , \labels[4][185] , \labels[4][184] , 
	\labels[4][183] , \labels[4][182] , \labels[4][181] , 
	\labels[4][180] , \labels[4][179] , \labels[4][178] , 
	\labels[4][177] , \labels[4][176] , \labels[4][175] , 
	\labels[4][174] , \labels[4][173] , \labels[4][172] , 
	\labels[4][171] , \labels[4][170] , \labels[4][169] }, 
	_zy_simnet_labels_131_w$[0:31]);
ixc_assign_32 _zz_strnp_121 ( { \labels[4][232] , \labels[4][231] , 
	\labels[4][230] , \labels[4][229] , \labels[4][228] , 
	\labels[4][227] , \labels[4][226] , \labels[4][225] , 
	\labels[4][224] , \labels[4][223] , \labels[4][222] , 
	\labels[4][221] , \labels[4][220] , \labels[4][219] , 
	\labels[4][218] , \labels[4][217] , \labels[4][216] , 
	\labels[4][215] , \labels[4][214] , \labels[4][213] , 
	\labels[4][212] , \labels[4][211] , \labels[4][210] , 
	\labels[4][209] , \labels[4][208] , \labels[4][207] , 
	\labels[4][206] , \labels[4][205] , \labels[4][204] , 
	\labels[4][203] , \labels[4][202] , \labels[4][201] }, 
	_zy_simnet_labels_130_w$[0:31]);
ixc_assign_32 _zz_strnp_120 ( { \labels[4][264] , \labels[4][263] , 
	\labels[4][262] , \labels[4][261] , \labels[4][260] , 
	\labels[4][259] , \labels[4][258] , \labels[4][257] , 
	\labels[4][256] , \labels[4][255] , \labels[4][254] , 
	\labels[4][253] , \labels[4][252] , \labels[4][251] , 
	\labels[4][250] , \labels[4][249] , \labels[4][248] , 
	\labels[4][247] , \labels[4][246] , \labels[4][245] , 
	\labels[4][244] , \labels[4][243] , \labels[4][242] , 
	\labels[4][241] , \labels[4][240] , \labels[4][239] , 
	\labels[4][238] , \labels[4][237] , \labels[4][236] , 
	\labels[4][235] , \labels[4][234] , \labels[4][233] }, 
	_zy_simnet_labels_129_w$[0:31]);
ixc_assign_16 _zz_strnp_119 ( { \labels[4][271] , \labels[4][270] , 
	\labels[4][269] , \labels[4][268] , \labels[4][267] , 
	\labels[4][266] , \labels[4][265] , \labels[4][8] , \labels[4][7] , 
	\labels[4][6] , \labels[4][5] , \labels[4][4] , \labels[4][3] , 
	\labels[4][2] , \labels[4][1] , \labels[4][0] }, 
	_zy_simnet_tvar_128[0:15]);
ixc_assign_32 _zz_strnp_118 ( { \labels[3][40] , \labels[3][39] , 
	\labels[3][38] , \labels[3][37] , \labels[3][36] , \labels[3][35] , 
	\labels[3][34] , \labels[3][33] , \labels[3][32] , \labels[3][31] , 
	\labels[3][30] , \labels[3][29] , \labels[3][28] , \labels[3][27] , 
	\labels[3][26] , \labels[3][25] , \labels[3][24] , \labels[3][23] , 
	\labels[3][22] , \labels[3][21] , \labels[3][20] , \labels[3][19] , 
	\labels[3][18] , \labels[3][17] , \labels[3][16] , \labels[3][15] , 
	\labels[3][14] , \labels[3][13] , \labels[3][12] , \labels[3][11] , 
	\labels[3][10] , \labels[3][9] }, _zy_simnet_labels_127_w$[0:31]);
ixc_assign_32 _zz_strnp_117 ( { \labels[3][72] , \labels[3][71] , 
	\labels[3][70] , \labels[3][69] , \labels[3][68] , \labels[3][67] , 
	\labels[3][66] , \labels[3][65] , \labels[3][64] , \labels[3][63] , 
	\labels[3][62] , \labels[3][61] , \labels[3][60] , \labels[3][59] , 
	\labels[3][58] , \labels[3][57] , \labels[3][56] , \labels[3][55] , 
	\labels[3][54] , \labels[3][53] , \labels[3][52] , \labels[3][51] , 
	\labels[3][50] , \labels[3][49] , \labels[3][48] , \labels[3][47] , 
	\labels[3][46] , \labels[3][45] , \labels[3][44] , \labels[3][43] , 
	\labels[3][42] , \labels[3][41] }, _zy_simnet_labels_126_w$[0:31]);
ixc_assign_32 _zz_strnp_116 ( { \labels[3][104] , \labels[3][103] , 
	\labels[3][102] , \labels[3][101] , \labels[3][100] , 
	\labels[3][99] , \labels[3][98] , \labels[3][97] , \labels[3][96] , 
	\labels[3][95] , \labels[3][94] , \labels[3][93] , \labels[3][92] , 
	\labels[3][91] , \labels[3][90] , \labels[3][89] , \labels[3][88] , 
	\labels[3][87] , \labels[3][86] , \labels[3][85] , \labels[3][84] , 
	\labels[3][83] , \labels[3][82] , \labels[3][81] , \labels[3][80] , 
	\labels[3][79] , \labels[3][78] , \labels[3][77] , \labels[3][76] , 
	\labels[3][75] , \labels[3][74] , \labels[3][73] }, 
	_zy_simnet_labels_125_w$[0:31]);
ixc_assign_32 _zz_strnp_115 ( { \labels[3][136] , \labels[3][135] , 
	\labels[3][134] , \labels[3][133] , \labels[3][132] , 
	\labels[3][131] , \labels[3][130] , \labels[3][129] , 
	\labels[3][128] , \labels[3][127] , \labels[3][126] , 
	\labels[3][125] , \labels[3][124] , \labels[3][123] , 
	\labels[3][122] , \labels[3][121] , \labels[3][120] , 
	\labels[3][119] , \labels[3][118] , \labels[3][117] , 
	\labels[3][116] , \labels[3][115] , \labels[3][114] , 
	\labels[3][113] , \labels[3][112] , \labels[3][111] , 
	\labels[3][110] , \labels[3][109] , \labels[3][108] , 
	\labels[3][107] , \labels[3][106] , \labels[3][105] }, 
	_zy_simnet_labels_124_w$[0:31]);
ixc_assign_32 _zz_strnp_114 ( { \labels[3][168] , \labels[3][167] , 
	\labels[3][166] , \labels[3][165] , \labels[3][164] , 
	\labels[3][163] , \labels[3][162] , \labels[3][161] , 
	\labels[3][160] , \labels[3][159] , \labels[3][158] , 
	\labels[3][157] , \labels[3][156] , \labels[3][155] , 
	\labels[3][154] , \labels[3][153] , \labels[3][152] , 
	\labels[3][151] , \labels[3][150] , \labels[3][149] , 
	\labels[3][148] , \labels[3][147] , \labels[3][146] , 
	\labels[3][145] , \labels[3][144] , \labels[3][143] , 
	\labels[3][142] , \labels[3][141] , \labels[3][140] , 
	\labels[3][139] , \labels[3][138] , \labels[3][137] }, 
	_zy_simnet_labels_123_w$[0:31]);
ixc_assign_32 _zz_strnp_113 ( { \labels[3][200] , \labels[3][199] , 
	\labels[3][198] , \labels[3][197] , \labels[3][196] , 
	\labels[3][195] , \labels[3][194] , \labels[3][193] , 
	\labels[3][192] , \labels[3][191] , \labels[3][190] , 
	\labels[3][189] , \labels[3][188] , \labels[3][187] , 
	\labels[3][186] , \labels[3][185] , \labels[3][184] , 
	\labels[3][183] , \labels[3][182] , \labels[3][181] , 
	\labels[3][180] , \labels[3][179] , \labels[3][178] , 
	\labels[3][177] , \labels[3][176] , \labels[3][175] , 
	\labels[3][174] , \labels[3][173] , \labels[3][172] , 
	\labels[3][171] , \labels[3][170] , \labels[3][169] }, 
	_zy_simnet_labels_122_w$[0:31]);
ixc_assign_32 _zz_strnp_112 ( { \labels[3][232] , \labels[3][231] , 
	\labels[3][230] , \labels[3][229] , \labels[3][228] , 
	\labels[3][227] , \labels[3][226] , \labels[3][225] , 
	\labels[3][224] , \labels[3][223] , \labels[3][222] , 
	\labels[3][221] , \labels[3][220] , \labels[3][219] , 
	\labels[3][218] , \labels[3][217] , \labels[3][216] , 
	\labels[3][215] , \labels[3][214] , \labels[3][213] , 
	\labels[3][212] , \labels[3][211] , \labels[3][210] , 
	\labels[3][209] , \labels[3][208] , \labels[3][207] , 
	\labels[3][206] , \labels[3][205] , \labels[3][204] , 
	\labels[3][203] , \labels[3][202] , \labels[3][201] }, 
	_zy_simnet_labels_121_w$[0:31]);
ixc_assign_32 _zz_strnp_111 ( { \labels[3][264] , \labels[3][263] , 
	\labels[3][262] , \labels[3][261] , \labels[3][260] , 
	\labels[3][259] , \labels[3][258] , \labels[3][257] , 
	\labels[3][256] , \labels[3][255] , \labels[3][254] , 
	\labels[3][253] , \labels[3][252] , \labels[3][251] , 
	\labels[3][250] , \labels[3][249] , \labels[3][248] , 
	\labels[3][247] , \labels[3][246] , \labels[3][245] , 
	\labels[3][244] , \labels[3][243] , \labels[3][242] , 
	\labels[3][241] , \labels[3][240] , \labels[3][239] , 
	\labels[3][238] , \labels[3][237] , \labels[3][236] , 
	\labels[3][235] , \labels[3][234] , \labels[3][233] }, 
	_zy_simnet_labels_120_w$[0:31]);
ixc_assign_16 _zz_strnp_110 ( { \labels[3][271] , \labels[3][270] , 
	\labels[3][269] , \labels[3][268] , \labels[3][267] , 
	\labels[3][266] , \labels[3][265] , \labels[3][8] , \labels[3][7] , 
	\labels[3][6] , \labels[3][5] , \labels[3][4] , \labels[3][3] , 
	\labels[3][2] , \labels[3][1] , \labels[3][0] }, 
	_zy_simnet_tvar_119[0:15]);
ixc_assign_32 _zz_strnp_109 ( { \labels[2][40] , \labels[2][39] , 
	\labels[2][38] , \labels[2][37] , \labels[2][36] , \labels[2][35] , 
	\labels[2][34] , \labels[2][33] , \labels[2][32] , \labels[2][31] , 
	\labels[2][30] , \labels[2][29] , \labels[2][28] , \labels[2][27] , 
	\labels[2][26] , \labels[2][25] , \labels[2][24] , \labels[2][23] , 
	\labels[2][22] , \labels[2][21] , \labels[2][20] , \labels[2][19] , 
	\labels[2][18] , \labels[2][17] , \labels[2][16] , \labels[2][15] , 
	\labels[2][14] , \labels[2][13] , \labels[2][12] , \labels[2][11] , 
	\labels[2][10] , \labels[2][9] }, _zy_simnet_labels_118_w$[0:31]);
ixc_assign_32 _zz_strnp_108 ( { \labels[2][72] , \labels[2][71] , 
	\labels[2][70] , \labels[2][69] , \labels[2][68] , \labels[2][67] , 
	\labels[2][66] , \labels[2][65] , \labels[2][64] , \labels[2][63] , 
	\labels[2][62] , \labels[2][61] , \labels[2][60] , \labels[2][59] , 
	\labels[2][58] , \labels[2][57] , \labels[2][56] , \labels[2][55] , 
	\labels[2][54] , \labels[2][53] , \labels[2][52] , \labels[2][51] , 
	\labels[2][50] , \labels[2][49] , \labels[2][48] , \labels[2][47] , 
	\labels[2][46] , \labels[2][45] , \labels[2][44] , \labels[2][43] , 
	\labels[2][42] , \labels[2][41] }, _zy_simnet_labels_117_w$[0:31]);
ixc_assign_32 _zz_strnp_107 ( { \labels[2][104] , \labels[2][103] , 
	\labels[2][102] , \labels[2][101] , \labels[2][100] , 
	\labels[2][99] , \labels[2][98] , \labels[2][97] , \labels[2][96] , 
	\labels[2][95] , \labels[2][94] , \labels[2][93] , \labels[2][92] , 
	\labels[2][91] , \labels[2][90] , \labels[2][89] , \labels[2][88] , 
	\labels[2][87] , \labels[2][86] , \labels[2][85] , \labels[2][84] , 
	\labels[2][83] , \labels[2][82] , \labels[2][81] , \labels[2][80] , 
	\labels[2][79] , \labels[2][78] , \labels[2][77] , \labels[2][76] , 
	\labels[2][75] , \labels[2][74] , \labels[2][73] }, 
	_zy_simnet_labels_116_w$[0:31]);
ixc_assign_32 _zz_strnp_106 ( { \labels[2][136] , \labels[2][135] , 
	\labels[2][134] , \labels[2][133] , \labels[2][132] , 
	\labels[2][131] , \labels[2][130] , \labels[2][129] , 
	\labels[2][128] , \labels[2][127] , \labels[2][126] , 
	\labels[2][125] , \labels[2][124] , \labels[2][123] , 
	\labels[2][122] , \labels[2][121] , \labels[2][120] , 
	\labels[2][119] , \labels[2][118] , \labels[2][117] , 
	\labels[2][116] , \labels[2][115] , \labels[2][114] , 
	\labels[2][113] , \labels[2][112] , \labels[2][111] , 
	\labels[2][110] , \labels[2][109] , \labels[2][108] , 
	\labels[2][107] , \labels[2][106] , \labels[2][105] }, 
	_zy_simnet_labels_115_w$[0:31]);
ixc_assign_32 _zz_strnp_105 ( { \labels[2][168] , \labels[2][167] , 
	\labels[2][166] , \labels[2][165] , \labels[2][164] , 
	\labels[2][163] , \labels[2][162] , \labels[2][161] , 
	\labels[2][160] , \labels[2][159] , \labels[2][158] , 
	\labels[2][157] , \labels[2][156] , \labels[2][155] , 
	\labels[2][154] , \labels[2][153] , \labels[2][152] , 
	\labels[2][151] , \labels[2][150] , \labels[2][149] , 
	\labels[2][148] , \labels[2][147] , \labels[2][146] , 
	\labels[2][145] , \labels[2][144] , \labels[2][143] , 
	\labels[2][142] , \labels[2][141] , \labels[2][140] , 
	\labels[2][139] , \labels[2][138] , \labels[2][137] }, 
	_zy_simnet_labels_114_w$[0:31]);
ixc_assign_32 _zz_strnp_104 ( { \labels[2][200] , \labels[2][199] , 
	\labels[2][198] , \labels[2][197] , \labels[2][196] , 
	\labels[2][195] , \labels[2][194] , \labels[2][193] , 
	\labels[2][192] , \labels[2][191] , \labels[2][190] , 
	\labels[2][189] , \labels[2][188] , \labels[2][187] , 
	\labels[2][186] , \labels[2][185] , \labels[2][184] , 
	\labels[2][183] , \labels[2][182] , \labels[2][181] , 
	\labels[2][180] , \labels[2][179] , \labels[2][178] , 
	\labels[2][177] , \labels[2][176] , \labels[2][175] , 
	\labels[2][174] , \labels[2][173] , \labels[2][172] , 
	\labels[2][171] , \labels[2][170] , \labels[2][169] }, 
	_zy_simnet_labels_113_w$[0:31]);
ixc_assign_32 _zz_strnp_103 ( { \labels[2][232] , \labels[2][231] , 
	\labels[2][230] , \labels[2][229] , \labels[2][228] , 
	\labels[2][227] , \labels[2][226] , \labels[2][225] , 
	\labels[2][224] , \labels[2][223] , \labels[2][222] , 
	\labels[2][221] , \labels[2][220] , \labels[2][219] , 
	\labels[2][218] , \labels[2][217] , \labels[2][216] , 
	\labels[2][215] , \labels[2][214] , \labels[2][213] , 
	\labels[2][212] , \labels[2][211] , \labels[2][210] , 
	\labels[2][209] , \labels[2][208] , \labels[2][207] , 
	\labels[2][206] , \labels[2][205] , \labels[2][204] , 
	\labels[2][203] , \labels[2][202] , \labels[2][201] }, 
	_zy_simnet_labels_112_w$[0:31]);
ixc_assign_32 _zz_strnp_102 ( { \labels[2][264] , \labels[2][263] , 
	\labels[2][262] , \labels[2][261] , \labels[2][260] , 
	\labels[2][259] , \labels[2][258] , \labels[2][257] , 
	\labels[2][256] , \labels[2][255] , \labels[2][254] , 
	\labels[2][253] , \labels[2][252] , \labels[2][251] , 
	\labels[2][250] , \labels[2][249] , \labels[2][248] , 
	\labels[2][247] , \labels[2][246] , \labels[2][245] , 
	\labels[2][244] , \labels[2][243] , \labels[2][242] , 
	\labels[2][241] , \labels[2][240] , \labels[2][239] , 
	\labels[2][238] , \labels[2][237] , \labels[2][236] , 
	\labels[2][235] , \labels[2][234] , \labels[2][233] }, 
	_zy_simnet_labels_111_w$[0:31]);
ixc_assign_16 _zz_strnp_101 ( { \labels[2][271] , \labels[2][270] , 
	\labels[2][269] , \labels[2][268] , \labels[2][267] , 
	\labels[2][266] , \labels[2][265] , \labels[2][8] , \labels[2][7] , 
	\labels[2][6] , \labels[2][5] , \labels[2][4] , \labels[2][3] , 
	\labels[2][2] , \labels[2][1] , \labels[2][0] }, 
	_zy_simnet_tvar_110[0:15]);
ixc_assign_32 _zz_strnp_100 ( { \labels[1][40] , \labels[1][39] , 
	\labels[1][38] , \labels[1][37] , \labels[1][36] , \labels[1][35] , 
	\labels[1][34] , \labels[1][33] , \labels[1][32] , \labels[1][31] , 
	\labels[1][30] , \labels[1][29] , \labels[1][28] , \labels[1][27] , 
	\labels[1][26] , \labels[1][25] , \labels[1][24] , \labels[1][23] , 
	\labels[1][22] , \labels[1][21] , \labels[1][20] , \labels[1][19] , 
	\labels[1][18] , \labels[1][17] , \labels[1][16] , \labels[1][15] , 
	\labels[1][14] , \labels[1][13] , \labels[1][12] , \labels[1][11] , 
	\labels[1][10] , \labels[1][9] }, _zy_simnet_labels_109_w$[0:31]);
ixc_assign_32 _zz_strnp_99 ( { \labels[1][72] , \labels[1][71] , 
	\labels[1][70] , \labels[1][69] , \labels[1][68] , \labels[1][67] , 
	\labels[1][66] , \labels[1][65] , \labels[1][64] , \labels[1][63] , 
	\labels[1][62] , \labels[1][61] , \labels[1][60] , \labels[1][59] , 
	\labels[1][58] , \labels[1][57] , \labels[1][56] , \labels[1][55] , 
	\labels[1][54] , \labels[1][53] , \labels[1][52] , \labels[1][51] , 
	\labels[1][50] , \labels[1][49] , \labels[1][48] , \labels[1][47] , 
	\labels[1][46] , \labels[1][45] , \labels[1][44] , \labels[1][43] , 
	\labels[1][42] , \labels[1][41] }, _zy_simnet_labels_108_w$[0:31]);
ixc_assign_32 _zz_strnp_98 ( { \labels[1][104] , \labels[1][103] , 
	\labels[1][102] , \labels[1][101] , \labels[1][100] , 
	\labels[1][99] , \labels[1][98] , \labels[1][97] , \labels[1][96] , 
	\labels[1][95] , \labels[1][94] , \labels[1][93] , \labels[1][92] , 
	\labels[1][91] , \labels[1][90] , \labels[1][89] , \labels[1][88] , 
	\labels[1][87] , \labels[1][86] , \labels[1][85] , \labels[1][84] , 
	\labels[1][83] , \labels[1][82] , \labels[1][81] , \labels[1][80] , 
	\labels[1][79] , \labels[1][78] , \labels[1][77] , \labels[1][76] , 
	\labels[1][75] , \labels[1][74] , \labels[1][73] }, 
	_zy_simnet_labels_107_w$[0:31]);
ixc_assign_32 _zz_strnp_97 ( { \labels[1][136] , \labels[1][135] , 
	\labels[1][134] , \labels[1][133] , \labels[1][132] , 
	\labels[1][131] , \labels[1][130] , \labels[1][129] , 
	\labels[1][128] , \labels[1][127] , \labels[1][126] , 
	\labels[1][125] , \labels[1][124] , \labels[1][123] , 
	\labels[1][122] , \labels[1][121] , \labels[1][120] , 
	\labels[1][119] , \labels[1][118] , \labels[1][117] , 
	\labels[1][116] , \labels[1][115] , \labels[1][114] , 
	\labels[1][113] , \labels[1][112] , \labels[1][111] , 
	\labels[1][110] , \labels[1][109] , \labels[1][108] , 
	\labels[1][107] , \labels[1][106] , \labels[1][105] }, 
	_zy_simnet_labels_106_w$[0:31]);
ixc_assign_32 _zz_strnp_96 ( { \labels[1][168] , \labels[1][167] , 
	\labels[1][166] , \labels[1][165] , \labels[1][164] , 
	\labels[1][163] , \labels[1][162] , \labels[1][161] , 
	\labels[1][160] , \labels[1][159] , \labels[1][158] , 
	\labels[1][157] , \labels[1][156] , \labels[1][155] , 
	\labels[1][154] , \labels[1][153] , \labels[1][152] , 
	\labels[1][151] , \labels[1][150] , \labels[1][149] , 
	\labels[1][148] , \labels[1][147] , \labels[1][146] , 
	\labels[1][145] , \labels[1][144] , \labels[1][143] , 
	\labels[1][142] , \labels[1][141] , \labels[1][140] , 
	\labels[1][139] , \labels[1][138] , \labels[1][137] }, 
	_zy_simnet_labels_105_w$[0:31]);
ixc_assign_32 _zz_strnp_95 ( { \labels[1][200] , \labels[1][199] , 
	\labels[1][198] , \labels[1][197] , \labels[1][196] , 
	\labels[1][195] , \labels[1][194] , \labels[1][193] , 
	\labels[1][192] , \labels[1][191] , \labels[1][190] , 
	\labels[1][189] , \labels[1][188] , \labels[1][187] , 
	\labels[1][186] , \labels[1][185] , \labels[1][184] , 
	\labels[1][183] , \labels[1][182] , \labels[1][181] , 
	\labels[1][180] , \labels[1][179] , \labels[1][178] , 
	\labels[1][177] , \labels[1][176] , \labels[1][175] , 
	\labels[1][174] , \labels[1][173] , \labels[1][172] , 
	\labels[1][171] , \labels[1][170] , \labels[1][169] }, 
	_zy_simnet_labels_104_w$[0:31]);
ixc_assign_32 _zz_strnp_94 ( { \labels[1][232] , \labels[1][231] , 
	\labels[1][230] , \labels[1][229] , \labels[1][228] , 
	\labels[1][227] , \labels[1][226] , \labels[1][225] , 
	\labels[1][224] , \labels[1][223] , \labels[1][222] , 
	\labels[1][221] , \labels[1][220] , \labels[1][219] , 
	\labels[1][218] , \labels[1][217] , \labels[1][216] , 
	\labels[1][215] , \labels[1][214] , \labels[1][213] , 
	\labels[1][212] , \labels[1][211] , \labels[1][210] , 
	\labels[1][209] , \labels[1][208] , \labels[1][207] , 
	\labels[1][206] , \labels[1][205] , \labels[1][204] , 
	\labels[1][203] , \labels[1][202] , \labels[1][201] }, 
	_zy_simnet_labels_103_w$[0:31]);
ixc_assign_32 _zz_strnp_93 ( { \labels[1][264] , \labels[1][263] , 
	\labels[1][262] , \labels[1][261] , \labels[1][260] , 
	\labels[1][259] , \labels[1][258] , \labels[1][257] , 
	\labels[1][256] , \labels[1][255] , \labels[1][254] , 
	\labels[1][253] , \labels[1][252] , \labels[1][251] , 
	\labels[1][250] , \labels[1][249] , \labels[1][248] , 
	\labels[1][247] , \labels[1][246] , \labels[1][245] , 
	\labels[1][244] , \labels[1][243] , \labels[1][242] , 
	\labels[1][241] , \labels[1][240] , \labels[1][239] , 
	\labels[1][238] , \labels[1][237] , \labels[1][236] , 
	\labels[1][235] , \labels[1][234] , \labels[1][233] }, 
	_zy_simnet_labels_102_w$[0:31]);
ixc_assign_16 _zz_strnp_92 ( { \labels[1][271] , \labels[1][270] , 
	\labels[1][269] , \labels[1][268] , \labels[1][267] , 
	\labels[1][266] , \labels[1][265] , \labels[1][8] , \labels[1][7] , 
	\labels[1][6] , \labels[1][5] , \labels[1][4] , \labels[1][3] , 
	\labels[1][2] , \labels[1][1] , \labels[1][0] }, 
	_zy_simnet_tvar_101[0:15]);
ixc_assign_32 _zz_strnp_91 ( { \labels[0][40] , \labels[0][39] , 
	\labels[0][38] , \labels[0][37] , \labels[0][36] , \labels[0][35] , 
	\labels[0][34] , \labels[0][33] , \labels[0][32] , \labels[0][31] , 
	\labels[0][30] , \labels[0][29] , \labels[0][28] , \labels[0][27] , 
	\labels[0][26] , \labels[0][25] , \labels[0][24] , \labels[0][23] , 
	\labels[0][22] , \labels[0][21] , \labels[0][20] , \labels[0][19] , 
	\labels[0][18] , \labels[0][17] , \labels[0][16] , \labels[0][15] , 
	\labels[0][14] , \labels[0][13] , \labels[0][12] , \labels[0][11] , 
	\labels[0][10] , \labels[0][9] }, _zy_simnet_labels_100_w$[0:31]);
ixc_assign_32 _zz_strnp_90 ( { \labels[0][72] , \labels[0][71] , 
	\labels[0][70] , \labels[0][69] , \labels[0][68] , \labels[0][67] , 
	\labels[0][66] , \labels[0][65] , \labels[0][64] , \labels[0][63] , 
	\labels[0][62] , \labels[0][61] , \labels[0][60] , \labels[0][59] , 
	\labels[0][58] , \labels[0][57] , \labels[0][56] , \labels[0][55] , 
	\labels[0][54] , \labels[0][53] , \labels[0][52] , \labels[0][51] , 
	\labels[0][50] , \labels[0][49] , \labels[0][48] , \labels[0][47] , 
	\labels[0][46] , \labels[0][45] , \labels[0][44] , \labels[0][43] , 
	\labels[0][42] , \labels[0][41] }, _zy_simnet_labels_99_w$[0:31]);
ixc_assign_32 _zz_strnp_89 ( { \labels[0][104] , \labels[0][103] , 
	\labels[0][102] , \labels[0][101] , \labels[0][100] , 
	\labels[0][99] , \labels[0][98] , \labels[0][97] , \labels[0][96] , 
	\labels[0][95] , \labels[0][94] , \labels[0][93] , \labels[0][92] , 
	\labels[0][91] , \labels[0][90] , \labels[0][89] , \labels[0][88] , 
	\labels[0][87] , \labels[0][86] , \labels[0][85] , \labels[0][84] , 
	\labels[0][83] , \labels[0][82] , \labels[0][81] , \labels[0][80] , 
	\labels[0][79] , \labels[0][78] , \labels[0][77] , \labels[0][76] , 
	\labels[0][75] , \labels[0][74] , \labels[0][73] }, 
	_zy_simnet_labels_98_w$[0:31]);
ixc_assign_32 _zz_strnp_88 ( { \labels[0][136] , \labels[0][135] , 
	\labels[0][134] , \labels[0][133] , \labels[0][132] , 
	\labels[0][131] , \labels[0][130] , \labels[0][129] , 
	\labels[0][128] , \labels[0][127] , \labels[0][126] , 
	\labels[0][125] , \labels[0][124] , \labels[0][123] , 
	\labels[0][122] , \labels[0][121] , \labels[0][120] , 
	\labels[0][119] , \labels[0][118] , \labels[0][117] , 
	\labels[0][116] , \labels[0][115] , \labels[0][114] , 
	\labels[0][113] , \labels[0][112] , \labels[0][111] , 
	\labels[0][110] , \labels[0][109] , \labels[0][108] , 
	\labels[0][107] , \labels[0][106] , \labels[0][105] }, 
	_zy_simnet_labels_97_w$[0:31]);
ixc_assign_32 _zz_strnp_87 ( { \labels[0][168] , \labels[0][167] , 
	\labels[0][166] , \labels[0][165] , \labels[0][164] , 
	\labels[0][163] , \labels[0][162] , \labels[0][161] , 
	\labels[0][160] , \labels[0][159] , \labels[0][158] , 
	\labels[0][157] , \labels[0][156] , \labels[0][155] , 
	\labels[0][154] , \labels[0][153] , \labels[0][152] , 
	\labels[0][151] , \labels[0][150] , \labels[0][149] , 
	\labels[0][148] , \labels[0][147] , \labels[0][146] , 
	\labels[0][145] , \labels[0][144] , \labels[0][143] , 
	\labels[0][142] , \labels[0][141] , \labels[0][140] , 
	\labels[0][139] , \labels[0][138] , \labels[0][137] }, 
	_zy_simnet_labels_96_w$[0:31]);
ixc_assign_32 _zz_strnp_86 ( { \labels[0][200] , \labels[0][199] , 
	\labels[0][198] , \labels[0][197] , \labels[0][196] , 
	\labels[0][195] , \labels[0][194] , \labels[0][193] , 
	\labels[0][192] , \labels[0][191] , \labels[0][190] , 
	\labels[0][189] , \labels[0][188] , \labels[0][187] , 
	\labels[0][186] , \labels[0][185] , \labels[0][184] , 
	\labels[0][183] , \labels[0][182] , \labels[0][181] , 
	\labels[0][180] , \labels[0][179] , \labels[0][178] , 
	\labels[0][177] , \labels[0][176] , \labels[0][175] , 
	\labels[0][174] , \labels[0][173] , \labels[0][172] , 
	\labels[0][171] , \labels[0][170] , \labels[0][169] }, 
	_zy_simnet_labels_95_w$[0:31]);
ixc_assign_32 _zz_strnp_85 ( { \labels[0][232] , \labels[0][231] , 
	\labels[0][230] , \labels[0][229] , \labels[0][228] , 
	\labels[0][227] , \labels[0][226] , \labels[0][225] , 
	\labels[0][224] , \labels[0][223] , \labels[0][222] , 
	\labels[0][221] , \labels[0][220] , \labels[0][219] , 
	\labels[0][218] , \labels[0][217] , \labels[0][216] , 
	\labels[0][215] , \labels[0][214] , \labels[0][213] , 
	\labels[0][212] , \labels[0][211] , \labels[0][210] , 
	\labels[0][209] , \labels[0][208] , \labels[0][207] , 
	\labels[0][206] , \labels[0][205] , \labels[0][204] , 
	\labels[0][203] , \labels[0][202] , \labels[0][201] }, 
	_zy_simnet_labels_94_w$[0:31]);
ixc_assign_32 _zz_strnp_84 ( { \labels[0][264] , \labels[0][263] , 
	\labels[0][262] , \labels[0][261] , \labels[0][260] , 
	\labels[0][259] , \labels[0][258] , \labels[0][257] , 
	\labels[0][256] , \labels[0][255] , \labels[0][254] , 
	\labels[0][253] , \labels[0][252] , \labels[0][251] , 
	\labels[0][250] , \labels[0][249] , \labels[0][248] , 
	\labels[0][247] , \labels[0][246] , \labels[0][245] , 
	\labels[0][244] , \labels[0][243] , \labels[0][242] , 
	\labels[0][241] , \labels[0][240] , \labels[0][239] , 
	\labels[0][238] , \labels[0][237] , \labels[0][236] , 
	\labels[0][235] , \labels[0][234] , \labels[0][233] }, 
	_zy_simnet_labels_93_w$[0:31]);
ixc_assign_16 _zz_strnp_83 ( { \labels[0][271] , \labels[0][270] , 
	\labels[0][269] , \labels[0][268] , \labels[0][267] , 
	\labels[0][266] , \labels[0][265] , \labels[0][8] , \labels[0][7] , 
	\labels[0][6] , \labels[0][5] , \labels[0][4] , \labels[0][3] , 
	\labels[0][2] , \labels[0][1] , \labels[0][0] }, 
	_zy_simnet_tvar_92[0:15]);
ixc_assign_18 _zz_strnp_82 ( o_kim_ia_config[17:0], 
	_zy_simnet_o_kim_ia_config_91_w$[0:17]);
ixc_assign_17 _zz_strnp_81 ( o_kim_ia_wdata_part1[16:0], 
	_zy_simnet_o_kim_ia_wdata_part1_90_w$[0:16]);
ixc_assign_21 _zz_strnp_80 ( o_kim_ia_wdata_part0[20:0], 
	_zy_simnet_o_kim_ia_wdata_part0_89_w$[0:20]);
ixc_assign_19 _zz_strnp_79 ( o_ckv_ia_config[18:0], 
	_zy_simnet_o_ckv_ia_config_88_w$[0:18]);
ixc_assign_32 _zz_strnp_78 ( o_ckv_ia_wdata_part1[31:0], 
	_zy_simnet_o_ckv_ia_wdata_part1_87_w$[0:31]);
ixc_assign_32 _zz_strnp_77 ( o_ckv_ia_wdata_part0[31:0], 
	_zy_simnet_o_ckv_ia_wdata_part0_86_w$[0:31]);
ixc_assign_12 _zz_strnp_76 ( cddip3_out_im_config[11:0], 
	_zy_simnet_cddip3_out_im_config_84_w$[0:11]);
ixc_assign_13 _zz_strnp_75 ( cddip3_out_ia_config[12:0], 
	_zy_simnet_cddip3_out_ia_config_83_w$[0:12]);
ixc_assign_32 _zz_strnp_74 ( cddip3_out_ia_wdata[95:64], 
	_zy_simnet_cddip3_out_ia_wdata_82_w$[0:31]);
ixc_assign_32 _zz_strnp_73 ( cddip3_out_ia_wdata[63:32], 
	_zy_simnet_cddip3_out_ia_wdata_81_w$[0:31]);
ixc_assign_32 _zz_strnp_72 ( cddip3_out_ia_wdata[31:0], 
	_zy_simnet_cddip3_out_ia_wdata_80_w$[0:31]);
ixc_assign_12 _zz_strnp_71 ( cddip2_out_im_config[11:0], 
	_zy_simnet_cddip2_out_im_config_78_w$[0:11]);
ixc_assign_13 _zz_strnp_70 ( cddip2_out_ia_config[12:0], 
	_zy_simnet_cddip2_out_ia_config_77_w$[0:12]);
ixc_assign_32 _zz_strnp_69 ( cddip2_out_ia_wdata[95:64], 
	_zy_simnet_cddip2_out_ia_wdata_76_w$[0:31]);
ixc_assign_32 _zz_strnp_68 ( cddip2_out_ia_wdata[63:32], 
	_zy_simnet_cddip2_out_ia_wdata_75_w$[0:31]);
ixc_assign_32 _zz_strnp_67 ( cddip2_out_ia_wdata[31:0], 
	_zy_simnet_cddip2_out_ia_wdata_74_w$[0:31]);
ixc_assign_12 _zz_strnp_66 ( cddip1_out_im_config[11:0], 
	_zy_simnet_cddip1_out_im_config_72_w$[0:11]);
ixc_assign_13 _zz_strnp_65 ( cddip1_out_ia_config[12:0], 
	_zy_simnet_cddip1_out_ia_config_71_w$[0:12]);
ixc_assign_32 _zz_strnp_64 ( cddip1_out_ia_wdata[95:64], 
	_zy_simnet_cddip1_out_ia_wdata_70_w$[0:31]);
ixc_assign_32 _zz_strnp_63 ( cddip1_out_ia_wdata[63:32], 
	_zy_simnet_cddip1_out_ia_wdata_69_w$[0:31]);
ixc_assign_32 _zz_strnp_62 ( cddip1_out_ia_wdata[31:0], 
	_zy_simnet_cddip1_out_ia_wdata_68_w$[0:31]);
ixc_assign_12 _zz_strnp_61 ( cddip0_out_im_config[11:0], 
	_zy_simnet_cddip0_out_im_config_66_w$[0:11]);
ixc_assign_13 _zz_strnp_60 ( cddip0_out_ia_config[12:0], 
	_zy_simnet_cddip0_out_ia_config_65_w$[0:12]);
ixc_assign_32 _zz_strnp_59 ( cddip0_out_ia_wdata[95:64], 
	_zy_simnet_cddip0_out_ia_wdata_64_w$[0:31]);
ixc_assign_32 _zz_strnp_58 ( cddip0_out_ia_wdata[63:32], 
	_zy_simnet_cddip0_out_ia_wdata_63_w$[0:31]);
ixc_assign_32 _zz_strnp_57 ( cddip0_out_ia_wdata[31:0], 
	_zy_simnet_cddip0_out_ia_wdata_62_w$[0:31]);
ixc_assign_12 _zz_strnp_56 ( cceip3_out_im_config[11:0], 
	_zy_simnet_cceip3_out_im_config_60_w$[0:11]);
ixc_assign_13 _zz_strnp_55 ( cceip3_out_ia_config[12:0], 
	_zy_simnet_cceip3_out_ia_config_59_w$[0:12]);
ixc_assign_32 _zz_strnp_54 ( cceip3_out_ia_wdata[95:64], 
	_zy_simnet_cceip3_out_ia_wdata_58_w$[0:31]);
ixc_assign_32 _zz_strnp_53 ( cceip3_out_ia_wdata[63:32], 
	_zy_simnet_cceip3_out_ia_wdata_57_w$[0:31]);
ixc_assign_32 _zz_strnp_52 ( cceip3_out_ia_wdata[31:0], 
	_zy_simnet_cceip3_out_ia_wdata_56_w$[0:31]);
ixc_assign_12 _zz_strnp_51 ( cceip2_out_im_config[11:0], 
	_zy_simnet_cceip2_out_im_config_54_w$[0:11]);
ixc_assign_13 _zz_strnp_50 ( cceip2_out_ia_config[12:0], 
	_zy_simnet_cceip2_out_ia_config_53_w$[0:12]);
ixc_assign_32 _zz_strnp_49 ( cceip2_out_ia_wdata[95:64], 
	_zy_simnet_cceip2_out_ia_wdata_52_w$[0:31]);
ixc_assign_32 _zz_strnp_48 ( cceip2_out_ia_wdata[63:32], 
	_zy_simnet_cceip2_out_ia_wdata_51_w$[0:31]);
ixc_assign_32 _zz_strnp_47 ( cceip2_out_ia_wdata[31:0], 
	_zy_simnet_cceip2_out_ia_wdata_50_w$[0:31]);
ixc_assign_12 _zz_strnp_46 ( cceip1_out_im_config[11:0], 
	_zy_simnet_cceip1_out_im_config_48_w$[0:11]);
ixc_assign_13 _zz_strnp_45 ( cceip1_out_ia_config[12:0], 
	_zy_simnet_cceip1_out_ia_config_47_w$[0:12]);
ixc_assign_32 _zz_strnp_44 ( cceip1_out_ia_wdata[95:64], 
	_zy_simnet_cceip1_out_ia_wdata_46_w$[0:31]);
ixc_assign_32 _zz_strnp_43 ( cceip1_out_ia_wdata[63:32], 
	_zy_simnet_cceip1_out_ia_wdata_45_w$[0:31]);
ixc_assign_32 _zz_strnp_42 ( cceip1_out_ia_wdata[31:0], 
	_zy_simnet_cceip1_out_ia_wdata_44_w$[0:31]);
ixc_assign_12 _zz_strnp_41 ( cceip0_out_im_config[11:0], 
	_zy_simnet_cceip0_out_im_config_42_w$[0:11]);
ixc_assign_13 _zz_strnp_40 ( cceip0_out_ia_config[12:0], 
	_zy_simnet_cceip0_out_ia_config_41_w$[0:12]);
ixc_assign_32 _zz_strnp_39 ( cceip0_out_ia_wdata[95:64], 
	_zy_simnet_cceip0_out_ia_wdata_40_w$[0:31]);
ixc_assign_32 _zz_strnp_38 ( cceip0_out_ia_wdata[63:32], 
	_zy_simnet_cceip0_out_ia_wdata_39_w$[0:31]);
ixc_assign_32 _zz_strnp_37 ( cceip0_out_ia_wdata[31:0], 
	_zy_simnet_cceip0_out_ia_wdata_38_w$[0:31]);
ixc_assign_32 _zz_strnp_36 ( { _zy_simnet_tvar_33[0], _zy_simnet_tvar_33[1], 
	_zy_simnet_tvar_33[2], _zy_simnet_tvar_33[3], _zy_simnet_tvar_33[4], 
	_zy_simnet_tvar_33[5], _zy_simnet_tvar_33[6], _zy_simnet_tvar_33[7], 
	_zy_simnet_tvar_33[8], _zy_simnet_tvar_33[9], _zy_simnet_tvar_33[10], 
	_zy_simnet_tvar_33[11], _zy_simnet_tvar_33[12], 
	_zy_simnet_tvar_33[13], _zy_simnet_tvar_33[14], 
	_zy_simnet_tvar_33[15], _zy_simnet_tvar_33[16], 
	_zy_simnet_tvar_33[17], _zy_simnet_tvar_33[18], 
	_zy_simnet_tvar_33[19], _zy_simnet_tvar_33[20], 
	_zy_simnet_tvar_33[21], _zy_simnet_tvar_33[22], 
	_zy_simnet_tvar_33[23], _zy_simnet_tvar_33[24], kdf_test_mode_en, 
	always_validate_kim_ref, manual_txc, _zy_simnet_tvar_34, 
	_zy_simnet_tvar_35, _zy_simnet_tvar_36, _zy_simnet_tvar_37}, 
	_zy_simnet_tvar_32[0:31]);
ixc_assign _zz_strnp_30 ( locl_err_ack, _zy_simnet_locl_err_ack_31_w$);
ixc_assign _zz_strnp_29 ( locl_ack, _zy_simnet_locl_ack_30_w$);
ixc_assign_32 _zz_strnp_28 ( locl_rd_data[31:0], 
	_zy_simnet_locl_rd_data_29_w$[0:31]);
ixc_assign _zz_strnp_27 ( _zy_simnet_locl_rd_strb_28_w$, locl_rd_strb);
ixc_assign_32 _zz_strnp_26 ( _zy_simnet_locl_wr_data_27_w$[0:31], 
	locl_wr_data[31:0]);
ixc_assign _zz_strnp_25 ( _zy_simnet_locl_wr_strb_26_w$, locl_wr_strb);
ixc_assign_11 _zz_strnp_24 ( _zy_simnet_locl_addr_25_w$[0:10], 
	locl_addr[10:0]);
ixc_assign_32 _zz_strnp_23 ( _zy_simnet_sa_global_ctrl_23_w$[0:31], 
	sa_global_ctrl[31:0]);
ixc_assign_7 _zz_strnp_22 ( 
	_zy_simnet_cddip_decrypt_kop_fifo_override_22_w$[0:6], 
	cddip_decrypt_kop_fifo_override[6:0]);
ixc_assign_7 _zz_strnp_21 ( 
	_zy_simnet_cceip_validate_kop_fifo_override_21_w$[0:6], 
	cceip_validate_kop_fifo_override[6:0]);
ixc_assign_7 _zz_strnp_20 ( 
	_zy_simnet_cceip_encrypt_kop_fifo_override_20_w$[0:6], 
	cceip_encrypt_kop_fifo_override[6:0]);
ixc_assign_9 _zz_strnp_19 ( _zy_simnet_tready_override_19_w$[0:8], 
	tready_override[8:0]);
ixc_assign_2176 _zz_strnp_18 ( _zy_simnet_labels_18_w$[0:2175], { 
	\labels[7][271] , \labels[7][270] , \labels[7][269] , 
	\labels[7][268] , \labels[7][267] , \labels[7][266] , 
	\labels[7][265] , \labels[7][264] , \labels[7][263] , 
	\labels[7][262] , \labels[7][261] , \labels[7][260] , 
	\labels[7][259] , \labels[7][258] , \labels[7][257] , 
	\labels[7][256] , \labels[7][255] , \labels[7][254] , 
	\labels[7][253] , \labels[7][252] , \labels[7][251] , 
	\labels[7][250] , \labels[7][249] , \labels[7][248] , 
	\labels[7][247] , \labels[7][246] , \labels[7][245] , 
	\labels[7][244] , \labels[7][243] , \labels[7][242] , 
	\labels[7][241] , \labels[7][240] , \labels[7][239] , 
	\labels[7][238] , \labels[7][237] , \labels[7][236] , 
	\labels[7][235] , \labels[7][234] , \labels[7][233] , 
	\labels[7][232] , \labels[7][231] , \labels[7][230] , 
	\labels[7][229] , \labels[7][228] , \labels[7][227] , 
	\labels[7][226] , \labels[7][225] , \labels[7][224] , 
	\labels[7][223] , \labels[7][222] , \labels[7][221] , 
	\labels[7][220] , \labels[7][219] , \labels[7][218] , 
	\labels[7][217] , \labels[7][216] , \labels[7][215] , 
	\labels[7][214] , \labels[7][213] , \labels[7][212] , 
	\labels[7][211] , \labels[7][210] , \labels[7][209] , 
	\labels[7][208] , \labels[7][207] , \labels[7][206] , 
	\labels[7][205] , \labels[7][204] , \labels[7][203] , 
	\labels[7][202] , \labels[7][201] , \labels[7][200] , 
	\labels[7][199] , \labels[7][198] , \labels[7][197] , 
	\labels[7][196] , \labels[7][195] , \labels[7][194] , 
	\labels[7][193] , \labels[7][192] , \labels[7][191] , 
	\labels[7][190] , \labels[7][189] , \labels[7][188] , 
	\labels[7][187] , \labels[7][186] , \labels[7][185] , 
	\labels[7][184] , \labels[7][183] , \labels[7][182] , 
	\labels[7][181] , \labels[7][180] , \labels[7][179] , 
	\labels[7][178] , \labels[7][177] , \labels[7][176] , 
	\labels[7][175] , \labels[7][174] , \labels[7][173] , 
	\labels[7][172] , \labels[7][171] , \labels[7][170] , 
	\labels[7][169] , \labels[7][168] , \labels[7][167] , 
	\labels[7][166] , \labels[7][165] , \labels[7][164] , 
	\labels[7][163] , \labels[7][162] , \labels[7][161] , 
	\labels[7][160] , \labels[7][159] , \labels[7][158] , 
	\labels[7][157] , \labels[7][156] , \labels[7][155] , 
	\labels[7][154] , \labels[7][153] , \labels[7][152] , 
	\labels[7][151] , \labels[7][150] , \labels[7][149] , 
	\labels[7][148] , \labels[7][147] , \labels[7][146] , 
	\labels[7][145] , \labels[7][144] , \labels[7][143] , 
	\labels[7][142] , \labels[7][141] , \labels[7][140] , 
	\labels[7][139] , \labels[7][138] , \labels[7][137] , 
	\labels[7][136] , \labels[7][135] , \labels[7][134] , 
	\labels[7][133] , \labels[7][132] , \labels[7][131] , 
	\labels[7][130] , \labels[7][129] , \labels[7][128] , 
	\labels[7][127] , \labels[7][126] , \labels[7][125] , 
	\labels[7][124] , \labels[7][123] , \labels[7][122] , 
	\labels[7][121] , \labels[7][120] , \labels[7][119] , 
	\labels[7][118] , \labels[7][117] , \labels[7][116] , 
	\labels[7][115] , \labels[7][114] , \labels[7][113] , 
	\labels[7][112] , \labels[7][111] , \labels[7][110] , 
	\labels[7][109] , \labels[7][108] , \labels[7][107] , 
	\labels[7][106] , \labels[7][105] , \labels[7][104] , 
	\labels[7][103] , \labels[7][102] , \labels[7][101] , 
	\labels[7][100] , \labels[7][99] , \labels[7][98] , \labels[7][97] , 
	\labels[7][96] , \labels[7][95] , \labels[7][94] , \labels[7][93] , 
	\labels[7][92] , \labels[7][91] , \labels[7][90] , \labels[7][89] , 
	\labels[7][88] , \labels[7][87] , \labels[7][86] , \labels[7][85] , 
	\labels[7][84] , \labels[7][83] , \labels[7][82] , \labels[7][81] , 
	\labels[7][80] , \labels[7][79] , \labels[7][78] , \labels[7][77] , 
	\labels[7][76] , \labels[7][75] , \labels[7][74] , \labels[7][73] , 
	\labels[7][72] , \labels[7][71] , \labels[7][70] , \labels[7][69] , 
	\labels[7][68] , \labels[7][67] , \labels[7][66] , \labels[7][65] , 
	\labels[7][64] , \labels[7][63] , \labels[7][62] , \labels[7][61] , 
	\labels[7][60] , \labels[7][59] , \labels[7][58] , \labels[7][57] , 
	\labels[7][56] , \labels[7][55] , \labels[7][54] , \labels[7][53] , 
	\labels[7][52] , \labels[7][51] , \labels[7][50] , \labels[7][49] , 
	\labels[7][48] , \labels[7][47] , \labels[7][46] , \labels[7][45] , 
	\labels[7][44] , \labels[7][43] , \labels[7][42] , \labels[7][41] , 
	\labels[7][40] , \labels[7][39] , \labels[7][38] , \labels[7][37] , 
	\labels[7][36] , \labels[7][35] , \labels[7][34] , \labels[7][33] , 
	\labels[7][32] , \labels[7][31] , \labels[7][30] , \labels[7][29] , 
	\labels[7][28] , \labels[7][27] , \labels[7][26] , \labels[7][25] , 
	\labels[7][24] , \labels[7][23] , \labels[7][22] , \labels[7][21] , 
	\labels[7][20] , \labels[7][19] , \labels[7][18] , \labels[7][17] , 
	\labels[7][16] , \labels[7][15] , \labels[7][14] , \labels[7][13] , 
	\labels[7][12] , \labels[7][11] , \labels[7][10] , \labels[7][9] , 
	\labels[7][8] , \labels[7][7] , \labels[7][6] , \labels[7][5] , 
	\labels[7][4] , \labels[7][3] , \labels[7][2] , \labels[7][1] , 
	\labels[7][0] , \labels[6][271] , \labels[6][270] , \labels[6][269] , 
	\labels[6][268] , \labels[6][267] , \labels[6][266] , 
	\labels[6][265] , \labels[6][264] , \labels[6][263] , 
	\labels[6][262] , \labels[6][261] , \labels[6][260] , 
	\labels[6][259] , \labels[6][258] , \labels[6][257] , 
	\labels[6][256] , \labels[6][255] , \labels[6][254] , 
	\labels[6][253] , \labels[6][252] , \labels[6][251] , 
	\labels[6][250] , \labels[6][249] , \labels[6][248] , 
	\labels[6][247] , \labels[6][246] , \labels[6][245] , 
	\labels[6][244] , \labels[6][243] , \labels[6][242] , 
	\labels[6][241] , \labels[6][240] , \labels[6][239] , 
	\labels[6][238] , \labels[6][237] , \labels[6][236] , 
	\labels[6][235] , \labels[6][234] , \labels[6][233] , 
	\labels[6][232] , \labels[6][231] , \labels[6][230] , 
	\labels[6][229] , \labels[6][228] , \labels[6][227] , 
	\labels[6][226] , \labels[6][225] , \labels[6][224] , 
	\labels[6][223] , \labels[6][222] , \labels[6][221] , 
	\labels[6][220] , \labels[6][219] , \labels[6][218] , 
	\labels[6][217] , \labels[6][216] , \labels[6][215] , 
	\labels[6][214] , \labels[6][213] , \labels[6][212] , 
	\labels[6][211] , \labels[6][210] , \labels[6][209] , 
	\labels[6][208] , \labels[6][207] , \labels[6][206] , 
	\labels[6][205] , \labels[6][204] , \labels[6][203] , 
	\labels[6][202] , \labels[6][201] , \labels[6][200] , 
	\labels[6][199] , \labels[6][198] , \labels[6][197] , 
	\labels[6][196] , \labels[6][195] , \labels[6][194] , 
	\labels[6][193] , \labels[6][192] , \labels[6][191] , 
	\labels[6][190] , \labels[6][189] , \labels[6][188] , 
	\labels[6][187] , \labels[6][186] , \labels[6][185] , 
	\labels[6][184] , \labels[6][183] , \labels[6][182] , 
	\labels[6][181] , \labels[6][180] , \labels[6][179] , 
	\labels[6][178] , \labels[6][177] , \labels[6][176] , 
	\labels[6][175] , \labels[6][174] , \labels[6][173] , 
	\labels[6][172] , \labels[6][171] , \labels[6][170] , 
	\labels[6][169] , \labels[6][168] , \labels[6][167] , 
	\labels[6][166] , \labels[6][165] , \labels[6][164] , 
	\labels[6][163] , \labels[6][162] , \labels[6][161] , 
	\labels[6][160] , \labels[6][159] , \labels[6][158] , 
	\labels[6][157] , \labels[6][156] , \labels[6][155] , 
	\labels[6][154] , \labels[6][153] , \labels[6][152] , 
	\labels[6][151] , \labels[6][150] , \labels[6][149] , 
	\labels[6][148] , \labels[6][147] , \labels[6][146] , 
	\labels[6][145] , \labels[6][144] , \labels[6][143] , 
	\labels[6][142] , \labels[6][141] , \labels[6][140] , 
	\labels[6][139] , \labels[6][138] , \labels[6][137] , 
	\labels[6][136] , \labels[6][135] , \labels[6][134] , 
	\labels[6][133] , \labels[6][132] , \labels[6][131] , 
	\labels[6][130] , \labels[6][129] , \labels[6][128] , 
	\labels[6][127] , \labels[6][126] , \labels[6][125] , 
	\labels[6][124] , \labels[6][123] , \labels[6][122] , 
	\labels[6][121] , \labels[6][120] , \labels[6][119] , 
	\labels[6][118] , \labels[6][117] , \labels[6][116] , 
	\labels[6][115] , \labels[6][114] , \labels[6][113] , 
	\labels[6][112] , \labels[6][111] , \labels[6][110] , 
	\labels[6][109] , \labels[6][108] , \labels[6][107] , 
	\labels[6][106] , \labels[6][105] , \labels[6][104] , 
	\labels[6][103] , \labels[6][102] , \labels[6][101] , 
	\labels[6][100] , \labels[6][99] , \labels[6][98] , \labels[6][97] , 
	\labels[6][96] , \labels[6][95] , \labels[6][94] , \labels[6][93] , 
	\labels[6][92] , \labels[6][91] , \labels[6][90] , \labels[6][89] , 
	\labels[6][88] , \labels[6][87] , \labels[6][86] , \labels[6][85] , 
	\labels[6][84] , \labels[6][83] , \labels[6][82] , \labels[6][81] , 
	\labels[6][80] , \labels[6][79] , \labels[6][78] , \labels[6][77] , 
	\labels[6][76] , \labels[6][75] , \labels[6][74] , \labels[6][73] , 
	\labels[6][72] , \labels[6][71] , \labels[6][70] , \labels[6][69] , 
	\labels[6][68] , \labels[6][67] , \labels[6][66] , \labels[6][65] , 
	\labels[6][64] , \labels[6][63] , \labels[6][62] , \labels[6][61] , 
	\labels[6][60] , \labels[6][59] , \labels[6][58] , \labels[6][57] , 
	\labels[6][56] , \labels[6][55] , \labels[6][54] , \labels[6][53] , 
	\labels[6][52] , \labels[6][51] , \labels[6][50] , \labels[6][49] , 
	\labels[6][48] , \labels[6][47] , \labels[6][46] , \labels[6][45] , 
	\labels[6][44] , \labels[6][43] , \labels[6][42] , \labels[6][41] , 
	\labels[6][40] , \labels[6][39] , \labels[6][38] , \labels[6][37] , 
	\labels[6][36] , \labels[6][35] , \labels[6][34] , \labels[6][33] , 
	\labels[6][32] , \labels[6][31] , \labels[6][30] , \labels[6][29] , 
	\labels[6][28] , \labels[6][27] , \labels[6][26] , \labels[6][25] , 
	\labels[6][24] , \labels[6][23] , \labels[6][22] , \labels[6][21] , 
	\labels[6][20] , \labels[6][19] , \labels[6][18] , \labels[6][17] , 
	\labels[6][16] , \labels[6][15] , \labels[6][14] , \labels[6][13] , 
	\labels[6][12] , \labels[6][11] , \labels[6][10] , \labels[6][9] , 
	\labels[6][8] , \labels[6][7] , \labels[6][6] , \labels[6][5] , 
	\labels[6][4] , \labels[6][3] , \labels[6][2] , \labels[6][1] , 
	\labels[6][0] , \labels[5][271] , \labels[5][270] , \labels[5][269] , 
	\labels[5][268] , \labels[5][267] , \labels[5][266] , 
	\labels[5][265] , \labels[5][264] , \labels[5][263] , 
	\labels[5][262] , \labels[5][261] , \labels[5][260] , 
	\labels[5][259] , \labels[5][258] , \labels[5][257] , 
	\labels[5][256] , \labels[5][255] , \labels[5][254] , 
	\labels[5][253] , \labels[5][252] , \labels[5][251] , 
	\labels[5][250] , \labels[5][249] , \labels[5][248] , 
	\labels[5][247] , \labels[5][246] , \labels[5][245] , 
	\labels[5][244] , \labels[5][243] , \labels[5][242] , 
	\labels[5][241] , \labels[5][240] , \labels[5][239] , 
	\labels[5][238] , \labels[5][237] , \labels[5][236] , 
	\labels[5][235] , \labels[5][234] , \labels[5][233] , 
	\labels[5][232] , \labels[5][231] , \labels[5][230] , 
	\labels[5][229] , \labels[5][228] , \labels[5][227] , 
	\labels[5][226] , \labels[5][225] , \labels[5][224] , 
	\labels[5][223] , \labels[5][222] , \labels[5][221] , 
	\labels[5][220] , \labels[5][219] , \labels[5][218] , 
	\labels[5][217] , \labels[5][216] , \labels[5][215] , 
	\labels[5][214] , \labels[5][213] , \labels[5][212] , 
	\labels[5][211] , \labels[5][210] , \labels[5][209] , 
	\labels[5][208] , \labels[5][207] , \labels[5][206] , 
	\labels[5][205] , \labels[5][204] , \labels[5][203] , 
	\labels[5][202] , \labels[5][201] , \labels[5][200] , 
	\labels[5][199] , \labels[5][198] , \labels[5][197] , 
	\labels[5][196] , \labels[5][195] , \labels[5][194] , 
	\labels[5][193] , \labels[5][192] , \labels[5][191] , 
	\labels[5][190] , \labels[5][189] , \labels[5][188] , 
	\labels[5][187] , \labels[5][186] , \labels[5][185] , 
	\labels[5][184] , \labels[5][183] , \labels[5][182] , 
	\labels[5][181] , \labels[5][180] , \labels[5][179] , 
	\labels[5][178] , \labels[5][177] , \labels[5][176] , 
	\labels[5][175] , \labels[5][174] , \labels[5][173] , 
	\labels[5][172] , \labels[5][171] , \labels[5][170] , 
	\labels[5][169] , \labels[5][168] , \labels[5][167] , 
	\labels[5][166] , \labels[5][165] , \labels[5][164] , 
	\labels[5][163] , \labels[5][162] , \labels[5][161] , 
	\labels[5][160] , \labels[5][159] , \labels[5][158] , 
	\labels[5][157] , \labels[5][156] , \labels[5][155] , 
	\labels[5][154] , \labels[5][153] , \labels[5][152] , 
	\labels[5][151] , \labels[5][150] , \labels[5][149] , 
	\labels[5][148] , \labels[5][147] , \labels[5][146] , 
	\labels[5][145] , \labels[5][144] , \labels[5][143] , 
	\labels[5][142] , \labels[5][141] , \labels[5][140] , 
	\labels[5][139] , \labels[5][138] , \labels[5][137] , 
	\labels[5][136] , \labels[5][135] , \labels[5][134] , 
	\labels[5][133] , \labels[5][132] , \labels[5][131] , 
	\labels[5][130] , \labels[5][129] , \labels[5][128] , 
	\labels[5][127] , \labels[5][126] , \labels[5][125] , 
	\labels[5][124] , \labels[5][123] , \labels[5][122] , 
	\labels[5][121] , \labels[5][120] , \labels[5][119] , 
	\labels[5][118] , \labels[5][117] , \labels[5][116] , 
	\labels[5][115] , \labels[5][114] , \labels[5][113] , 
	\labels[5][112] , \labels[5][111] , \labels[5][110] , 
	\labels[5][109] , \labels[5][108] , \labels[5][107] , 
	\labels[5][106] , \labels[5][105] , \labels[5][104] , 
	\labels[5][103] , \labels[5][102] , \labels[5][101] , 
	\labels[5][100] , \labels[5][99] , \labels[5][98] , \labels[5][97] , 
	\labels[5][96] , \labels[5][95] , \labels[5][94] , \labels[5][93] , 
	\labels[5][92] , \labels[5][91] , \labels[5][90] , \labels[5][89] , 
	\labels[5][88] , \labels[5][87] , \labels[5][86] , \labels[5][85] , 
	\labels[5][84] , \labels[5][83] , \labels[5][82] , \labels[5][81] , 
	\labels[5][80] , \labels[5][79] , \labels[5][78] , \labels[5][77] , 
	\labels[5][76] , \labels[5][75] , \labels[5][74] , \labels[5][73] , 
	\labels[5][72] , \labels[5][71] , \labels[5][70] , \labels[5][69] , 
	\labels[5][68] , \labels[5][67] , \labels[5][66] , \labels[5][65] , 
	\labels[5][64] , \labels[5][63] , \labels[5][62] , \labels[5][61] , 
	\labels[5][60] , \labels[5][59] , \labels[5][58] , \labels[5][57] , 
	\labels[5][56] , \labels[5][55] , \labels[5][54] , \labels[5][53] , 
	\labels[5][52] , \labels[5][51] , \labels[5][50] , \labels[5][49] , 
	\labels[5][48] , \labels[5][47] , \labels[5][46] , \labels[5][45] , 
	\labels[5][44] , \labels[5][43] , \labels[5][42] , \labels[5][41] , 
	\labels[5][40] , \labels[5][39] , \labels[5][38] , \labels[5][37] , 
	\labels[5][36] , \labels[5][35] , \labels[5][34] , \labels[5][33] , 
	\labels[5][32] , \labels[5][31] , \labels[5][30] , \labels[5][29] , 
	\labels[5][28] , \labels[5][27] , \labels[5][26] , \labels[5][25] , 
	\labels[5][24] , \labels[5][23] , \labels[5][22] , \labels[5][21] , 
	\labels[5][20] , \labels[5][19] , \labels[5][18] , \labels[5][17] , 
	\labels[5][16] , \labels[5][15] , \labels[5][14] , \labels[5][13] , 
	\labels[5][12] , \labels[5][11] , \labels[5][10] , \labels[5][9] , 
	\labels[5][8] , \labels[5][7] , \labels[5][6] , \labels[5][5] , 
	\labels[5][4] , \labels[5][3] , \labels[5][2] , \labels[5][1] , 
	\labels[5][0] , \labels[4][271] , \labels[4][270] , \labels[4][269] , 
	\labels[4][268] , \labels[4][267] , \labels[4][266] , 
	\labels[4][265] , \labels[4][264] , \labels[4][263] , 
	\labels[4][262] , \labels[4][261] , \labels[4][260] , 
	\labels[4][259] , \labels[4][258] , \labels[4][257] , 
	\labels[4][256] , \labels[4][255] , \labels[4][254] , 
	\labels[4][253] , \labels[4][252] , \labels[4][251] , 
	\labels[4][250] , \labels[4][249] , \labels[4][248] , 
	\labels[4][247] , \labels[4][246] , \labels[4][245] , 
	\labels[4][244] , \labels[4][243] , \labels[4][242] , 
	\labels[4][241] , \labels[4][240] , \labels[4][239] , 
	\labels[4][238] , \labels[4][237] , \labels[4][236] , 
	\labels[4][235] , \labels[4][234] , \labels[4][233] , 
	\labels[4][232] , \labels[4][231] , \labels[4][230] , 
	\labels[4][229] , \labels[4][228] , \labels[4][227] , 
	\labels[4][226] , \labels[4][225] , \labels[4][224] , 
	\labels[4][223] , \labels[4][222] , \labels[4][221] , 
	\labels[4][220] , \labels[4][219] , \labels[4][218] , 
	\labels[4][217] , \labels[4][216] , \labels[4][215] , 
	\labels[4][214] , \labels[4][213] , \labels[4][212] , 
	\labels[4][211] , \labels[4][210] , \labels[4][209] , 
	\labels[4][208] , \labels[4][207] , \labels[4][206] , 
	\labels[4][205] , \labels[4][204] , \labels[4][203] , 
	\labels[4][202] , \labels[4][201] , \labels[4][200] , 
	\labels[4][199] , \labels[4][198] , \labels[4][197] , 
	\labels[4][196] , \labels[4][195] , \labels[4][194] , 
	\labels[4][193] , \labels[4][192] , \labels[4][191] , 
	\labels[4][190] , \labels[4][189] , \labels[4][188] , 
	\labels[4][187] , \labels[4][186] , \labels[4][185] , 
	\labels[4][184] , \labels[4][183] , \labels[4][182] , 
	\labels[4][181] , \labels[4][180] , \labels[4][179] , 
	\labels[4][178] , \labels[4][177] , \labels[4][176] , 
	\labels[4][175] , \labels[4][174] , \labels[4][173] , 
	\labels[4][172] , \labels[4][171] , \labels[4][170] , 
	\labels[4][169] , \labels[4][168] , \labels[4][167] , 
	\labels[4][166] , \labels[4][165] , \labels[4][164] , 
	\labels[4][163] , \labels[4][162] , \labels[4][161] , 
	\labels[4][160] , \labels[4][159] , \labels[4][158] , 
	\labels[4][157] , \labels[4][156] , \labels[4][155] , 
	\labels[4][154] , \labels[4][153] , \labels[4][152] , 
	\labels[4][151] , \labels[4][150] , \labels[4][149] , 
	\labels[4][148] , \labels[4][147] , \labels[4][146] , 
	\labels[4][145] , \labels[4][144] , \labels[4][143] , 
	\labels[4][142] , \labels[4][141] , \labels[4][140] , 
	\labels[4][139] , \labels[4][138] , \labels[4][137] , 
	\labels[4][136] , \labels[4][135] , \labels[4][134] , 
	\labels[4][133] , \labels[4][132] , \labels[4][131] , 
	\labels[4][130] , \labels[4][129] , \labels[4][128] , 
	\labels[4][127] , \labels[4][126] , \labels[4][125] , 
	\labels[4][124] , \labels[4][123] , \labels[4][122] , 
	\labels[4][121] , \labels[4][120] , \labels[4][119] , 
	\labels[4][118] , \labels[4][117] , \labels[4][116] , 
	\labels[4][115] , \labels[4][114] , \labels[4][113] , 
	\labels[4][112] , \labels[4][111] , \labels[4][110] , 
	\labels[4][109] , \labels[4][108] , \labels[4][107] , 
	\labels[4][106] , \labels[4][105] , \labels[4][104] , 
	\labels[4][103] , \labels[4][102] , \labels[4][101] , 
	\labels[4][100] , \labels[4][99] , \labels[4][98] , \labels[4][97] , 
	\labels[4][96] , \labels[4][95] , \labels[4][94] , \labels[4][93] , 
	\labels[4][92] , \labels[4][91] , \labels[4][90] , \labels[4][89] , 
	\labels[4][88] , \labels[4][87] , \labels[4][86] , \labels[4][85] , 
	\labels[4][84] , \labels[4][83] , \labels[4][82] , \labels[4][81] , 
	\labels[4][80] , \labels[4][79] , \labels[4][78] , \labels[4][77] , 
	\labels[4][76] , \labels[4][75] , \labels[4][74] , \labels[4][73] , 
	\labels[4][72] , \labels[4][71] , \labels[4][70] , \labels[4][69] , 
	\labels[4][68] , \labels[4][67] , \labels[4][66] , \labels[4][65] , 
	\labels[4][64] , \labels[4][63] , \labels[4][62] , \labels[4][61] , 
	\labels[4][60] , \labels[4][59] , \labels[4][58] , \labels[4][57] , 
	\labels[4][56] , \labels[4][55] , \labels[4][54] , \labels[4][53] , 
	\labels[4][52] , \labels[4][51] , \labels[4][50] , \labels[4][49] , 
	\labels[4][48] , \labels[4][47] , \labels[4][46] , \labels[4][45] , 
	\labels[4][44] , \labels[4][43] , \labels[4][42] , \labels[4][41] , 
	\labels[4][40] , \labels[4][39] , \labels[4][38] , \labels[4][37] , 
	\labels[4][36] , \labels[4][35] , \labels[4][34] , \labels[4][33] , 
	\labels[4][32] , \labels[4][31] , \labels[4][30] , \labels[4][29] , 
	\labels[4][28] , \labels[4][27] , \labels[4][26] , \labels[4][25] , 
	\labels[4][24] , \labels[4][23] , \labels[4][22] , \labels[4][21] , 
	\labels[4][20] , \labels[4][19] , \labels[4][18] , \labels[4][17] , 
	\labels[4][16] , \labels[4][15] , \labels[4][14] , \labels[4][13] , 
	\labels[4][12] , \labels[4][11] , \labels[4][10] , \labels[4][9] , 
	\labels[4][8] , \labels[4][7] , \labels[4][6] , \labels[4][5] , 
	\labels[4][4] , \labels[4][3] , \labels[4][2] , \labels[4][1] , 
	\labels[4][0] , \labels[3][271] , \labels[3][270] , \labels[3][269] , 
	\labels[3][268] , \labels[3][267] , \labels[3][266] , 
	\labels[3][265] , \labels[3][264] , \labels[3][263] , 
	\labels[3][262] , \labels[3][261] , \labels[3][260] , 
	\labels[3][259] , \labels[3][258] , \labels[3][257] , 
	\labels[3][256] , \labels[3][255] , \labels[3][254] , 
	\labels[3][253] , \labels[3][252] , \labels[3][251] , 
	\labels[3][250] , \labels[3][249] , \labels[3][248] , 
	\labels[3][247] , \labels[3][246] , \labels[3][245] , 
	\labels[3][244] , \labels[3][243] , \labels[3][242] , 
	\labels[3][241] , \labels[3][240] , \labels[3][239] , 
	\labels[3][238] , \labels[3][237] , \labels[3][236] , 
	\labels[3][235] , \labels[3][234] , \labels[3][233] , 
	\labels[3][232] , \labels[3][231] , \labels[3][230] , 
	\labels[3][229] , \labels[3][228] , \labels[3][227] , 
	\labels[3][226] , \labels[3][225] , \labels[3][224] , 
	\labels[3][223] , \labels[3][222] , \labels[3][221] , 
	\labels[3][220] , \labels[3][219] , \labels[3][218] , 
	\labels[3][217] , \labels[3][216] , \labels[3][215] , 
	\labels[3][214] , \labels[3][213] , \labels[3][212] , 
	\labels[3][211] , \labels[3][210] , \labels[3][209] , 
	\labels[3][208] , \labels[3][207] , \labels[3][206] , 
	\labels[3][205] , \labels[3][204] , \labels[3][203] , 
	\labels[3][202] , \labels[3][201] , \labels[3][200] , 
	\labels[3][199] , \labels[3][198] , \labels[3][197] , 
	\labels[3][196] , \labels[3][195] , \labels[3][194] , 
	\labels[3][193] , \labels[3][192] , \labels[3][191] , 
	\labels[3][190] , \labels[3][189] , \labels[3][188] , 
	\labels[3][187] , \labels[3][186] , \labels[3][185] , 
	\labels[3][184] , \labels[3][183] , \labels[3][182] , 
	\labels[3][181] , \labels[3][180] , \labels[3][179] , 
	\labels[3][178] , \labels[3][177] , \labels[3][176] , 
	\labels[3][175] , \labels[3][174] , \labels[3][173] , 
	\labels[3][172] , \labels[3][171] , \labels[3][170] , 
	\labels[3][169] , \labels[3][168] , \labels[3][167] , 
	\labels[3][166] , \labels[3][165] , \labels[3][164] , 
	\labels[3][163] , \labels[3][162] , \labels[3][161] , 
	\labels[3][160] , \labels[3][159] , \labels[3][158] , 
	\labels[3][157] , \labels[3][156] , \labels[3][155] , 
	\labels[3][154] , \labels[3][153] , \labels[3][152] , 
	\labels[3][151] , \labels[3][150] , \labels[3][149] , 
	\labels[3][148] , \labels[3][147] , \labels[3][146] , 
	\labels[3][145] , \labels[3][144] , \labels[3][143] , 
	\labels[3][142] , \labels[3][141] , \labels[3][140] , 
	\labels[3][139] , \labels[3][138] , \labels[3][137] , 
	\labels[3][136] , \labels[3][135] , \labels[3][134] , 
	\labels[3][133] , \labels[3][132] , \labels[3][131] , 
	\labels[3][130] , \labels[3][129] , \labels[3][128] , 
	\labels[3][127] , \labels[3][126] , \labels[3][125] , 
	\labels[3][124] , \labels[3][123] , \labels[3][122] , 
	\labels[3][121] , \labels[3][120] , \labels[3][119] , 
	\labels[3][118] , \labels[3][117] , \labels[3][116] , 
	\labels[3][115] , \labels[3][114] , \labels[3][113] , 
	\labels[3][112] , \labels[3][111] , \labels[3][110] , 
	\labels[3][109] , \labels[3][108] , \labels[3][107] , 
	\labels[3][106] , \labels[3][105] , \labels[3][104] , 
	\labels[3][103] , \labels[3][102] , \labels[3][101] , 
	\labels[3][100] , \labels[3][99] , \labels[3][98] , \labels[3][97] , 
	\labels[3][96] , \labels[3][95] , \labels[3][94] , \labels[3][93] , 
	\labels[3][92] , \labels[3][91] , \labels[3][90] , \labels[3][89] , 
	\labels[3][88] , \labels[3][87] , \labels[3][86] , \labels[3][85] , 
	\labels[3][84] , \labels[3][83] , \labels[3][82] , \labels[3][81] , 
	\labels[3][80] , \labels[3][79] , \labels[3][78] , \labels[3][77] , 
	\labels[3][76] , \labels[3][75] , \labels[3][74] , \labels[3][73] , 
	\labels[3][72] , \labels[3][71] , \labels[3][70] , \labels[3][69] , 
	\labels[3][68] , \labels[3][67] , \labels[3][66] , \labels[3][65] , 
	\labels[3][64] , \labels[3][63] , \labels[3][62] , \labels[3][61] , 
	\labels[3][60] , \labels[3][59] , \labels[3][58] , \labels[3][57] , 
	\labels[3][56] , \labels[3][55] , \labels[3][54] , \labels[3][53] , 
	\labels[3][52] , \labels[3][51] , \labels[3][50] , \labels[3][49] , 
	\labels[3][48] , \labels[3][47] , \labels[3][46] , \labels[3][45] , 
	\labels[3][44] , \labels[3][43] , \labels[3][42] , \labels[3][41] , 
	\labels[3][40] , \labels[3][39] , \labels[3][38] , \labels[3][37] , 
	\labels[3][36] , \labels[3][35] , \labels[3][34] , \labels[3][33] , 
	\labels[3][32] , \labels[3][31] , \labels[3][30] , \labels[3][29] , 
	\labels[3][28] , \labels[3][27] , \labels[3][26] , \labels[3][25] , 
	\labels[3][24] , \labels[3][23] , \labels[3][22] , \labels[3][21] , 
	\labels[3][20] , \labels[3][19] , \labels[3][18] , \labels[3][17] , 
	\labels[3][16] , \labels[3][15] , \labels[3][14] , \labels[3][13] , 
	\labels[3][12] , \labels[3][11] , \labels[3][10] , \labels[3][9] , 
	\labels[3][8] , \labels[3][7] , \labels[3][6] , \labels[3][5] , 
	\labels[3][4] , \labels[3][3] , \labels[3][2] , \labels[3][1] , 
	\labels[3][0] , \labels[2][271] , \labels[2][270] , \labels[2][269] , 
	\labels[2][268] , \labels[2][267] , \labels[2][266] , 
	\labels[2][265] , \labels[2][264] , \labels[2][263] , 
	\labels[2][262] , \labels[2][261] , \labels[2][260] , 
	\labels[2][259] , \labels[2][258] , \labels[2][257] , 
	\labels[2][256] , \labels[2][255] , \labels[2][254] , 
	\labels[2][253] , \labels[2][252] , \labels[2][251] , 
	\labels[2][250] , \labels[2][249] , \labels[2][248] , 
	\labels[2][247] , \labels[2][246] , \labels[2][245] , 
	\labels[2][244] , \labels[2][243] , \labels[2][242] , 
	\labels[2][241] , \labels[2][240] , \labels[2][239] , 
	\labels[2][238] , \labels[2][237] , \labels[2][236] , 
	\labels[2][235] , \labels[2][234] , \labels[2][233] , 
	\labels[2][232] , \labels[2][231] , \labels[2][230] , 
	\labels[2][229] , \labels[2][228] , \labels[2][227] , 
	\labels[2][226] , \labels[2][225] , \labels[2][224] , 
	\labels[2][223] , \labels[2][222] , \labels[2][221] , 
	\labels[2][220] , \labels[2][219] , \labels[2][218] , 
	\labels[2][217] , \labels[2][216] , \labels[2][215] , 
	\labels[2][214] , \labels[2][213] , \labels[2][212] , 
	\labels[2][211] , \labels[2][210] , \labels[2][209] , 
	\labels[2][208] , \labels[2][207] , \labels[2][206] , 
	\labels[2][205] , \labels[2][204] , \labels[2][203] , 
	\labels[2][202] , \labels[2][201] , \labels[2][200] , 
	\labels[2][199] , \labels[2][198] , \labels[2][197] , 
	\labels[2][196] , \labels[2][195] , \labels[2][194] , 
	\labels[2][193] , \labels[2][192] , \labels[2][191] , 
	\labels[2][190] , \labels[2][189] , \labels[2][188] , 
	\labels[2][187] , \labels[2][186] , \labels[2][185] , 
	\labels[2][184] , \labels[2][183] , \labels[2][182] , 
	\labels[2][181] , \labels[2][180] , \labels[2][179] , 
	\labels[2][178] , \labels[2][177] , \labels[2][176] , 
	\labels[2][175] , \labels[2][174] , \labels[2][173] , 
	\labels[2][172] , \labels[2][171] , \labels[2][170] , 
	\labels[2][169] , \labels[2][168] , \labels[2][167] , 
	\labels[2][166] , \labels[2][165] , \labels[2][164] , 
	\labels[2][163] , \labels[2][162] , \labels[2][161] , 
	\labels[2][160] , \labels[2][159] , \labels[2][158] , 
	\labels[2][157] , \labels[2][156] , \labels[2][155] , 
	\labels[2][154] , \labels[2][153] , \labels[2][152] , 
	\labels[2][151] , \labels[2][150] , \labels[2][149] , 
	\labels[2][148] , \labels[2][147] , \labels[2][146] , 
	\labels[2][145] , \labels[2][144] , \labels[2][143] , 
	\labels[2][142] , \labels[2][141] , \labels[2][140] , 
	\labels[2][139] , \labels[2][138] , \labels[2][137] , 
	\labels[2][136] , \labels[2][135] , \labels[2][134] , 
	\labels[2][133] , \labels[2][132] , \labels[2][131] , 
	\labels[2][130] , \labels[2][129] , \labels[2][128] , 
	\labels[2][127] , \labels[2][126] , \labels[2][125] , 
	\labels[2][124] , \labels[2][123] , \labels[2][122] , 
	\labels[2][121] , \labels[2][120] , \labels[2][119] , 
	\labels[2][118] , \labels[2][117] , \labels[2][116] , 
	\labels[2][115] , \labels[2][114] , \labels[2][113] , 
	\labels[2][112] , \labels[2][111] , \labels[2][110] , 
	\labels[2][109] , \labels[2][108] , \labels[2][107] , 
	\labels[2][106] , \labels[2][105] , \labels[2][104] , 
	\labels[2][103] , \labels[2][102] , \labels[2][101] , 
	\labels[2][100] , \labels[2][99] , \labels[2][98] , \labels[2][97] , 
	\labels[2][96] , \labels[2][95] , \labels[2][94] , \labels[2][93] , 
	\labels[2][92] , \labels[2][91] , \labels[2][90] , \labels[2][89] , 
	\labels[2][88] , \labels[2][87] , \labels[2][86] , \labels[2][85] , 
	\labels[2][84] , \labels[2][83] , \labels[2][82] , \labels[2][81] , 
	\labels[2][80] , \labels[2][79] , \labels[2][78] , \labels[2][77] , 
	\labels[2][76] , \labels[2][75] , \labels[2][74] , \labels[2][73] , 
	\labels[2][72] , \labels[2][71] , \labels[2][70] , \labels[2][69] , 
	\labels[2][68] , \labels[2][67] , \labels[2][66] , \labels[2][65] , 
	\labels[2][64] , \labels[2][63] , \labels[2][62] , \labels[2][61] , 
	\labels[2][60] , \labels[2][59] , \labels[2][58] , \labels[2][57] , 
	\labels[2][56] , \labels[2][55] , \labels[2][54] , \labels[2][53] , 
	\labels[2][52] , \labels[2][51] , \labels[2][50] , \labels[2][49] , 
	\labels[2][48] , \labels[2][47] , \labels[2][46] , \labels[2][45] , 
	\labels[2][44] , \labels[2][43] , \labels[2][42] , \labels[2][41] , 
	\labels[2][40] , \labels[2][39] , \labels[2][38] , \labels[2][37] , 
	\labels[2][36] , \labels[2][35] , \labels[2][34] , \labels[2][33] , 
	\labels[2][32] , \labels[2][31] , \labels[2][30] , \labels[2][29] , 
	\labels[2][28] , \labels[2][27] , \labels[2][26] , \labels[2][25] , 
	\labels[2][24] , \labels[2][23] , \labels[2][22] , \labels[2][21] , 
	\labels[2][20] , \labels[2][19] , \labels[2][18] , \labels[2][17] , 
	\labels[2][16] , \labels[2][15] , \labels[2][14] , \labels[2][13] , 
	\labels[2][12] , \labels[2][11] , \labels[2][10] , \labels[2][9] , 
	\labels[2][8] , \labels[2][7] , \labels[2][6] , \labels[2][5] , 
	\labels[2][4] , \labels[2][3] , \labels[2][2] , \labels[2][1] , 
	\labels[2][0] , \labels[1][271] , \labels[1][270] , \labels[1][269] , 
	\labels[1][268] , \labels[1][267] , \labels[1][266] , 
	\labels[1][265] , \labels[1][264] , \labels[1][263] , 
	\labels[1][262] , \labels[1][261] , \labels[1][260] , 
	\labels[1][259] , \labels[1][258] , \labels[1][257] , 
	\labels[1][256] , \labels[1][255] , \labels[1][254] , 
	\labels[1][253] , \labels[1][252] , \labels[1][251] , 
	\labels[1][250] , \labels[1][249] , \labels[1][248] , 
	\labels[1][247] , \labels[1][246] , \labels[1][245] , 
	\labels[1][244] , \labels[1][243] , \labels[1][242] , 
	\labels[1][241] , \labels[1][240] , \labels[1][239] , 
	\labels[1][238] , \labels[1][237] , \labels[1][236] , 
	\labels[1][235] , \labels[1][234] , \labels[1][233] , 
	\labels[1][232] , \labels[1][231] , \labels[1][230] , 
	\labels[1][229] , \labels[1][228] , \labels[1][227] , 
	\labels[1][226] , \labels[1][225] , \labels[1][224] , 
	\labels[1][223] , \labels[1][222] , \labels[1][221] , 
	\labels[1][220] , \labels[1][219] , \labels[1][218] , 
	\labels[1][217] , \labels[1][216] , \labels[1][215] , 
	\labels[1][214] , \labels[1][213] , \labels[1][212] , 
	\labels[1][211] , \labels[1][210] , \labels[1][209] , 
	\labels[1][208] , \labels[1][207] , \labels[1][206] , 
	\labels[1][205] , \labels[1][204] , \labels[1][203] , 
	\labels[1][202] , \labels[1][201] , \labels[1][200] , 
	\labels[1][199] , \labels[1][198] , \labels[1][197] , 
	\labels[1][196] , \labels[1][195] , \labels[1][194] , 
	\labels[1][193] , \labels[1][192] , \labels[1][191] , 
	\labels[1][190] , \labels[1][189] , \labels[1][188] , 
	\labels[1][187] , \labels[1][186] , \labels[1][185] , 
	\labels[1][184] , \labels[1][183] , \labels[1][182] , 
	\labels[1][181] , \labels[1][180] , \labels[1][179] , 
	\labels[1][178] , \labels[1][177] , \labels[1][176] , 
	\labels[1][175] , \labels[1][174] , \labels[1][173] , 
	\labels[1][172] , \labels[1][171] , \labels[1][170] , 
	\labels[1][169] , \labels[1][168] , \labels[1][167] , 
	\labels[1][166] , \labels[1][165] , \labels[1][164] , 
	\labels[1][163] , \labels[1][162] , \labels[1][161] , 
	\labels[1][160] , \labels[1][159] , \labels[1][158] , 
	\labels[1][157] , \labels[1][156] , \labels[1][155] , 
	\labels[1][154] , \labels[1][153] , \labels[1][152] , 
	\labels[1][151] , \labels[1][150] , \labels[1][149] , 
	\labels[1][148] , \labels[1][147] , \labels[1][146] , 
	\labels[1][145] , \labels[1][144] , \labels[1][143] , 
	\labels[1][142] , \labels[1][141] , \labels[1][140] , 
	\labels[1][139] , \labels[1][138] , \labels[1][137] , 
	\labels[1][136] , \labels[1][135] , \labels[1][134] , 
	\labels[1][133] , \labels[1][132] , \labels[1][131] , 
	\labels[1][130] , \labels[1][129] , \labels[1][128] , 
	\labels[1][127] , \labels[1][126] , \labels[1][125] , 
	\labels[1][124] , \labels[1][123] , \labels[1][122] , 
	\labels[1][121] , \labels[1][120] , \labels[1][119] , 
	\labels[1][118] , \labels[1][117] , \labels[1][116] , 
	\labels[1][115] , \labels[1][114] , \labels[1][113] , 
	\labels[1][112] , \labels[1][111] , \labels[1][110] , 
	\labels[1][109] , \labels[1][108] , \labels[1][107] , 
	\labels[1][106] , \labels[1][105] , \labels[1][104] , 
	\labels[1][103] , \labels[1][102] , \labels[1][101] , 
	\labels[1][100] , \labels[1][99] , \labels[1][98] , \labels[1][97] , 
	\labels[1][96] , \labels[1][95] , \labels[1][94] , \labels[1][93] , 
	\labels[1][92] , \labels[1][91] , \labels[1][90] , \labels[1][89] , 
	\labels[1][88] , \labels[1][87] , \labels[1][86] , \labels[1][85] , 
	\labels[1][84] , \labels[1][83] , \labels[1][82] , \labels[1][81] , 
	\labels[1][80] , \labels[1][79] , \labels[1][78] , \labels[1][77] , 
	\labels[1][76] , \labels[1][75] , \labels[1][74] , \labels[1][73] , 
	\labels[1][72] , \labels[1][71] , \labels[1][70] , \labels[1][69] , 
	\labels[1][68] , \labels[1][67] , \labels[1][66] , \labels[1][65] , 
	\labels[1][64] , \labels[1][63] , \labels[1][62] , \labels[1][61] , 
	\labels[1][60] , \labels[1][59] , \labels[1][58] , \labels[1][57] , 
	\labels[1][56] , \labels[1][55] , \labels[1][54] , \labels[1][53] , 
	\labels[1][52] , \labels[1][51] , \labels[1][50] , \labels[1][49] , 
	\labels[1][48] , \labels[1][47] , \labels[1][46] , \labels[1][45] , 
	\labels[1][44] , \labels[1][43] , \labels[1][42] , \labels[1][41] , 
	\labels[1][40] , \labels[1][39] , \labels[1][38] , \labels[1][37] , 
	\labels[1][36] , \labels[1][35] , \labels[1][34] , \labels[1][33] , 
	\labels[1][32] , \labels[1][31] , \labels[1][30] , \labels[1][29] , 
	\labels[1][28] , \labels[1][27] , \labels[1][26] , \labels[1][25] , 
	\labels[1][24] , \labels[1][23] , \labels[1][22] , \labels[1][21] , 
	\labels[1][20] , \labels[1][19] , \labels[1][18] , \labels[1][17] , 
	\labels[1][16] , \labels[1][15] , \labels[1][14] , \labels[1][13] , 
	\labels[1][12] , \labels[1][11] , \labels[1][10] , \labels[1][9] , 
	\labels[1][8] , \labels[1][7] , \labels[1][6] , \labels[1][5] , 
	\labels[1][4] , \labels[1][3] , \labels[1][2] , \labels[1][1] , 
	\labels[1][0] , \labels[0][271] , \labels[0][270] , \labels[0][269] , 
	\labels[0][268] , \labels[0][267] , \labels[0][266] , 
	\labels[0][265] , \labels[0][264] , \labels[0][263] , 
	\labels[0][262] , \labels[0][261] , \labels[0][260] , 
	\labels[0][259] , \labels[0][258] , \labels[0][257] , 
	\labels[0][256] , \labels[0][255] , \labels[0][254] , 
	\labels[0][253] , \labels[0][252] , \labels[0][251] , 
	\labels[0][250] , \labels[0][249] , \labels[0][248] , 
	\labels[0][247] , \labels[0][246] , \labels[0][245] , 
	\labels[0][244] , \labels[0][243] , \labels[0][242] , 
	\labels[0][241] , \labels[0][240] , \labels[0][239] , 
	\labels[0][238] , \labels[0][237] , \labels[0][236] , 
	\labels[0][235] , \labels[0][234] , \labels[0][233] , 
	\labels[0][232] , \labels[0][231] , \labels[0][230] , 
	\labels[0][229] , \labels[0][228] , \labels[0][227] , 
	\labels[0][226] , \labels[0][225] , \labels[0][224] , 
	\labels[0][223] , \labels[0][222] , \labels[0][221] , 
	\labels[0][220] , \labels[0][219] , \labels[0][218] , 
	\labels[0][217] , \labels[0][216] , \labels[0][215] , 
	\labels[0][214] , \labels[0][213] , \labels[0][212] , 
	\labels[0][211] , \labels[0][210] , \labels[0][209] , 
	\labels[0][208] , \labels[0][207] , \labels[0][206] , 
	\labels[0][205] , \labels[0][204] , \labels[0][203] , 
	\labels[0][202] , \labels[0][201] , \labels[0][200] , 
	\labels[0][199] , \labels[0][198] , \labels[0][197] , 
	\labels[0][196] , \labels[0][195] , \labels[0][194] , 
	\labels[0][193] , \labels[0][192] , \labels[0][191] , 
	\labels[0][190] , \labels[0][189] , \labels[0][188] , 
	\labels[0][187] , \labels[0][186] , \labels[0][185] , 
	\labels[0][184] , \labels[0][183] , \labels[0][182] , 
	\labels[0][181] , \labels[0][180] , \labels[0][179] , 
	\labels[0][178] , \labels[0][177] , \labels[0][176] , 
	\labels[0][175] , \labels[0][174] , \labels[0][173] , 
	\labels[0][172] , \labels[0][171] , \labels[0][170] , 
	\labels[0][169] , \labels[0][168] , \labels[0][167] , 
	\labels[0][166] , \labels[0][165] , \labels[0][164] , 
	\labels[0][163] , \labels[0][162] , \labels[0][161] , 
	\labels[0][160] , \labels[0][159] , \labels[0][158] , 
	\labels[0][157] , \labels[0][156] , \labels[0][155] , 
	\labels[0][154] , \labels[0][153] , \labels[0][152] , 
	\labels[0][151] , \labels[0][150] , \labels[0][149] , 
	\labels[0][148] , \labels[0][147] , \labels[0][146] , 
	\labels[0][145] , \labels[0][144] , \labels[0][143] , 
	\labels[0][142] , \labels[0][141] , \labels[0][140] , 
	\labels[0][139] , \labels[0][138] , \labels[0][137] , 
	\labels[0][136] , \labels[0][135] , \labels[0][134] , 
	\labels[0][133] , \labels[0][132] , \labels[0][131] , 
	\labels[0][130] , \labels[0][129] , \labels[0][128] , 
	\labels[0][127] , \labels[0][126] , \labels[0][125] , 
	\labels[0][124] , \labels[0][123] , \labels[0][122] , 
	\labels[0][121] , \labels[0][120] , \labels[0][119] , 
	\labels[0][118] , \labels[0][117] , \labels[0][116] , 
	\labels[0][115] , \labels[0][114] , \labels[0][113] , 
	\labels[0][112] , \labels[0][111] , \labels[0][110] , 
	\labels[0][109] , \labels[0][108] , \labels[0][107] , 
	\labels[0][106] , \labels[0][105] , \labels[0][104] , 
	\labels[0][103] , \labels[0][102] , \labels[0][101] , 
	\labels[0][100] , \labels[0][99] , \labels[0][98] , \labels[0][97] , 
	\labels[0][96] , \labels[0][95] , \labels[0][94] , \labels[0][93] , 
	\labels[0][92] , \labels[0][91] , \labels[0][90] , \labels[0][89] , 
	\labels[0][88] , \labels[0][87] , \labels[0][86] , \labels[0][85] , 
	\labels[0][84] , \labels[0][83] , \labels[0][82] , \labels[0][81] , 
	\labels[0][80] , \labels[0][79] , \labels[0][78] , \labels[0][77] , 
	\labels[0][76] , \labels[0][75] , \labels[0][74] , \labels[0][73] , 
	\labels[0][72] , \labels[0][71] , \labels[0][70] , \labels[0][69] , 
	\labels[0][68] , \labels[0][67] , \labels[0][66] , \labels[0][65] , 
	\labels[0][64] , \labels[0][63] , \labels[0][62] , \labels[0][61] , 
	\labels[0][60] , \labels[0][59] , \labels[0][58] , \labels[0][57] , 
	\labels[0][56] , \labels[0][55] , \labels[0][54] , \labels[0][53] , 
	\labels[0][52] , \labels[0][51] , \labels[0][50] , \labels[0][49] , 
	\labels[0][48] , \labels[0][47] , \labels[0][46] , \labels[0][45] , 
	\labels[0][44] , \labels[0][43] , \labels[0][42] , \labels[0][41] , 
	\labels[0][40] , \labels[0][39] , \labels[0][38] , \labels[0][37] , 
	\labels[0][36] , \labels[0][35] , \labels[0][34] , \labels[0][33] , 
	\labels[0][32] , \labels[0][31] , \labels[0][30] , \labels[0][29] , 
	\labels[0][28] , \labels[0][27] , \labels[0][26] , \labels[0][25] , 
	\labels[0][24] , \labels[0][23] , \labels[0][22] , \labels[0][21] , 
	\labels[0][20] , \labels[0][19] , \labels[0][18] , \labels[0][17] , 
	\labels[0][16] , \labels[0][15] , \labels[0][14] , \labels[0][13] , 
	\labels[0][12] , \labels[0][11] , \labels[0][10] , \labels[0][9] , 
	\labels[0][8] , \labels[0][7] , \labels[0][6] , \labels[0][5] , 
	\labels[0][4] , \labels[0][3] , \labels[0][2] , \labels[0][1] , 
	\labels[0][0] });
ixc_assign_38 _zz_strnp_17 ( _zy_simnet_kim_dout_17_w$[0:37], kim_dout[37:0]);
ixc_assign _zz_strnp_16 ( _zy_simnet_kme_cddip3_ob_in_mod_16_w$, 
	kme_cddip3_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_15 ( _zy_simnet_kme_cddip3_ob_out_15_w$[0:82], 
	kme_cddip3_ob_out[82:0]);
ixc_assign _zz_strnp_14 ( _zy_simnet_kme_cddip2_ob_in_mod_14_w$, 
	kme_cddip2_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_13 ( _zy_simnet_kme_cddip2_ob_out_13_w$[0:82], 
	kme_cddip2_ob_out[82:0]);
ixc_assign _zz_strnp_12 ( _zy_simnet_kme_cddip1_ob_in_mod_12_w$, 
	kme_cddip1_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_11 ( _zy_simnet_kme_cddip1_ob_out_11_w$[0:82], 
	kme_cddip1_ob_out[82:0]);
ixc_assign _zz_strnp_10 ( _zy_simnet_kme_cddip0_ob_in_mod_10_w$, 
	kme_cddip0_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_9 ( _zy_simnet_kme_cddip0_ob_out_9_w$[0:82], 
	kme_cddip0_ob_out[82:0]);
ixc_assign _zz_strnp_8 ( _zy_simnet_kme_cceip3_ob_in_mod_8_w$, 
	kme_cceip3_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_7 ( _zy_simnet_kme_cceip3_ob_out_7_w$[0:82], 
	kme_cceip3_ob_out[82:0]);
ixc_assign _zz_strnp_6 ( _zy_simnet_kme_cceip2_ob_in_mod_6_w$, 
	kme_cceip2_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_5 ( _zy_simnet_kme_cceip2_ob_out_5_w$[0:82], 
	kme_cceip2_ob_out[82:0]);
ixc_assign _zz_strnp_4 ( _zy_simnet_kme_cceip1_ob_in_mod_4_w$, 
	kme_cceip1_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_3 ( _zy_simnet_kme_cceip1_ob_out_3_w$[0:82], 
	kme_cceip1_ob_out[82:0]);
ixc_assign _zz_strnp_2 ( _zy_simnet_kme_cceip0_ob_in_mod_2_w$, 
	kme_cceip0_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_1 ( _zy_simnet_kme_cceip0_ob_out_1_w$[0:82], 
	kme_cceip0_ob_out[82:0]);
Q_AN02 U2849 ( .A0(n3), .A1(cceip0_out_ia_rdata[0]), .Z(_zy_simnet_tvar_229[31]));
Q_AN02 U2850 ( .A0(n3), .A1(cceip0_out_ia_rdata[1]), .Z(_zy_simnet_tvar_229[30]));
Q_AN02 U2851 ( .A0(n3), .A1(cceip0_out_ia_rdata[2]), .Z(_zy_simnet_tvar_229[29]));
Q_AN02 U2852 ( .A0(n3), .A1(cceip0_out_ia_rdata[3]), .Z(_zy_simnet_tvar_229[28]));
Q_AN02 U2853 ( .A0(n3), .A1(cceip0_out_ia_rdata[4]), .Z(_zy_simnet_tvar_229[27]));
Q_AN02 U2854 ( .A0(n3), .A1(cceip0_out_ia_rdata[5]), .Z(_zy_simnet_tvar_229[26]));
Q_AN02 U2855 ( .A0(n3), .A1(cceip0_out_ia_rdata[6]), .Z(_zy_simnet_tvar_229[25]));
Q_AN02 U2856 ( .A0(n3), .A1(cceip0_out_ia_rdata[7]), .Z(_zy_simnet_tvar_229[24]));
Q_AN02 U2857 ( .A0(n3), .A1(cceip0_out_ia_rdata[8]), .Z(_zy_simnet_tvar_229[23]));
Q_AN02 U2858 ( .A0(n3), .A1(cceip0_out_ia_rdata[9]), .Z(_zy_simnet_tvar_229[22]));
Q_AN02 U2859 ( .A0(n3), .A1(cceip0_out_ia_rdata[10]), .Z(_zy_simnet_tvar_229[21]));
Q_AN02 U2860 ( .A0(n3), .A1(cceip0_out_ia_rdata[11]), .Z(_zy_simnet_tvar_229[20]));
Q_AN02 U2861 ( .A0(n3), .A1(cceip0_out_ia_rdata[12]), .Z(_zy_simnet_tvar_229[19]));
Q_AN02 U2862 ( .A0(n3), .A1(cceip0_out_ia_rdata[13]), .Z(_zy_simnet_tvar_229[18]));
Q_AN02 U2863 ( .A0(n3), .A1(cceip0_out_ia_rdata[14]), .Z(_zy_simnet_tvar_229[17]));
Q_AN02 U2864 ( .A0(n3), .A1(cceip0_out_ia_rdata[15]), .Z(_zy_simnet_tvar_229[16]));
Q_AN02 U2865 ( .A0(n3), .A1(cceip0_out_ia_rdata[16]), .Z(_zy_simnet_tvar_229[15]));
Q_AN02 U2866 ( .A0(n3), .A1(cceip0_out_ia_rdata[17]), .Z(_zy_simnet_tvar_229[14]));
Q_AN02 U2867 ( .A0(n3), .A1(cceip0_out_ia_rdata[18]), .Z(_zy_simnet_tvar_229[13]));
Q_AN02 U2868 ( .A0(n3), .A1(cceip0_out_ia_rdata[19]), .Z(_zy_simnet_tvar_229[12]));
Q_AN02 U2869 ( .A0(n3), .A1(cceip0_out_ia_rdata[20]), .Z(_zy_simnet_tvar_229[11]));
Q_AN02 U2870 ( .A0(n3), .A1(cceip0_out_ia_rdata[21]), .Z(_zy_simnet_tvar_229[10]));
Q_AN02 U2871 ( .A0(n3), .A1(cceip0_out_ia_rdata[22]), .Z(_zy_simnet_tvar_229[9]));
Q_AN02 U2872 ( .A0(n3), .A1(cceip0_out_ia_rdata[23]), .Z(_zy_simnet_tvar_229[8]));
Q_AN02 U2873 ( .A0(n3), .A1(cceip0_out_ia_rdata[24]), .Z(_zy_simnet_tvar_229[7]));
Q_AN02 U2874 ( .A0(n3), .A1(cceip0_out_ia_rdata[25]), .Z(_zy_simnet_tvar_229[6]));
Q_AN02 U2875 ( .A0(n3), .A1(cceip0_out_ia_rdata[26]), .Z(_zy_simnet_tvar_229[5]));
Q_AN02 U2876 ( .A0(n3), .A1(cceip0_out_ia_rdata[27]), .Z(_zy_simnet_tvar_229[4]));
Q_AN02 U2877 ( .A0(n3), .A1(cceip0_out_ia_rdata[28]), .Z(_zy_simnet_tvar_229[3]));
Q_AN02 U2878 ( .A0(n3), .A1(cceip0_out_ia_rdata[29]), .Z(_zy_simnet_tvar_229[2]));
Q_AN02 U2879 ( .A0(n3), .A1(cceip0_out_ia_rdata[30]), .Z(_zy_simnet_tvar_229[1]));
Q_AN02 U2880 ( .A0(n3), .A1(cceip0_out_ia_rdata[31]), .Z(_zy_simnet_tvar_229[0]));
Q_INV U2881 ( .A(disable_ckv_kim_ism_reads), .Z(n3));
Q_AN02 U2882 ( .A0(n3), .A1(cceip0_out_ia_rdata[32]), .Z(_zy_simnet_tvar_230[31]));
Q_AN02 U2883 ( .A0(n3), .A1(cceip0_out_ia_rdata[33]), .Z(_zy_simnet_tvar_230[30]));
Q_AN02 U2884 ( .A0(n3), .A1(cceip0_out_ia_rdata[34]), .Z(_zy_simnet_tvar_230[29]));
Q_AN02 U2885 ( .A0(n3), .A1(cceip0_out_ia_rdata[35]), .Z(_zy_simnet_tvar_230[28]));
Q_AN02 U2886 ( .A0(n3), .A1(cceip0_out_ia_rdata[36]), .Z(_zy_simnet_tvar_230[27]));
Q_AN02 U2887 ( .A0(n3), .A1(cceip0_out_ia_rdata[37]), .Z(_zy_simnet_tvar_230[26]));
Q_AN02 U2888 ( .A0(n3), .A1(cceip0_out_ia_rdata[38]), .Z(_zy_simnet_tvar_230[25]));
Q_AN02 U2889 ( .A0(n3), .A1(cceip0_out_ia_rdata[39]), .Z(_zy_simnet_tvar_230[24]));
Q_AN02 U2890 ( .A0(n3), .A1(cceip0_out_ia_rdata[40]), .Z(_zy_simnet_tvar_230[23]));
Q_AN02 U2891 ( .A0(n3), .A1(cceip0_out_ia_rdata[41]), .Z(_zy_simnet_tvar_230[22]));
Q_AN02 U2892 ( .A0(n3), .A1(cceip0_out_ia_rdata[42]), .Z(_zy_simnet_tvar_230[21]));
Q_AN02 U2893 ( .A0(n3), .A1(cceip0_out_ia_rdata[43]), .Z(_zy_simnet_tvar_230[20]));
Q_AN02 U2894 ( .A0(n3), .A1(cceip0_out_ia_rdata[44]), .Z(_zy_simnet_tvar_230[19]));
Q_AN02 U2895 ( .A0(n3), .A1(cceip0_out_ia_rdata[45]), .Z(_zy_simnet_tvar_230[18]));
Q_AN02 U2896 ( .A0(n3), .A1(cceip0_out_ia_rdata[46]), .Z(_zy_simnet_tvar_230[17]));
Q_AN02 U2897 ( .A0(n3), .A1(cceip0_out_ia_rdata[47]), .Z(_zy_simnet_tvar_230[16]));
Q_AN02 U2898 ( .A0(n3), .A1(cceip0_out_ia_rdata[48]), .Z(_zy_simnet_tvar_230[15]));
Q_AN02 U2899 ( .A0(n3), .A1(cceip0_out_ia_rdata[49]), .Z(_zy_simnet_tvar_230[14]));
Q_AN02 U2900 ( .A0(n3), .A1(cceip0_out_ia_rdata[50]), .Z(_zy_simnet_tvar_230[13]));
Q_AN02 U2901 ( .A0(n3), .A1(cceip0_out_ia_rdata[51]), .Z(_zy_simnet_tvar_230[12]));
Q_AN02 U2902 ( .A0(n3), .A1(cceip0_out_ia_rdata[52]), .Z(_zy_simnet_tvar_230[11]));
Q_AN02 U2903 ( .A0(n3), .A1(cceip0_out_ia_rdata[53]), .Z(_zy_simnet_tvar_230[10]));
Q_AN02 U2904 ( .A0(n3), .A1(cceip0_out_ia_rdata[54]), .Z(_zy_simnet_tvar_230[9]));
Q_AN02 U2905 ( .A0(n3), .A1(cceip0_out_ia_rdata[55]), .Z(_zy_simnet_tvar_230[8]));
Q_AN02 U2906 ( .A0(n3), .A1(cceip0_out_ia_rdata[56]), .Z(_zy_simnet_tvar_230[7]));
Q_AN02 U2907 ( .A0(n3), .A1(cceip0_out_ia_rdata[57]), .Z(_zy_simnet_tvar_230[6]));
Q_AN02 U2908 ( .A0(n3), .A1(cceip0_out_ia_rdata[58]), .Z(_zy_simnet_tvar_230[5]));
Q_AN02 U2909 ( .A0(n3), .A1(cceip0_out_ia_rdata[59]), .Z(_zy_simnet_tvar_230[4]));
Q_AN02 U2910 ( .A0(n3), .A1(cceip0_out_ia_rdata[60]), .Z(_zy_simnet_tvar_230[3]));
Q_AN02 U2911 ( .A0(n3), .A1(cceip0_out_ia_rdata[61]), .Z(_zy_simnet_tvar_230[2]));
Q_AN02 U2912 ( .A0(n3), .A1(cceip0_out_ia_rdata[62]), .Z(_zy_simnet_tvar_230[1]));
Q_AN02 U2913 ( .A0(n3), .A1(cceip0_out_ia_rdata[63]), .Z(_zy_simnet_tvar_230[0]));
Q_AN02 U2914 ( .A0(n3), .A1(cceip0_out_ia_rdata[64]), .Z(_zy_simnet_tvar_231[31]));
Q_AN02 U2915 ( .A0(n3), .A1(cceip0_out_ia_rdata[65]), .Z(_zy_simnet_tvar_231[30]));
Q_AN02 U2916 ( .A0(n3), .A1(cceip0_out_ia_rdata[66]), .Z(_zy_simnet_tvar_231[29]));
Q_AN02 U2917 ( .A0(n3), .A1(cceip0_out_ia_rdata[67]), .Z(_zy_simnet_tvar_231[28]));
Q_AN02 U2918 ( .A0(n3), .A1(cceip0_out_ia_rdata[68]), .Z(_zy_simnet_tvar_231[27]));
Q_AN02 U2919 ( .A0(n3), .A1(cceip0_out_ia_rdata[69]), .Z(_zy_simnet_tvar_231[26]));
Q_AN02 U2920 ( .A0(n3), .A1(cceip0_out_ia_rdata[70]), .Z(_zy_simnet_tvar_231[25]));
Q_AN02 U2921 ( .A0(n3), .A1(cceip0_out_ia_rdata[71]), .Z(_zy_simnet_tvar_231[24]));
Q_AN02 U2922 ( .A0(n3), .A1(cceip0_out_ia_rdata[72]), .Z(_zy_simnet_tvar_231[23]));
Q_AN02 U2923 ( .A0(n3), .A1(cceip0_out_ia_rdata[73]), .Z(_zy_simnet_tvar_231[22]));
Q_AN02 U2924 ( .A0(n3), .A1(cceip0_out_ia_rdata[74]), .Z(_zy_simnet_tvar_231[21]));
Q_AN02 U2925 ( .A0(n3), .A1(cceip0_out_ia_rdata[75]), .Z(_zy_simnet_tvar_231[20]));
Q_AN02 U2926 ( .A0(n3), .A1(cceip0_out_ia_rdata[76]), .Z(_zy_simnet_tvar_231[19]));
Q_AN02 U2927 ( .A0(n3), .A1(cceip0_out_ia_rdata[77]), .Z(_zy_simnet_tvar_231[18]));
Q_AN02 U2928 ( .A0(n3), .A1(cceip0_out_ia_rdata[78]), .Z(_zy_simnet_tvar_231[17]));
Q_AN02 U2929 ( .A0(n3), .A1(cceip0_out_ia_rdata[79]), .Z(_zy_simnet_tvar_231[16]));
Q_AN02 U2930 ( .A0(n3), .A1(cceip0_out_ia_rdata[80]), .Z(_zy_simnet_tvar_231[15]));
Q_AN02 U2931 ( .A0(n3), .A1(cceip0_out_ia_rdata[81]), .Z(_zy_simnet_tvar_231[14]));
Q_AN02 U2932 ( .A0(n3), .A1(cceip0_out_ia_rdata[82]), .Z(_zy_simnet_tvar_231[13]));
Q_AN02 U2933 ( .A0(n3), .A1(cceip0_out_ia_rdata[83]), .Z(_zy_simnet_tvar_231[12]));
Q_AN02 U2934 ( .A0(n3), .A1(cceip0_out_ia_rdata[84]), .Z(_zy_simnet_tvar_231[11]));
Q_AN02 U2935 ( .A0(n3), .A1(cceip0_out_ia_rdata[85]), .Z(_zy_simnet_tvar_231[10]));
Q_AN02 U2936 ( .A0(n3), .A1(cceip0_out_ia_rdata[86]), .Z(_zy_simnet_tvar_231[9]));
Q_AN02 U2937 ( .A0(n3), .A1(cceip0_out_ia_rdata[87]), .Z(_zy_simnet_tvar_231[8]));
Q_AN02 U2938 ( .A0(n3), .A1(cceip0_out_ia_rdata[88]), .Z(_zy_simnet_tvar_231[7]));
Q_AN02 U2939 ( .A0(n3), .A1(cceip0_out_ia_rdata[89]), .Z(_zy_simnet_tvar_231[6]));
Q_AN02 U2940 ( .A0(n3), .A1(cceip0_out_ia_rdata[90]), .Z(_zy_simnet_tvar_231[5]));
Q_AN02 U2941 ( .A0(n3), .A1(cceip0_out_ia_rdata[91]), .Z(_zy_simnet_tvar_231[4]));
Q_AN02 U2942 ( .A0(n3), .A1(cceip0_out_ia_rdata[92]), .Z(_zy_simnet_tvar_231[3]));
Q_AN02 U2943 ( .A0(n3), .A1(cceip0_out_ia_rdata[93]), .Z(_zy_simnet_tvar_231[2]));
Q_AN02 U2944 ( .A0(n3), .A1(cceip0_out_ia_rdata[94]), .Z(_zy_simnet_tvar_231[1]));
Q_AN02 U2945 ( .A0(n3), .A1(cceip0_out_ia_rdata[95]), .Z(_zy_simnet_tvar_231[0]));
Q_AN02 U2946 ( .A0(n3), .A1(cceip1_out_ia_rdata[0]), .Z(_zy_simnet_tvar_236[31]));
Q_AN02 U2947 ( .A0(n3), .A1(cceip1_out_ia_rdata[1]), .Z(_zy_simnet_tvar_236[30]));
Q_AN02 U2948 ( .A0(n3), .A1(cceip1_out_ia_rdata[2]), .Z(_zy_simnet_tvar_236[29]));
Q_AN02 U2949 ( .A0(n3), .A1(cceip1_out_ia_rdata[3]), .Z(_zy_simnet_tvar_236[28]));
Q_AN02 U2950 ( .A0(n3), .A1(cceip1_out_ia_rdata[4]), .Z(_zy_simnet_tvar_236[27]));
Q_AN02 U2951 ( .A0(n3), .A1(cceip1_out_ia_rdata[5]), .Z(_zy_simnet_tvar_236[26]));
Q_AN02 U2952 ( .A0(n3), .A1(cceip1_out_ia_rdata[6]), .Z(_zy_simnet_tvar_236[25]));
Q_AN02 U2953 ( .A0(n3), .A1(cceip1_out_ia_rdata[7]), .Z(_zy_simnet_tvar_236[24]));
Q_AN02 U2954 ( .A0(n3), .A1(cceip1_out_ia_rdata[8]), .Z(_zy_simnet_tvar_236[23]));
Q_AN02 U2955 ( .A0(n3), .A1(cceip1_out_ia_rdata[9]), .Z(_zy_simnet_tvar_236[22]));
Q_AN02 U2956 ( .A0(n3), .A1(cceip1_out_ia_rdata[10]), .Z(_zy_simnet_tvar_236[21]));
Q_AN02 U2957 ( .A0(n3), .A1(cceip1_out_ia_rdata[11]), .Z(_zy_simnet_tvar_236[20]));
Q_AN02 U2958 ( .A0(n3), .A1(cceip1_out_ia_rdata[12]), .Z(_zy_simnet_tvar_236[19]));
Q_AN02 U2959 ( .A0(n3), .A1(cceip1_out_ia_rdata[13]), .Z(_zy_simnet_tvar_236[18]));
Q_AN02 U2960 ( .A0(n3), .A1(cceip1_out_ia_rdata[14]), .Z(_zy_simnet_tvar_236[17]));
Q_AN02 U2961 ( .A0(n3), .A1(cceip1_out_ia_rdata[15]), .Z(_zy_simnet_tvar_236[16]));
Q_AN02 U2962 ( .A0(n3), .A1(cceip1_out_ia_rdata[16]), .Z(_zy_simnet_tvar_236[15]));
Q_AN02 U2963 ( .A0(n3), .A1(cceip1_out_ia_rdata[17]), .Z(_zy_simnet_tvar_236[14]));
Q_AN02 U2964 ( .A0(n3), .A1(cceip1_out_ia_rdata[18]), .Z(_zy_simnet_tvar_236[13]));
Q_AN02 U2965 ( .A0(n3), .A1(cceip1_out_ia_rdata[19]), .Z(_zy_simnet_tvar_236[12]));
Q_AN02 U2966 ( .A0(n3), .A1(cceip1_out_ia_rdata[20]), .Z(_zy_simnet_tvar_236[11]));
Q_AN02 U2967 ( .A0(n3), .A1(cceip1_out_ia_rdata[21]), .Z(_zy_simnet_tvar_236[10]));
Q_AN02 U2968 ( .A0(n3), .A1(cceip1_out_ia_rdata[22]), .Z(_zy_simnet_tvar_236[9]));
Q_AN02 U2969 ( .A0(n3), .A1(cceip1_out_ia_rdata[23]), .Z(_zy_simnet_tvar_236[8]));
Q_AN02 U2970 ( .A0(n3), .A1(cceip1_out_ia_rdata[24]), .Z(_zy_simnet_tvar_236[7]));
Q_AN02 U2971 ( .A0(n3), .A1(cceip1_out_ia_rdata[25]), .Z(_zy_simnet_tvar_236[6]));
Q_AN02 U2972 ( .A0(n3), .A1(cceip1_out_ia_rdata[26]), .Z(_zy_simnet_tvar_236[5]));
Q_AN02 U2973 ( .A0(n3), .A1(cceip1_out_ia_rdata[27]), .Z(_zy_simnet_tvar_236[4]));
Q_AN02 U2974 ( .A0(n3), .A1(cceip1_out_ia_rdata[28]), .Z(_zy_simnet_tvar_236[3]));
Q_AN02 U2975 ( .A0(n3), .A1(cceip1_out_ia_rdata[29]), .Z(_zy_simnet_tvar_236[2]));
Q_AN02 U2976 ( .A0(n3), .A1(cceip1_out_ia_rdata[30]), .Z(_zy_simnet_tvar_236[1]));
Q_AN02 U2977 ( .A0(n3), .A1(cceip1_out_ia_rdata[31]), .Z(_zy_simnet_tvar_236[0]));
Q_AN02 U2978 ( .A0(n3), .A1(cceip1_out_ia_rdata[32]), .Z(_zy_simnet_tvar_237[31]));
Q_AN02 U2979 ( .A0(n3), .A1(cceip1_out_ia_rdata[33]), .Z(_zy_simnet_tvar_237[30]));
Q_AN02 U2980 ( .A0(n3), .A1(cceip1_out_ia_rdata[34]), .Z(_zy_simnet_tvar_237[29]));
Q_AN02 U2981 ( .A0(n3), .A1(cceip1_out_ia_rdata[35]), .Z(_zy_simnet_tvar_237[28]));
Q_AN02 U2982 ( .A0(n3), .A1(cceip1_out_ia_rdata[36]), .Z(_zy_simnet_tvar_237[27]));
Q_AN02 U2983 ( .A0(n3), .A1(cceip1_out_ia_rdata[37]), .Z(_zy_simnet_tvar_237[26]));
Q_AN02 U2984 ( .A0(n3), .A1(cceip1_out_ia_rdata[38]), .Z(_zy_simnet_tvar_237[25]));
Q_AN02 U2985 ( .A0(n3), .A1(cceip1_out_ia_rdata[39]), .Z(_zy_simnet_tvar_237[24]));
Q_AN02 U2986 ( .A0(n3), .A1(cceip1_out_ia_rdata[40]), .Z(_zy_simnet_tvar_237[23]));
Q_AN02 U2987 ( .A0(n3), .A1(cceip1_out_ia_rdata[41]), .Z(_zy_simnet_tvar_237[22]));
Q_AN02 U2988 ( .A0(n3), .A1(cceip1_out_ia_rdata[42]), .Z(_zy_simnet_tvar_237[21]));
Q_AN02 U2989 ( .A0(n3), .A1(cceip1_out_ia_rdata[43]), .Z(_zy_simnet_tvar_237[20]));
Q_AN02 U2990 ( .A0(n3), .A1(cceip1_out_ia_rdata[44]), .Z(_zy_simnet_tvar_237[19]));
Q_AN02 U2991 ( .A0(n3), .A1(cceip1_out_ia_rdata[45]), .Z(_zy_simnet_tvar_237[18]));
Q_AN02 U2992 ( .A0(n3), .A1(cceip1_out_ia_rdata[46]), .Z(_zy_simnet_tvar_237[17]));
Q_AN02 U2993 ( .A0(n3), .A1(cceip1_out_ia_rdata[47]), .Z(_zy_simnet_tvar_237[16]));
Q_AN02 U2994 ( .A0(n3), .A1(cceip1_out_ia_rdata[48]), .Z(_zy_simnet_tvar_237[15]));
Q_AN02 U2995 ( .A0(n3), .A1(cceip1_out_ia_rdata[49]), .Z(_zy_simnet_tvar_237[14]));
Q_AN02 U2996 ( .A0(n3), .A1(cceip1_out_ia_rdata[50]), .Z(_zy_simnet_tvar_237[13]));
Q_AN02 U2997 ( .A0(n3), .A1(cceip1_out_ia_rdata[51]), .Z(_zy_simnet_tvar_237[12]));
Q_AN02 U2998 ( .A0(n3), .A1(cceip1_out_ia_rdata[52]), .Z(_zy_simnet_tvar_237[11]));
Q_AN02 U2999 ( .A0(n3), .A1(cceip1_out_ia_rdata[53]), .Z(_zy_simnet_tvar_237[10]));
Q_AN02 U3000 ( .A0(n3), .A1(cceip1_out_ia_rdata[54]), .Z(_zy_simnet_tvar_237[9]));
Q_AN02 U3001 ( .A0(n3), .A1(cceip1_out_ia_rdata[55]), .Z(_zy_simnet_tvar_237[8]));
Q_AN02 U3002 ( .A0(n3), .A1(cceip1_out_ia_rdata[56]), .Z(_zy_simnet_tvar_237[7]));
Q_AN02 U3003 ( .A0(n3), .A1(cceip1_out_ia_rdata[57]), .Z(_zy_simnet_tvar_237[6]));
Q_AN02 U3004 ( .A0(n3), .A1(cceip1_out_ia_rdata[58]), .Z(_zy_simnet_tvar_237[5]));
Q_AN02 U3005 ( .A0(n3), .A1(cceip1_out_ia_rdata[59]), .Z(_zy_simnet_tvar_237[4]));
Q_AN02 U3006 ( .A0(n3), .A1(cceip1_out_ia_rdata[60]), .Z(_zy_simnet_tvar_237[3]));
Q_AN02 U3007 ( .A0(n3), .A1(cceip1_out_ia_rdata[61]), .Z(_zy_simnet_tvar_237[2]));
Q_AN02 U3008 ( .A0(n3), .A1(cceip1_out_ia_rdata[62]), .Z(_zy_simnet_tvar_237[1]));
Q_AN02 U3009 ( .A0(n3), .A1(cceip1_out_ia_rdata[63]), .Z(_zy_simnet_tvar_237[0]));
Q_AN02 U3010 ( .A0(n3), .A1(cceip1_out_ia_rdata[64]), .Z(_zy_simnet_tvar_238[31]));
Q_AN02 U3011 ( .A0(n3), .A1(cceip1_out_ia_rdata[65]), .Z(_zy_simnet_tvar_238[30]));
Q_AN02 U3012 ( .A0(n3), .A1(cceip1_out_ia_rdata[66]), .Z(_zy_simnet_tvar_238[29]));
Q_AN02 U3013 ( .A0(n3), .A1(cceip1_out_ia_rdata[67]), .Z(_zy_simnet_tvar_238[28]));
Q_AN02 U3014 ( .A0(n3), .A1(cceip1_out_ia_rdata[68]), .Z(_zy_simnet_tvar_238[27]));
Q_AN02 U3015 ( .A0(n3), .A1(cceip1_out_ia_rdata[69]), .Z(_zy_simnet_tvar_238[26]));
Q_AN02 U3016 ( .A0(n3), .A1(cceip1_out_ia_rdata[70]), .Z(_zy_simnet_tvar_238[25]));
Q_AN02 U3017 ( .A0(n3), .A1(cceip1_out_ia_rdata[71]), .Z(_zy_simnet_tvar_238[24]));
Q_AN02 U3018 ( .A0(n3), .A1(cceip1_out_ia_rdata[72]), .Z(_zy_simnet_tvar_238[23]));
Q_AN02 U3019 ( .A0(n3), .A1(cceip1_out_ia_rdata[73]), .Z(_zy_simnet_tvar_238[22]));
Q_AN02 U3020 ( .A0(n3), .A1(cceip1_out_ia_rdata[74]), .Z(_zy_simnet_tvar_238[21]));
Q_AN02 U3021 ( .A0(n3), .A1(cceip1_out_ia_rdata[75]), .Z(_zy_simnet_tvar_238[20]));
Q_AN02 U3022 ( .A0(n3), .A1(cceip1_out_ia_rdata[76]), .Z(_zy_simnet_tvar_238[19]));
Q_AN02 U3023 ( .A0(n3), .A1(cceip1_out_ia_rdata[77]), .Z(_zy_simnet_tvar_238[18]));
Q_AN02 U3024 ( .A0(n3), .A1(cceip1_out_ia_rdata[78]), .Z(_zy_simnet_tvar_238[17]));
Q_AN02 U3025 ( .A0(n3), .A1(cceip1_out_ia_rdata[79]), .Z(_zy_simnet_tvar_238[16]));
Q_AN02 U3026 ( .A0(n3), .A1(cceip1_out_ia_rdata[80]), .Z(_zy_simnet_tvar_238[15]));
Q_AN02 U3027 ( .A0(n3), .A1(cceip1_out_ia_rdata[81]), .Z(_zy_simnet_tvar_238[14]));
Q_AN02 U3028 ( .A0(n3), .A1(cceip1_out_ia_rdata[82]), .Z(_zy_simnet_tvar_238[13]));
Q_AN02 U3029 ( .A0(n3), .A1(cceip1_out_ia_rdata[83]), .Z(_zy_simnet_tvar_238[12]));
Q_AN02 U3030 ( .A0(n3), .A1(cceip1_out_ia_rdata[84]), .Z(_zy_simnet_tvar_238[11]));
Q_AN02 U3031 ( .A0(n3), .A1(cceip1_out_ia_rdata[85]), .Z(_zy_simnet_tvar_238[10]));
Q_AN02 U3032 ( .A0(n3), .A1(cceip1_out_ia_rdata[86]), .Z(_zy_simnet_tvar_238[9]));
Q_AN02 U3033 ( .A0(n3), .A1(cceip1_out_ia_rdata[87]), .Z(_zy_simnet_tvar_238[8]));
Q_AN02 U3034 ( .A0(n3), .A1(cceip1_out_ia_rdata[88]), .Z(_zy_simnet_tvar_238[7]));
Q_AN02 U3035 ( .A0(n3), .A1(cceip1_out_ia_rdata[89]), .Z(_zy_simnet_tvar_238[6]));
Q_AN02 U3036 ( .A0(n3), .A1(cceip1_out_ia_rdata[90]), .Z(_zy_simnet_tvar_238[5]));
Q_AN02 U3037 ( .A0(n3), .A1(cceip1_out_ia_rdata[91]), .Z(_zy_simnet_tvar_238[4]));
Q_AN02 U3038 ( .A0(n3), .A1(cceip1_out_ia_rdata[92]), .Z(_zy_simnet_tvar_238[3]));
Q_AN02 U3039 ( .A0(n3), .A1(cceip1_out_ia_rdata[93]), .Z(_zy_simnet_tvar_238[2]));
Q_AN02 U3040 ( .A0(n3), .A1(cceip1_out_ia_rdata[94]), .Z(_zy_simnet_tvar_238[1]));
Q_AN02 U3041 ( .A0(n3), .A1(cceip1_out_ia_rdata[95]), .Z(_zy_simnet_tvar_238[0]));
Q_AN02 U3042 ( .A0(n3), .A1(cceip2_out_ia_rdata[0]), .Z(_zy_simnet_tvar_243[31]));
Q_AN02 U3043 ( .A0(n3), .A1(cceip2_out_ia_rdata[1]), .Z(_zy_simnet_tvar_243[30]));
Q_AN02 U3044 ( .A0(n3), .A1(cceip2_out_ia_rdata[2]), .Z(_zy_simnet_tvar_243[29]));
Q_AN02 U3045 ( .A0(n3), .A1(cceip2_out_ia_rdata[3]), .Z(_zy_simnet_tvar_243[28]));
Q_AN02 U3046 ( .A0(n3), .A1(cceip2_out_ia_rdata[4]), .Z(_zy_simnet_tvar_243[27]));
Q_AN02 U3047 ( .A0(n3), .A1(cceip2_out_ia_rdata[5]), .Z(_zy_simnet_tvar_243[26]));
Q_AN02 U3048 ( .A0(n3), .A1(cceip2_out_ia_rdata[6]), .Z(_zy_simnet_tvar_243[25]));
Q_AN02 U3049 ( .A0(n3), .A1(cceip2_out_ia_rdata[7]), .Z(_zy_simnet_tvar_243[24]));
Q_AN02 U3050 ( .A0(n3), .A1(cceip2_out_ia_rdata[8]), .Z(_zy_simnet_tvar_243[23]));
Q_AN02 U3051 ( .A0(n3), .A1(cceip2_out_ia_rdata[9]), .Z(_zy_simnet_tvar_243[22]));
Q_AN02 U3052 ( .A0(n3), .A1(cceip2_out_ia_rdata[10]), .Z(_zy_simnet_tvar_243[21]));
Q_AN02 U3053 ( .A0(n3), .A1(cceip2_out_ia_rdata[11]), .Z(_zy_simnet_tvar_243[20]));
Q_AN02 U3054 ( .A0(n3), .A1(cceip2_out_ia_rdata[12]), .Z(_zy_simnet_tvar_243[19]));
Q_AN02 U3055 ( .A0(n3), .A1(cceip2_out_ia_rdata[13]), .Z(_zy_simnet_tvar_243[18]));
Q_AN02 U3056 ( .A0(n3), .A1(cceip2_out_ia_rdata[14]), .Z(_zy_simnet_tvar_243[17]));
Q_AN02 U3057 ( .A0(n3), .A1(cceip2_out_ia_rdata[15]), .Z(_zy_simnet_tvar_243[16]));
Q_AN02 U3058 ( .A0(n3), .A1(cceip2_out_ia_rdata[16]), .Z(_zy_simnet_tvar_243[15]));
Q_AN02 U3059 ( .A0(n3), .A1(cceip2_out_ia_rdata[17]), .Z(_zy_simnet_tvar_243[14]));
Q_AN02 U3060 ( .A0(n3), .A1(cceip2_out_ia_rdata[18]), .Z(_zy_simnet_tvar_243[13]));
Q_AN02 U3061 ( .A0(n3), .A1(cceip2_out_ia_rdata[19]), .Z(_zy_simnet_tvar_243[12]));
Q_AN02 U3062 ( .A0(n3), .A1(cceip2_out_ia_rdata[20]), .Z(_zy_simnet_tvar_243[11]));
Q_AN02 U3063 ( .A0(n3), .A1(cceip2_out_ia_rdata[21]), .Z(_zy_simnet_tvar_243[10]));
Q_AN02 U3064 ( .A0(n3), .A1(cceip2_out_ia_rdata[22]), .Z(_zy_simnet_tvar_243[9]));
Q_AN02 U3065 ( .A0(n3), .A1(cceip2_out_ia_rdata[23]), .Z(_zy_simnet_tvar_243[8]));
Q_AN02 U3066 ( .A0(n3), .A1(cceip2_out_ia_rdata[24]), .Z(_zy_simnet_tvar_243[7]));
Q_AN02 U3067 ( .A0(n3), .A1(cceip2_out_ia_rdata[25]), .Z(_zy_simnet_tvar_243[6]));
Q_AN02 U3068 ( .A0(n3), .A1(cceip2_out_ia_rdata[26]), .Z(_zy_simnet_tvar_243[5]));
Q_AN02 U3069 ( .A0(n3), .A1(cceip2_out_ia_rdata[27]), .Z(_zy_simnet_tvar_243[4]));
Q_AN02 U3070 ( .A0(n3), .A1(cceip2_out_ia_rdata[28]), .Z(_zy_simnet_tvar_243[3]));
Q_AN02 U3071 ( .A0(n3), .A1(cceip2_out_ia_rdata[29]), .Z(_zy_simnet_tvar_243[2]));
Q_AN02 U3072 ( .A0(n3), .A1(cceip2_out_ia_rdata[30]), .Z(_zy_simnet_tvar_243[1]));
Q_AN02 U3073 ( .A0(n3), .A1(cceip2_out_ia_rdata[31]), .Z(_zy_simnet_tvar_243[0]));
Q_AN02 U3074 ( .A0(n3), .A1(cceip2_out_ia_rdata[32]), .Z(_zy_simnet_tvar_244[31]));
Q_AN02 U3075 ( .A0(n3), .A1(cceip2_out_ia_rdata[33]), .Z(_zy_simnet_tvar_244[30]));
Q_AN02 U3076 ( .A0(n3), .A1(cceip2_out_ia_rdata[34]), .Z(_zy_simnet_tvar_244[29]));
Q_AN02 U3077 ( .A0(n3), .A1(cceip2_out_ia_rdata[35]), .Z(_zy_simnet_tvar_244[28]));
Q_AN02 U3078 ( .A0(n3), .A1(cceip2_out_ia_rdata[36]), .Z(_zy_simnet_tvar_244[27]));
Q_AN02 U3079 ( .A0(n3), .A1(cceip2_out_ia_rdata[37]), .Z(_zy_simnet_tvar_244[26]));
Q_AN02 U3080 ( .A0(n3), .A1(cceip2_out_ia_rdata[38]), .Z(_zy_simnet_tvar_244[25]));
Q_AN02 U3081 ( .A0(n3), .A1(cceip2_out_ia_rdata[39]), .Z(_zy_simnet_tvar_244[24]));
Q_AN02 U3082 ( .A0(n3), .A1(cceip2_out_ia_rdata[40]), .Z(_zy_simnet_tvar_244[23]));
Q_AN02 U3083 ( .A0(n3), .A1(cceip2_out_ia_rdata[41]), .Z(_zy_simnet_tvar_244[22]));
Q_AN02 U3084 ( .A0(n3), .A1(cceip2_out_ia_rdata[42]), .Z(_zy_simnet_tvar_244[21]));
Q_AN02 U3085 ( .A0(n3), .A1(cceip2_out_ia_rdata[43]), .Z(_zy_simnet_tvar_244[20]));
Q_AN02 U3086 ( .A0(n3), .A1(cceip2_out_ia_rdata[44]), .Z(_zy_simnet_tvar_244[19]));
Q_AN02 U3087 ( .A0(n3), .A1(cceip2_out_ia_rdata[45]), .Z(_zy_simnet_tvar_244[18]));
Q_AN02 U3088 ( .A0(n3), .A1(cceip2_out_ia_rdata[46]), .Z(_zy_simnet_tvar_244[17]));
Q_AN02 U3089 ( .A0(n3), .A1(cceip2_out_ia_rdata[47]), .Z(_zy_simnet_tvar_244[16]));
Q_AN02 U3090 ( .A0(n3), .A1(cceip2_out_ia_rdata[48]), .Z(_zy_simnet_tvar_244[15]));
Q_AN02 U3091 ( .A0(n3), .A1(cceip2_out_ia_rdata[49]), .Z(_zy_simnet_tvar_244[14]));
Q_AN02 U3092 ( .A0(n3), .A1(cceip2_out_ia_rdata[50]), .Z(_zy_simnet_tvar_244[13]));
Q_AN02 U3093 ( .A0(n3), .A1(cceip2_out_ia_rdata[51]), .Z(_zy_simnet_tvar_244[12]));
Q_AN02 U3094 ( .A0(n3), .A1(cceip2_out_ia_rdata[52]), .Z(_zy_simnet_tvar_244[11]));
Q_AN02 U3095 ( .A0(n3), .A1(cceip2_out_ia_rdata[53]), .Z(_zy_simnet_tvar_244[10]));
Q_AN02 U3096 ( .A0(n3), .A1(cceip2_out_ia_rdata[54]), .Z(_zy_simnet_tvar_244[9]));
Q_AN02 U3097 ( .A0(n3), .A1(cceip2_out_ia_rdata[55]), .Z(_zy_simnet_tvar_244[8]));
Q_AN02 U3098 ( .A0(n3), .A1(cceip2_out_ia_rdata[56]), .Z(_zy_simnet_tvar_244[7]));
Q_AN02 U3099 ( .A0(n3), .A1(cceip2_out_ia_rdata[57]), .Z(_zy_simnet_tvar_244[6]));
Q_AN02 U3100 ( .A0(n3), .A1(cceip2_out_ia_rdata[58]), .Z(_zy_simnet_tvar_244[5]));
Q_AN02 U3101 ( .A0(n3), .A1(cceip2_out_ia_rdata[59]), .Z(_zy_simnet_tvar_244[4]));
Q_AN02 U3102 ( .A0(n3), .A1(cceip2_out_ia_rdata[60]), .Z(_zy_simnet_tvar_244[3]));
Q_AN02 U3103 ( .A0(n3), .A1(cceip2_out_ia_rdata[61]), .Z(_zy_simnet_tvar_244[2]));
Q_AN02 U3104 ( .A0(n3), .A1(cceip2_out_ia_rdata[62]), .Z(_zy_simnet_tvar_244[1]));
Q_AN02 U3105 ( .A0(n3), .A1(cceip2_out_ia_rdata[63]), .Z(_zy_simnet_tvar_244[0]));
Q_AN02 U3106 ( .A0(n3), .A1(cceip2_out_ia_rdata[64]), .Z(_zy_simnet_tvar_245[31]));
Q_AN02 U3107 ( .A0(n3), .A1(cceip2_out_ia_rdata[65]), .Z(_zy_simnet_tvar_245[30]));
Q_AN02 U3108 ( .A0(n3), .A1(cceip2_out_ia_rdata[66]), .Z(_zy_simnet_tvar_245[29]));
Q_AN02 U3109 ( .A0(n3), .A1(cceip2_out_ia_rdata[67]), .Z(_zy_simnet_tvar_245[28]));
Q_AN02 U3110 ( .A0(n3), .A1(cceip2_out_ia_rdata[68]), .Z(_zy_simnet_tvar_245[27]));
Q_AN02 U3111 ( .A0(n3), .A1(cceip2_out_ia_rdata[69]), .Z(_zy_simnet_tvar_245[26]));
Q_AN02 U3112 ( .A0(n3), .A1(cceip2_out_ia_rdata[70]), .Z(_zy_simnet_tvar_245[25]));
Q_AN02 U3113 ( .A0(n3), .A1(cceip2_out_ia_rdata[71]), .Z(_zy_simnet_tvar_245[24]));
Q_AN02 U3114 ( .A0(n3), .A1(cceip2_out_ia_rdata[72]), .Z(_zy_simnet_tvar_245[23]));
Q_AN02 U3115 ( .A0(n3), .A1(cceip2_out_ia_rdata[73]), .Z(_zy_simnet_tvar_245[22]));
Q_AN02 U3116 ( .A0(n3), .A1(cceip2_out_ia_rdata[74]), .Z(_zy_simnet_tvar_245[21]));
Q_AN02 U3117 ( .A0(n3), .A1(cceip2_out_ia_rdata[75]), .Z(_zy_simnet_tvar_245[20]));
Q_AN02 U3118 ( .A0(n3), .A1(cceip2_out_ia_rdata[76]), .Z(_zy_simnet_tvar_245[19]));
Q_AN02 U3119 ( .A0(n3), .A1(cceip2_out_ia_rdata[77]), .Z(_zy_simnet_tvar_245[18]));
Q_AN02 U3120 ( .A0(n3), .A1(cceip2_out_ia_rdata[78]), .Z(_zy_simnet_tvar_245[17]));
Q_AN02 U3121 ( .A0(n3), .A1(cceip2_out_ia_rdata[79]), .Z(_zy_simnet_tvar_245[16]));
Q_AN02 U3122 ( .A0(n3), .A1(cceip2_out_ia_rdata[80]), .Z(_zy_simnet_tvar_245[15]));
Q_AN02 U3123 ( .A0(n3), .A1(cceip2_out_ia_rdata[81]), .Z(_zy_simnet_tvar_245[14]));
Q_AN02 U3124 ( .A0(n3), .A1(cceip2_out_ia_rdata[82]), .Z(_zy_simnet_tvar_245[13]));
Q_AN02 U3125 ( .A0(n3), .A1(cceip2_out_ia_rdata[83]), .Z(_zy_simnet_tvar_245[12]));
Q_AN02 U3126 ( .A0(n3), .A1(cceip2_out_ia_rdata[84]), .Z(_zy_simnet_tvar_245[11]));
Q_AN02 U3127 ( .A0(n3), .A1(cceip2_out_ia_rdata[85]), .Z(_zy_simnet_tvar_245[10]));
Q_AN02 U3128 ( .A0(n3), .A1(cceip2_out_ia_rdata[86]), .Z(_zy_simnet_tvar_245[9]));
Q_AN02 U3129 ( .A0(n3), .A1(cceip2_out_ia_rdata[87]), .Z(_zy_simnet_tvar_245[8]));
Q_AN02 U3130 ( .A0(n3), .A1(cceip2_out_ia_rdata[88]), .Z(_zy_simnet_tvar_245[7]));
Q_AN02 U3131 ( .A0(n3), .A1(cceip2_out_ia_rdata[89]), .Z(_zy_simnet_tvar_245[6]));
Q_AN02 U3132 ( .A0(n3), .A1(cceip2_out_ia_rdata[90]), .Z(_zy_simnet_tvar_245[5]));
Q_AN02 U3133 ( .A0(n3), .A1(cceip2_out_ia_rdata[91]), .Z(_zy_simnet_tvar_245[4]));
Q_AN02 U3134 ( .A0(n3), .A1(cceip2_out_ia_rdata[92]), .Z(_zy_simnet_tvar_245[3]));
Q_AN02 U3135 ( .A0(n3), .A1(cceip2_out_ia_rdata[93]), .Z(_zy_simnet_tvar_245[2]));
Q_AN02 U3136 ( .A0(n3), .A1(cceip2_out_ia_rdata[94]), .Z(_zy_simnet_tvar_245[1]));
Q_AN02 U3137 ( .A0(n3), .A1(cceip2_out_ia_rdata[95]), .Z(_zy_simnet_tvar_245[0]));
Q_AN02 U3138 ( .A0(n3), .A1(cceip3_out_ia_rdata[0]), .Z(_zy_simnet_tvar_250[31]));
Q_AN02 U3139 ( .A0(n3), .A1(cceip3_out_ia_rdata[1]), .Z(_zy_simnet_tvar_250[30]));
Q_AN02 U3140 ( .A0(n3), .A1(cceip3_out_ia_rdata[2]), .Z(_zy_simnet_tvar_250[29]));
Q_AN02 U3141 ( .A0(n3), .A1(cceip3_out_ia_rdata[3]), .Z(_zy_simnet_tvar_250[28]));
Q_AN02 U3142 ( .A0(n3), .A1(cceip3_out_ia_rdata[4]), .Z(_zy_simnet_tvar_250[27]));
Q_AN02 U3143 ( .A0(n3), .A1(cceip3_out_ia_rdata[5]), .Z(_zy_simnet_tvar_250[26]));
Q_AN02 U3144 ( .A0(n3), .A1(cceip3_out_ia_rdata[6]), .Z(_zy_simnet_tvar_250[25]));
Q_AN02 U3145 ( .A0(n3), .A1(cceip3_out_ia_rdata[7]), .Z(_zy_simnet_tvar_250[24]));
Q_AN02 U3146 ( .A0(n3), .A1(cceip3_out_ia_rdata[8]), .Z(_zy_simnet_tvar_250[23]));
Q_AN02 U3147 ( .A0(n3), .A1(cceip3_out_ia_rdata[9]), .Z(_zy_simnet_tvar_250[22]));
Q_AN02 U3148 ( .A0(n3), .A1(cceip3_out_ia_rdata[10]), .Z(_zy_simnet_tvar_250[21]));
Q_AN02 U3149 ( .A0(n3), .A1(cceip3_out_ia_rdata[11]), .Z(_zy_simnet_tvar_250[20]));
Q_AN02 U3150 ( .A0(n3), .A1(cceip3_out_ia_rdata[12]), .Z(_zy_simnet_tvar_250[19]));
Q_AN02 U3151 ( .A0(n3), .A1(cceip3_out_ia_rdata[13]), .Z(_zy_simnet_tvar_250[18]));
Q_AN02 U3152 ( .A0(n3), .A1(cceip3_out_ia_rdata[14]), .Z(_zy_simnet_tvar_250[17]));
Q_AN02 U3153 ( .A0(n3), .A1(cceip3_out_ia_rdata[15]), .Z(_zy_simnet_tvar_250[16]));
Q_AN02 U3154 ( .A0(n3), .A1(cceip3_out_ia_rdata[16]), .Z(_zy_simnet_tvar_250[15]));
Q_AN02 U3155 ( .A0(n3), .A1(cceip3_out_ia_rdata[17]), .Z(_zy_simnet_tvar_250[14]));
Q_AN02 U3156 ( .A0(n3), .A1(cceip3_out_ia_rdata[18]), .Z(_zy_simnet_tvar_250[13]));
Q_AN02 U3157 ( .A0(n3), .A1(cceip3_out_ia_rdata[19]), .Z(_zy_simnet_tvar_250[12]));
Q_AN02 U3158 ( .A0(n3), .A1(cceip3_out_ia_rdata[20]), .Z(_zy_simnet_tvar_250[11]));
Q_AN02 U3159 ( .A0(n3), .A1(cceip3_out_ia_rdata[21]), .Z(_zy_simnet_tvar_250[10]));
Q_AN02 U3160 ( .A0(n3), .A1(cceip3_out_ia_rdata[22]), .Z(_zy_simnet_tvar_250[9]));
Q_AN02 U3161 ( .A0(n3), .A1(cceip3_out_ia_rdata[23]), .Z(_zy_simnet_tvar_250[8]));
Q_AN02 U3162 ( .A0(n3), .A1(cceip3_out_ia_rdata[24]), .Z(_zy_simnet_tvar_250[7]));
Q_AN02 U3163 ( .A0(n3), .A1(cceip3_out_ia_rdata[25]), .Z(_zy_simnet_tvar_250[6]));
Q_AN02 U3164 ( .A0(n3), .A1(cceip3_out_ia_rdata[26]), .Z(_zy_simnet_tvar_250[5]));
Q_AN02 U3165 ( .A0(n3), .A1(cceip3_out_ia_rdata[27]), .Z(_zy_simnet_tvar_250[4]));
Q_AN02 U3166 ( .A0(n3), .A1(cceip3_out_ia_rdata[28]), .Z(_zy_simnet_tvar_250[3]));
Q_AN02 U3167 ( .A0(n3), .A1(cceip3_out_ia_rdata[29]), .Z(_zy_simnet_tvar_250[2]));
Q_AN02 U3168 ( .A0(n3), .A1(cceip3_out_ia_rdata[30]), .Z(_zy_simnet_tvar_250[1]));
Q_AN02 U3169 ( .A0(n3), .A1(cceip3_out_ia_rdata[31]), .Z(_zy_simnet_tvar_250[0]));
Q_AN02 U3170 ( .A0(n3), .A1(cceip3_out_ia_rdata[32]), .Z(_zy_simnet_tvar_251[31]));
Q_AN02 U3171 ( .A0(n3), .A1(cceip3_out_ia_rdata[33]), .Z(_zy_simnet_tvar_251[30]));
Q_AN02 U3172 ( .A0(n3), .A1(cceip3_out_ia_rdata[34]), .Z(_zy_simnet_tvar_251[29]));
Q_AN02 U3173 ( .A0(n3), .A1(cceip3_out_ia_rdata[35]), .Z(_zy_simnet_tvar_251[28]));
Q_AN02 U3174 ( .A0(n3), .A1(cceip3_out_ia_rdata[36]), .Z(_zy_simnet_tvar_251[27]));
Q_AN02 U3175 ( .A0(n3), .A1(cceip3_out_ia_rdata[37]), .Z(_zy_simnet_tvar_251[26]));
Q_AN02 U3176 ( .A0(n3), .A1(cceip3_out_ia_rdata[38]), .Z(_zy_simnet_tvar_251[25]));
Q_AN02 U3177 ( .A0(n3), .A1(cceip3_out_ia_rdata[39]), .Z(_zy_simnet_tvar_251[24]));
Q_AN02 U3178 ( .A0(n3), .A1(cceip3_out_ia_rdata[40]), .Z(_zy_simnet_tvar_251[23]));
Q_AN02 U3179 ( .A0(n3), .A1(cceip3_out_ia_rdata[41]), .Z(_zy_simnet_tvar_251[22]));
Q_AN02 U3180 ( .A0(n3), .A1(cceip3_out_ia_rdata[42]), .Z(_zy_simnet_tvar_251[21]));
Q_AN02 U3181 ( .A0(n3), .A1(cceip3_out_ia_rdata[43]), .Z(_zy_simnet_tvar_251[20]));
Q_AN02 U3182 ( .A0(n3), .A1(cceip3_out_ia_rdata[44]), .Z(_zy_simnet_tvar_251[19]));
Q_AN02 U3183 ( .A0(n3), .A1(cceip3_out_ia_rdata[45]), .Z(_zy_simnet_tvar_251[18]));
Q_AN02 U3184 ( .A0(n3), .A1(cceip3_out_ia_rdata[46]), .Z(_zy_simnet_tvar_251[17]));
Q_AN02 U3185 ( .A0(n3), .A1(cceip3_out_ia_rdata[47]), .Z(_zy_simnet_tvar_251[16]));
Q_AN02 U3186 ( .A0(n3), .A1(cceip3_out_ia_rdata[48]), .Z(_zy_simnet_tvar_251[15]));
Q_AN02 U3187 ( .A0(n3), .A1(cceip3_out_ia_rdata[49]), .Z(_zy_simnet_tvar_251[14]));
Q_AN02 U3188 ( .A0(n3), .A1(cceip3_out_ia_rdata[50]), .Z(_zy_simnet_tvar_251[13]));
Q_AN02 U3189 ( .A0(n3), .A1(cceip3_out_ia_rdata[51]), .Z(_zy_simnet_tvar_251[12]));
Q_AN02 U3190 ( .A0(n3), .A1(cceip3_out_ia_rdata[52]), .Z(_zy_simnet_tvar_251[11]));
Q_AN02 U3191 ( .A0(n3), .A1(cceip3_out_ia_rdata[53]), .Z(_zy_simnet_tvar_251[10]));
Q_AN02 U3192 ( .A0(n3), .A1(cceip3_out_ia_rdata[54]), .Z(_zy_simnet_tvar_251[9]));
Q_AN02 U3193 ( .A0(n3), .A1(cceip3_out_ia_rdata[55]), .Z(_zy_simnet_tvar_251[8]));
Q_AN02 U3194 ( .A0(n3), .A1(cceip3_out_ia_rdata[56]), .Z(_zy_simnet_tvar_251[7]));
Q_AN02 U3195 ( .A0(n3), .A1(cceip3_out_ia_rdata[57]), .Z(_zy_simnet_tvar_251[6]));
Q_AN02 U3196 ( .A0(n3), .A1(cceip3_out_ia_rdata[58]), .Z(_zy_simnet_tvar_251[5]));
Q_AN02 U3197 ( .A0(n3), .A1(cceip3_out_ia_rdata[59]), .Z(_zy_simnet_tvar_251[4]));
Q_AN02 U3198 ( .A0(n3), .A1(cceip3_out_ia_rdata[60]), .Z(_zy_simnet_tvar_251[3]));
Q_AN02 U3199 ( .A0(n3), .A1(cceip3_out_ia_rdata[61]), .Z(_zy_simnet_tvar_251[2]));
Q_AN02 U3200 ( .A0(n3), .A1(cceip3_out_ia_rdata[62]), .Z(_zy_simnet_tvar_251[1]));
Q_AN02 U3201 ( .A0(n3), .A1(cceip3_out_ia_rdata[63]), .Z(_zy_simnet_tvar_251[0]));
Q_AN02 U3202 ( .A0(n3), .A1(cceip3_out_ia_rdata[64]), .Z(_zy_simnet_tvar_252[31]));
Q_AN02 U3203 ( .A0(n3), .A1(cceip3_out_ia_rdata[65]), .Z(_zy_simnet_tvar_252[30]));
Q_AN02 U3204 ( .A0(n3), .A1(cceip3_out_ia_rdata[66]), .Z(_zy_simnet_tvar_252[29]));
Q_AN02 U3205 ( .A0(n3), .A1(cceip3_out_ia_rdata[67]), .Z(_zy_simnet_tvar_252[28]));
Q_AN02 U3206 ( .A0(n3), .A1(cceip3_out_ia_rdata[68]), .Z(_zy_simnet_tvar_252[27]));
Q_AN02 U3207 ( .A0(n3), .A1(cceip3_out_ia_rdata[69]), .Z(_zy_simnet_tvar_252[26]));
Q_AN02 U3208 ( .A0(n3), .A1(cceip3_out_ia_rdata[70]), .Z(_zy_simnet_tvar_252[25]));
Q_AN02 U3209 ( .A0(n3), .A1(cceip3_out_ia_rdata[71]), .Z(_zy_simnet_tvar_252[24]));
Q_AN02 U3210 ( .A0(n3), .A1(cceip3_out_ia_rdata[72]), .Z(_zy_simnet_tvar_252[23]));
Q_AN02 U3211 ( .A0(n3), .A1(cceip3_out_ia_rdata[73]), .Z(_zy_simnet_tvar_252[22]));
Q_AN02 U3212 ( .A0(n3), .A1(cceip3_out_ia_rdata[74]), .Z(_zy_simnet_tvar_252[21]));
Q_AN02 U3213 ( .A0(n3), .A1(cceip3_out_ia_rdata[75]), .Z(_zy_simnet_tvar_252[20]));
Q_AN02 U3214 ( .A0(n3), .A1(cceip3_out_ia_rdata[76]), .Z(_zy_simnet_tvar_252[19]));
Q_AN02 U3215 ( .A0(n3), .A1(cceip3_out_ia_rdata[77]), .Z(_zy_simnet_tvar_252[18]));
Q_AN02 U3216 ( .A0(n3), .A1(cceip3_out_ia_rdata[78]), .Z(_zy_simnet_tvar_252[17]));
Q_AN02 U3217 ( .A0(n3), .A1(cceip3_out_ia_rdata[79]), .Z(_zy_simnet_tvar_252[16]));
Q_AN02 U3218 ( .A0(n3), .A1(cceip3_out_ia_rdata[80]), .Z(_zy_simnet_tvar_252[15]));
Q_AN02 U3219 ( .A0(n3), .A1(cceip3_out_ia_rdata[81]), .Z(_zy_simnet_tvar_252[14]));
Q_AN02 U3220 ( .A0(n3), .A1(cceip3_out_ia_rdata[82]), .Z(_zy_simnet_tvar_252[13]));
Q_AN02 U3221 ( .A0(n3), .A1(cceip3_out_ia_rdata[83]), .Z(_zy_simnet_tvar_252[12]));
Q_AN02 U3222 ( .A0(n3), .A1(cceip3_out_ia_rdata[84]), .Z(_zy_simnet_tvar_252[11]));
Q_AN02 U3223 ( .A0(n3), .A1(cceip3_out_ia_rdata[85]), .Z(_zy_simnet_tvar_252[10]));
Q_AN02 U3224 ( .A0(n3), .A1(cceip3_out_ia_rdata[86]), .Z(_zy_simnet_tvar_252[9]));
Q_AN02 U3225 ( .A0(n3), .A1(cceip3_out_ia_rdata[87]), .Z(_zy_simnet_tvar_252[8]));
Q_AN02 U3226 ( .A0(n3), .A1(cceip3_out_ia_rdata[88]), .Z(_zy_simnet_tvar_252[7]));
Q_AN02 U3227 ( .A0(n3), .A1(cceip3_out_ia_rdata[89]), .Z(_zy_simnet_tvar_252[6]));
Q_AN02 U3228 ( .A0(n3), .A1(cceip3_out_ia_rdata[90]), .Z(_zy_simnet_tvar_252[5]));
Q_AN02 U3229 ( .A0(n3), .A1(cceip3_out_ia_rdata[91]), .Z(_zy_simnet_tvar_252[4]));
Q_AN02 U3230 ( .A0(n3), .A1(cceip3_out_ia_rdata[92]), .Z(_zy_simnet_tvar_252[3]));
Q_AN02 U3231 ( .A0(n3), .A1(cceip3_out_ia_rdata[93]), .Z(_zy_simnet_tvar_252[2]));
Q_AN02 U3232 ( .A0(n3), .A1(cceip3_out_ia_rdata[94]), .Z(_zy_simnet_tvar_252[1]));
Q_AN02 U3233 ( .A0(n3), .A1(cceip3_out_ia_rdata[95]), .Z(_zy_simnet_tvar_252[0]));
Q_AN02 U3234 ( .A0(n3), .A1(cddip0_out_ia_rdata[0]), .Z(_zy_simnet_tvar_257[31]));
Q_AN02 U3235 ( .A0(n3), .A1(cddip0_out_ia_rdata[1]), .Z(_zy_simnet_tvar_257[30]));
Q_AN02 U3236 ( .A0(n3), .A1(cddip0_out_ia_rdata[2]), .Z(_zy_simnet_tvar_257[29]));
Q_AN02 U3237 ( .A0(n3), .A1(cddip0_out_ia_rdata[3]), .Z(_zy_simnet_tvar_257[28]));
Q_AN02 U3238 ( .A0(n3), .A1(cddip0_out_ia_rdata[4]), .Z(_zy_simnet_tvar_257[27]));
Q_AN02 U3239 ( .A0(n3), .A1(cddip0_out_ia_rdata[5]), .Z(_zy_simnet_tvar_257[26]));
Q_AN02 U3240 ( .A0(n3), .A1(cddip0_out_ia_rdata[6]), .Z(_zy_simnet_tvar_257[25]));
Q_AN02 U3241 ( .A0(n3), .A1(cddip0_out_ia_rdata[7]), .Z(_zy_simnet_tvar_257[24]));
Q_AN02 U3242 ( .A0(n3), .A1(cddip0_out_ia_rdata[8]), .Z(_zy_simnet_tvar_257[23]));
Q_AN02 U3243 ( .A0(n3), .A1(cddip0_out_ia_rdata[9]), .Z(_zy_simnet_tvar_257[22]));
Q_AN02 U3244 ( .A0(n3), .A1(cddip0_out_ia_rdata[10]), .Z(_zy_simnet_tvar_257[21]));
Q_AN02 U3245 ( .A0(n3), .A1(cddip0_out_ia_rdata[11]), .Z(_zy_simnet_tvar_257[20]));
Q_AN02 U3246 ( .A0(n3), .A1(cddip0_out_ia_rdata[12]), .Z(_zy_simnet_tvar_257[19]));
Q_AN02 U3247 ( .A0(n3), .A1(cddip0_out_ia_rdata[13]), .Z(_zy_simnet_tvar_257[18]));
Q_AN02 U3248 ( .A0(n3), .A1(cddip0_out_ia_rdata[14]), .Z(_zy_simnet_tvar_257[17]));
Q_AN02 U3249 ( .A0(n3), .A1(cddip0_out_ia_rdata[15]), .Z(_zy_simnet_tvar_257[16]));
Q_AN02 U3250 ( .A0(n3), .A1(cddip0_out_ia_rdata[16]), .Z(_zy_simnet_tvar_257[15]));
Q_AN02 U3251 ( .A0(n3), .A1(cddip0_out_ia_rdata[17]), .Z(_zy_simnet_tvar_257[14]));
Q_AN02 U3252 ( .A0(n3), .A1(cddip0_out_ia_rdata[18]), .Z(_zy_simnet_tvar_257[13]));
Q_AN02 U3253 ( .A0(n3), .A1(cddip0_out_ia_rdata[19]), .Z(_zy_simnet_tvar_257[12]));
Q_AN02 U3254 ( .A0(n3), .A1(cddip0_out_ia_rdata[20]), .Z(_zy_simnet_tvar_257[11]));
Q_AN02 U3255 ( .A0(n3), .A1(cddip0_out_ia_rdata[21]), .Z(_zy_simnet_tvar_257[10]));
Q_AN02 U3256 ( .A0(n3), .A1(cddip0_out_ia_rdata[22]), .Z(_zy_simnet_tvar_257[9]));
Q_AN02 U3257 ( .A0(n3), .A1(cddip0_out_ia_rdata[23]), .Z(_zy_simnet_tvar_257[8]));
Q_AN02 U3258 ( .A0(n3), .A1(cddip0_out_ia_rdata[24]), .Z(_zy_simnet_tvar_257[7]));
Q_AN02 U3259 ( .A0(n3), .A1(cddip0_out_ia_rdata[25]), .Z(_zy_simnet_tvar_257[6]));
Q_AN02 U3260 ( .A0(n3), .A1(cddip0_out_ia_rdata[26]), .Z(_zy_simnet_tvar_257[5]));
Q_AN02 U3261 ( .A0(n3), .A1(cddip0_out_ia_rdata[27]), .Z(_zy_simnet_tvar_257[4]));
Q_AN02 U3262 ( .A0(n3), .A1(cddip0_out_ia_rdata[28]), .Z(_zy_simnet_tvar_257[3]));
Q_AN02 U3263 ( .A0(n3), .A1(cddip0_out_ia_rdata[29]), .Z(_zy_simnet_tvar_257[2]));
Q_AN02 U3264 ( .A0(n3), .A1(cddip0_out_ia_rdata[30]), .Z(_zy_simnet_tvar_257[1]));
Q_AN02 U3265 ( .A0(n3), .A1(cddip0_out_ia_rdata[31]), .Z(_zy_simnet_tvar_257[0]));
Q_AN02 U3266 ( .A0(n3), .A1(cddip0_out_ia_rdata[32]), .Z(_zy_simnet_tvar_258[31]));
Q_AN02 U3267 ( .A0(n3), .A1(cddip0_out_ia_rdata[33]), .Z(_zy_simnet_tvar_258[30]));
Q_AN02 U3268 ( .A0(n3), .A1(cddip0_out_ia_rdata[34]), .Z(_zy_simnet_tvar_258[29]));
Q_AN02 U3269 ( .A0(n3), .A1(cddip0_out_ia_rdata[35]), .Z(_zy_simnet_tvar_258[28]));
Q_AN02 U3270 ( .A0(n3), .A1(cddip0_out_ia_rdata[36]), .Z(_zy_simnet_tvar_258[27]));
Q_AN02 U3271 ( .A0(n3), .A1(cddip0_out_ia_rdata[37]), .Z(_zy_simnet_tvar_258[26]));
Q_AN02 U3272 ( .A0(n3), .A1(cddip0_out_ia_rdata[38]), .Z(_zy_simnet_tvar_258[25]));
Q_AN02 U3273 ( .A0(n3), .A1(cddip0_out_ia_rdata[39]), .Z(_zy_simnet_tvar_258[24]));
Q_AN02 U3274 ( .A0(n3), .A1(cddip0_out_ia_rdata[40]), .Z(_zy_simnet_tvar_258[23]));
Q_AN02 U3275 ( .A0(n3), .A1(cddip0_out_ia_rdata[41]), .Z(_zy_simnet_tvar_258[22]));
Q_AN02 U3276 ( .A0(n3), .A1(cddip0_out_ia_rdata[42]), .Z(_zy_simnet_tvar_258[21]));
Q_AN02 U3277 ( .A0(n3), .A1(cddip0_out_ia_rdata[43]), .Z(_zy_simnet_tvar_258[20]));
Q_AN02 U3278 ( .A0(n3), .A1(cddip0_out_ia_rdata[44]), .Z(_zy_simnet_tvar_258[19]));
Q_AN02 U3279 ( .A0(n3), .A1(cddip0_out_ia_rdata[45]), .Z(_zy_simnet_tvar_258[18]));
Q_AN02 U3280 ( .A0(n3), .A1(cddip0_out_ia_rdata[46]), .Z(_zy_simnet_tvar_258[17]));
Q_AN02 U3281 ( .A0(n3), .A1(cddip0_out_ia_rdata[47]), .Z(_zy_simnet_tvar_258[16]));
Q_AN02 U3282 ( .A0(n3), .A1(cddip0_out_ia_rdata[48]), .Z(_zy_simnet_tvar_258[15]));
Q_AN02 U3283 ( .A0(n3), .A1(cddip0_out_ia_rdata[49]), .Z(_zy_simnet_tvar_258[14]));
Q_AN02 U3284 ( .A0(n3), .A1(cddip0_out_ia_rdata[50]), .Z(_zy_simnet_tvar_258[13]));
Q_AN02 U3285 ( .A0(n3), .A1(cddip0_out_ia_rdata[51]), .Z(_zy_simnet_tvar_258[12]));
Q_AN02 U3286 ( .A0(n3), .A1(cddip0_out_ia_rdata[52]), .Z(_zy_simnet_tvar_258[11]));
Q_AN02 U3287 ( .A0(n3), .A1(cddip0_out_ia_rdata[53]), .Z(_zy_simnet_tvar_258[10]));
Q_AN02 U3288 ( .A0(n3), .A1(cddip0_out_ia_rdata[54]), .Z(_zy_simnet_tvar_258[9]));
Q_AN02 U3289 ( .A0(n3), .A1(cddip0_out_ia_rdata[55]), .Z(_zy_simnet_tvar_258[8]));
Q_AN02 U3290 ( .A0(n3), .A1(cddip0_out_ia_rdata[56]), .Z(_zy_simnet_tvar_258[7]));
Q_AN02 U3291 ( .A0(n3), .A1(cddip0_out_ia_rdata[57]), .Z(_zy_simnet_tvar_258[6]));
Q_AN02 U3292 ( .A0(n3), .A1(cddip0_out_ia_rdata[58]), .Z(_zy_simnet_tvar_258[5]));
Q_AN02 U3293 ( .A0(n3), .A1(cddip0_out_ia_rdata[59]), .Z(_zy_simnet_tvar_258[4]));
Q_AN02 U3294 ( .A0(n3), .A1(cddip0_out_ia_rdata[60]), .Z(_zy_simnet_tvar_258[3]));
Q_AN02 U3295 ( .A0(n3), .A1(cddip0_out_ia_rdata[61]), .Z(_zy_simnet_tvar_258[2]));
Q_AN02 U3296 ( .A0(n3), .A1(cddip0_out_ia_rdata[62]), .Z(_zy_simnet_tvar_258[1]));
Q_AN02 U3297 ( .A0(n3), .A1(cddip0_out_ia_rdata[63]), .Z(_zy_simnet_tvar_258[0]));
Q_AN02 U3298 ( .A0(n3), .A1(cddip0_out_ia_rdata[64]), .Z(_zy_simnet_tvar_259[31]));
Q_AN02 U3299 ( .A0(n3), .A1(cddip0_out_ia_rdata[65]), .Z(_zy_simnet_tvar_259[30]));
Q_AN02 U3300 ( .A0(n3), .A1(cddip0_out_ia_rdata[66]), .Z(_zy_simnet_tvar_259[29]));
Q_AN02 U3301 ( .A0(n3), .A1(cddip0_out_ia_rdata[67]), .Z(_zy_simnet_tvar_259[28]));
Q_AN02 U3302 ( .A0(n3), .A1(cddip0_out_ia_rdata[68]), .Z(_zy_simnet_tvar_259[27]));
Q_AN02 U3303 ( .A0(n3), .A1(cddip0_out_ia_rdata[69]), .Z(_zy_simnet_tvar_259[26]));
Q_AN02 U3304 ( .A0(n3), .A1(cddip0_out_ia_rdata[70]), .Z(_zy_simnet_tvar_259[25]));
Q_AN02 U3305 ( .A0(n3), .A1(cddip0_out_ia_rdata[71]), .Z(_zy_simnet_tvar_259[24]));
Q_AN02 U3306 ( .A0(n3), .A1(cddip0_out_ia_rdata[72]), .Z(_zy_simnet_tvar_259[23]));
Q_AN02 U3307 ( .A0(n3), .A1(cddip0_out_ia_rdata[73]), .Z(_zy_simnet_tvar_259[22]));
Q_AN02 U3308 ( .A0(n3), .A1(cddip0_out_ia_rdata[74]), .Z(_zy_simnet_tvar_259[21]));
Q_AN02 U3309 ( .A0(n3), .A1(cddip0_out_ia_rdata[75]), .Z(_zy_simnet_tvar_259[20]));
Q_AN02 U3310 ( .A0(n3), .A1(cddip0_out_ia_rdata[76]), .Z(_zy_simnet_tvar_259[19]));
Q_AN02 U3311 ( .A0(n3), .A1(cddip0_out_ia_rdata[77]), .Z(_zy_simnet_tvar_259[18]));
Q_AN02 U3312 ( .A0(n3), .A1(cddip0_out_ia_rdata[78]), .Z(_zy_simnet_tvar_259[17]));
Q_AN02 U3313 ( .A0(n3), .A1(cddip0_out_ia_rdata[79]), .Z(_zy_simnet_tvar_259[16]));
Q_AN02 U3314 ( .A0(n3), .A1(cddip0_out_ia_rdata[80]), .Z(_zy_simnet_tvar_259[15]));
Q_AN02 U3315 ( .A0(n3), .A1(cddip0_out_ia_rdata[81]), .Z(_zy_simnet_tvar_259[14]));
Q_AN02 U3316 ( .A0(n3), .A1(cddip0_out_ia_rdata[82]), .Z(_zy_simnet_tvar_259[13]));
Q_AN02 U3317 ( .A0(n3), .A1(cddip0_out_ia_rdata[83]), .Z(_zy_simnet_tvar_259[12]));
Q_AN02 U3318 ( .A0(n3), .A1(cddip0_out_ia_rdata[84]), .Z(_zy_simnet_tvar_259[11]));
Q_AN02 U3319 ( .A0(n3), .A1(cddip0_out_ia_rdata[85]), .Z(_zy_simnet_tvar_259[10]));
Q_AN02 U3320 ( .A0(n3), .A1(cddip0_out_ia_rdata[86]), .Z(_zy_simnet_tvar_259[9]));
Q_AN02 U3321 ( .A0(n3), .A1(cddip0_out_ia_rdata[87]), .Z(_zy_simnet_tvar_259[8]));
Q_AN02 U3322 ( .A0(n3), .A1(cddip0_out_ia_rdata[88]), .Z(_zy_simnet_tvar_259[7]));
Q_AN02 U3323 ( .A0(n3), .A1(cddip0_out_ia_rdata[89]), .Z(_zy_simnet_tvar_259[6]));
Q_AN02 U3324 ( .A0(n3), .A1(cddip0_out_ia_rdata[90]), .Z(_zy_simnet_tvar_259[5]));
Q_AN02 U3325 ( .A0(n3), .A1(cddip0_out_ia_rdata[91]), .Z(_zy_simnet_tvar_259[4]));
Q_AN02 U3326 ( .A0(n3), .A1(cddip0_out_ia_rdata[92]), .Z(_zy_simnet_tvar_259[3]));
Q_AN02 U3327 ( .A0(n3), .A1(cddip0_out_ia_rdata[93]), .Z(_zy_simnet_tvar_259[2]));
Q_AN02 U3328 ( .A0(n3), .A1(cddip0_out_ia_rdata[94]), .Z(_zy_simnet_tvar_259[1]));
Q_AN02 U3329 ( .A0(n3), .A1(cddip0_out_ia_rdata[95]), .Z(_zy_simnet_tvar_259[0]));
Q_AN02 U3330 ( .A0(n3), .A1(cddip1_out_ia_rdata[0]), .Z(_zy_simnet_tvar_264[31]));
Q_AN02 U3331 ( .A0(n3), .A1(cddip1_out_ia_rdata[1]), .Z(_zy_simnet_tvar_264[30]));
Q_AN02 U3332 ( .A0(n3), .A1(cddip1_out_ia_rdata[2]), .Z(_zy_simnet_tvar_264[29]));
Q_AN02 U3333 ( .A0(n3), .A1(cddip1_out_ia_rdata[3]), .Z(_zy_simnet_tvar_264[28]));
Q_AN02 U3334 ( .A0(n3), .A1(cddip1_out_ia_rdata[4]), .Z(_zy_simnet_tvar_264[27]));
Q_AN02 U3335 ( .A0(n3), .A1(cddip1_out_ia_rdata[5]), .Z(_zy_simnet_tvar_264[26]));
Q_AN02 U3336 ( .A0(n3), .A1(cddip1_out_ia_rdata[6]), .Z(_zy_simnet_tvar_264[25]));
Q_AN02 U3337 ( .A0(n3), .A1(cddip1_out_ia_rdata[7]), .Z(_zy_simnet_tvar_264[24]));
Q_AN02 U3338 ( .A0(n3), .A1(cddip1_out_ia_rdata[8]), .Z(_zy_simnet_tvar_264[23]));
Q_AN02 U3339 ( .A0(n3), .A1(cddip1_out_ia_rdata[9]), .Z(_zy_simnet_tvar_264[22]));
Q_AN02 U3340 ( .A0(n3), .A1(cddip1_out_ia_rdata[10]), .Z(_zy_simnet_tvar_264[21]));
Q_AN02 U3341 ( .A0(n3), .A1(cddip1_out_ia_rdata[11]), .Z(_zy_simnet_tvar_264[20]));
Q_AN02 U3342 ( .A0(n3), .A1(cddip1_out_ia_rdata[12]), .Z(_zy_simnet_tvar_264[19]));
Q_AN02 U3343 ( .A0(n3), .A1(cddip1_out_ia_rdata[13]), .Z(_zy_simnet_tvar_264[18]));
Q_AN02 U3344 ( .A0(n3), .A1(cddip1_out_ia_rdata[14]), .Z(_zy_simnet_tvar_264[17]));
Q_AN02 U3345 ( .A0(n3), .A1(cddip1_out_ia_rdata[15]), .Z(_zy_simnet_tvar_264[16]));
Q_AN02 U3346 ( .A0(n3), .A1(cddip1_out_ia_rdata[16]), .Z(_zy_simnet_tvar_264[15]));
Q_AN02 U3347 ( .A0(n3), .A1(cddip1_out_ia_rdata[17]), .Z(_zy_simnet_tvar_264[14]));
Q_AN02 U3348 ( .A0(n3), .A1(cddip1_out_ia_rdata[18]), .Z(_zy_simnet_tvar_264[13]));
Q_AN02 U3349 ( .A0(n3), .A1(cddip1_out_ia_rdata[19]), .Z(_zy_simnet_tvar_264[12]));
Q_AN02 U3350 ( .A0(n3), .A1(cddip1_out_ia_rdata[20]), .Z(_zy_simnet_tvar_264[11]));
Q_AN02 U3351 ( .A0(n3), .A1(cddip1_out_ia_rdata[21]), .Z(_zy_simnet_tvar_264[10]));
Q_AN02 U3352 ( .A0(n3), .A1(cddip1_out_ia_rdata[22]), .Z(_zy_simnet_tvar_264[9]));
Q_AN02 U3353 ( .A0(n3), .A1(cddip1_out_ia_rdata[23]), .Z(_zy_simnet_tvar_264[8]));
Q_AN02 U3354 ( .A0(n3), .A1(cddip1_out_ia_rdata[24]), .Z(_zy_simnet_tvar_264[7]));
Q_AN02 U3355 ( .A0(n3), .A1(cddip1_out_ia_rdata[25]), .Z(_zy_simnet_tvar_264[6]));
Q_AN02 U3356 ( .A0(n3), .A1(cddip1_out_ia_rdata[26]), .Z(_zy_simnet_tvar_264[5]));
Q_AN02 U3357 ( .A0(n3), .A1(cddip1_out_ia_rdata[27]), .Z(_zy_simnet_tvar_264[4]));
Q_AN02 U3358 ( .A0(n3), .A1(cddip1_out_ia_rdata[28]), .Z(_zy_simnet_tvar_264[3]));
Q_AN02 U3359 ( .A0(n3), .A1(cddip1_out_ia_rdata[29]), .Z(_zy_simnet_tvar_264[2]));
Q_AN02 U3360 ( .A0(n3), .A1(cddip1_out_ia_rdata[30]), .Z(_zy_simnet_tvar_264[1]));
Q_AN02 U3361 ( .A0(n3), .A1(cddip1_out_ia_rdata[31]), .Z(_zy_simnet_tvar_264[0]));
Q_AN02 U3362 ( .A0(n3), .A1(cddip1_out_ia_rdata[32]), .Z(_zy_simnet_tvar_265[31]));
Q_AN02 U3363 ( .A0(n3), .A1(cddip1_out_ia_rdata[33]), .Z(_zy_simnet_tvar_265[30]));
Q_AN02 U3364 ( .A0(n3), .A1(cddip1_out_ia_rdata[34]), .Z(_zy_simnet_tvar_265[29]));
Q_AN02 U3365 ( .A0(n3), .A1(cddip1_out_ia_rdata[35]), .Z(_zy_simnet_tvar_265[28]));
Q_AN02 U3366 ( .A0(n3), .A1(cddip1_out_ia_rdata[36]), .Z(_zy_simnet_tvar_265[27]));
Q_AN02 U3367 ( .A0(n3), .A1(cddip1_out_ia_rdata[37]), .Z(_zy_simnet_tvar_265[26]));
Q_AN02 U3368 ( .A0(n3), .A1(cddip1_out_ia_rdata[38]), .Z(_zy_simnet_tvar_265[25]));
Q_AN02 U3369 ( .A0(n3), .A1(cddip1_out_ia_rdata[39]), .Z(_zy_simnet_tvar_265[24]));
Q_AN02 U3370 ( .A0(n3), .A1(cddip1_out_ia_rdata[40]), .Z(_zy_simnet_tvar_265[23]));
Q_AN02 U3371 ( .A0(n3), .A1(cddip1_out_ia_rdata[41]), .Z(_zy_simnet_tvar_265[22]));
Q_AN02 U3372 ( .A0(n3), .A1(cddip1_out_ia_rdata[42]), .Z(_zy_simnet_tvar_265[21]));
Q_AN02 U3373 ( .A0(n3), .A1(cddip1_out_ia_rdata[43]), .Z(_zy_simnet_tvar_265[20]));
Q_AN02 U3374 ( .A0(n3), .A1(cddip1_out_ia_rdata[44]), .Z(_zy_simnet_tvar_265[19]));
Q_AN02 U3375 ( .A0(n3), .A1(cddip1_out_ia_rdata[45]), .Z(_zy_simnet_tvar_265[18]));
Q_AN02 U3376 ( .A0(n3), .A1(cddip1_out_ia_rdata[46]), .Z(_zy_simnet_tvar_265[17]));
Q_AN02 U3377 ( .A0(n3), .A1(cddip1_out_ia_rdata[47]), .Z(_zy_simnet_tvar_265[16]));
Q_AN02 U3378 ( .A0(n3), .A1(cddip1_out_ia_rdata[48]), .Z(_zy_simnet_tvar_265[15]));
Q_AN02 U3379 ( .A0(n3), .A1(cddip1_out_ia_rdata[49]), .Z(_zy_simnet_tvar_265[14]));
Q_AN02 U3380 ( .A0(n3), .A1(cddip1_out_ia_rdata[50]), .Z(_zy_simnet_tvar_265[13]));
Q_AN02 U3381 ( .A0(n3), .A1(cddip1_out_ia_rdata[51]), .Z(_zy_simnet_tvar_265[12]));
Q_AN02 U3382 ( .A0(n3), .A1(cddip1_out_ia_rdata[52]), .Z(_zy_simnet_tvar_265[11]));
Q_AN02 U3383 ( .A0(n3), .A1(cddip1_out_ia_rdata[53]), .Z(_zy_simnet_tvar_265[10]));
Q_AN02 U3384 ( .A0(n3), .A1(cddip1_out_ia_rdata[54]), .Z(_zy_simnet_tvar_265[9]));
Q_AN02 U3385 ( .A0(n3), .A1(cddip1_out_ia_rdata[55]), .Z(_zy_simnet_tvar_265[8]));
Q_AN02 U3386 ( .A0(n3), .A1(cddip1_out_ia_rdata[56]), .Z(_zy_simnet_tvar_265[7]));
Q_AN02 U3387 ( .A0(n3), .A1(cddip1_out_ia_rdata[57]), .Z(_zy_simnet_tvar_265[6]));
Q_AN02 U3388 ( .A0(n3), .A1(cddip1_out_ia_rdata[58]), .Z(_zy_simnet_tvar_265[5]));
Q_AN02 U3389 ( .A0(n3), .A1(cddip1_out_ia_rdata[59]), .Z(_zy_simnet_tvar_265[4]));
Q_AN02 U3390 ( .A0(n3), .A1(cddip1_out_ia_rdata[60]), .Z(_zy_simnet_tvar_265[3]));
Q_AN02 U3391 ( .A0(n3), .A1(cddip1_out_ia_rdata[61]), .Z(_zy_simnet_tvar_265[2]));
Q_AN02 U3392 ( .A0(n3), .A1(cddip1_out_ia_rdata[62]), .Z(_zy_simnet_tvar_265[1]));
Q_AN02 U3393 ( .A0(n3), .A1(cddip1_out_ia_rdata[63]), .Z(_zy_simnet_tvar_265[0]));
Q_AN02 U3394 ( .A0(n3), .A1(cddip1_out_ia_rdata[64]), .Z(_zy_simnet_tvar_266[31]));
Q_AN02 U3395 ( .A0(n3), .A1(cddip1_out_ia_rdata[65]), .Z(_zy_simnet_tvar_266[30]));
Q_AN02 U3396 ( .A0(n3), .A1(cddip1_out_ia_rdata[66]), .Z(_zy_simnet_tvar_266[29]));
Q_AN02 U3397 ( .A0(n3), .A1(cddip1_out_ia_rdata[67]), .Z(_zy_simnet_tvar_266[28]));
Q_AN02 U3398 ( .A0(n3), .A1(cddip1_out_ia_rdata[68]), .Z(_zy_simnet_tvar_266[27]));
Q_AN02 U3399 ( .A0(n3), .A1(cddip1_out_ia_rdata[69]), .Z(_zy_simnet_tvar_266[26]));
Q_AN02 U3400 ( .A0(n3), .A1(cddip1_out_ia_rdata[70]), .Z(_zy_simnet_tvar_266[25]));
Q_AN02 U3401 ( .A0(n3), .A1(cddip1_out_ia_rdata[71]), .Z(_zy_simnet_tvar_266[24]));
Q_AN02 U3402 ( .A0(n3), .A1(cddip1_out_ia_rdata[72]), .Z(_zy_simnet_tvar_266[23]));
Q_AN02 U3403 ( .A0(n3), .A1(cddip1_out_ia_rdata[73]), .Z(_zy_simnet_tvar_266[22]));
Q_AN02 U3404 ( .A0(n3), .A1(cddip1_out_ia_rdata[74]), .Z(_zy_simnet_tvar_266[21]));
Q_AN02 U3405 ( .A0(n3), .A1(cddip1_out_ia_rdata[75]), .Z(_zy_simnet_tvar_266[20]));
Q_AN02 U3406 ( .A0(n3), .A1(cddip1_out_ia_rdata[76]), .Z(_zy_simnet_tvar_266[19]));
Q_AN02 U3407 ( .A0(n3), .A1(cddip1_out_ia_rdata[77]), .Z(_zy_simnet_tvar_266[18]));
Q_AN02 U3408 ( .A0(n3), .A1(cddip1_out_ia_rdata[78]), .Z(_zy_simnet_tvar_266[17]));
Q_AN02 U3409 ( .A0(n3), .A1(cddip1_out_ia_rdata[79]), .Z(_zy_simnet_tvar_266[16]));
Q_AN02 U3410 ( .A0(n3), .A1(cddip1_out_ia_rdata[80]), .Z(_zy_simnet_tvar_266[15]));
Q_AN02 U3411 ( .A0(n3), .A1(cddip1_out_ia_rdata[81]), .Z(_zy_simnet_tvar_266[14]));
Q_AN02 U3412 ( .A0(n3), .A1(cddip1_out_ia_rdata[82]), .Z(_zy_simnet_tvar_266[13]));
Q_AN02 U3413 ( .A0(n3), .A1(cddip1_out_ia_rdata[83]), .Z(_zy_simnet_tvar_266[12]));
Q_AN02 U3414 ( .A0(n3), .A1(cddip1_out_ia_rdata[84]), .Z(_zy_simnet_tvar_266[11]));
Q_AN02 U3415 ( .A0(n3), .A1(cddip1_out_ia_rdata[85]), .Z(_zy_simnet_tvar_266[10]));
Q_AN02 U3416 ( .A0(n3), .A1(cddip1_out_ia_rdata[86]), .Z(_zy_simnet_tvar_266[9]));
Q_AN02 U3417 ( .A0(n3), .A1(cddip1_out_ia_rdata[87]), .Z(_zy_simnet_tvar_266[8]));
Q_AN02 U3418 ( .A0(n3), .A1(cddip1_out_ia_rdata[88]), .Z(_zy_simnet_tvar_266[7]));
Q_AN02 U3419 ( .A0(n3), .A1(cddip1_out_ia_rdata[89]), .Z(_zy_simnet_tvar_266[6]));
Q_AN02 U3420 ( .A0(n3), .A1(cddip1_out_ia_rdata[90]), .Z(_zy_simnet_tvar_266[5]));
Q_AN02 U3421 ( .A0(n3), .A1(cddip1_out_ia_rdata[91]), .Z(_zy_simnet_tvar_266[4]));
Q_AN02 U3422 ( .A0(n3), .A1(cddip1_out_ia_rdata[92]), .Z(_zy_simnet_tvar_266[3]));
Q_AN02 U3423 ( .A0(n3), .A1(cddip1_out_ia_rdata[93]), .Z(_zy_simnet_tvar_266[2]));
Q_AN02 U3424 ( .A0(n3), .A1(cddip1_out_ia_rdata[94]), .Z(_zy_simnet_tvar_266[1]));
Q_AN02 U3425 ( .A0(n3), .A1(cddip1_out_ia_rdata[95]), .Z(_zy_simnet_tvar_266[0]));
Q_AN02 U3426 ( .A0(n3), .A1(cddip2_out_ia_rdata[0]), .Z(_zy_simnet_tvar_271[31]));
Q_AN02 U3427 ( .A0(n3), .A1(cddip2_out_ia_rdata[1]), .Z(_zy_simnet_tvar_271[30]));
Q_AN02 U3428 ( .A0(n3), .A1(cddip2_out_ia_rdata[2]), .Z(_zy_simnet_tvar_271[29]));
Q_AN02 U3429 ( .A0(n3), .A1(cddip2_out_ia_rdata[3]), .Z(_zy_simnet_tvar_271[28]));
Q_AN02 U3430 ( .A0(n3), .A1(cddip2_out_ia_rdata[4]), .Z(_zy_simnet_tvar_271[27]));
Q_AN02 U3431 ( .A0(n3), .A1(cddip2_out_ia_rdata[5]), .Z(_zy_simnet_tvar_271[26]));
Q_AN02 U3432 ( .A0(n3), .A1(cddip2_out_ia_rdata[6]), .Z(_zy_simnet_tvar_271[25]));
Q_AN02 U3433 ( .A0(n3), .A1(cddip2_out_ia_rdata[7]), .Z(_zy_simnet_tvar_271[24]));
Q_AN02 U3434 ( .A0(n3), .A1(cddip2_out_ia_rdata[8]), .Z(_zy_simnet_tvar_271[23]));
Q_AN02 U3435 ( .A0(n3), .A1(cddip2_out_ia_rdata[9]), .Z(_zy_simnet_tvar_271[22]));
Q_AN02 U3436 ( .A0(n3), .A1(cddip2_out_ia_rdata[10]), .Z(_zy_simnet_tvar_271[21]));
Q_AN02 U3437 ( .A0(n3), .A1(cddip2_out_ia_rdata[11]), .Z(_zy_simnet_tvar_271[20]));
Q_AN02 U3438 ( .A0(n3), .A1(cddip2_out_ia_rdata[12]), .Z(_zy_simnet_tvar_271[19]));
Q_AN02 U3439 ( .A0(n3), .A1(cddip2_out_ia_rdata[13]), .Z(_zy_simnet_tvar_271[18]));
Q_AN02 U3440 ( .A0(n3), .A1(cddip2_out_ia_rdata[14]), .Z(_zy_simnet_tvar_271[17]));
Q_AN02 U3441 ( .A0(n3), .A1(cddip2_out_ia_rdata[15]), .Z(_zy_simnet_tvar_271[16]));
Q_AN02 U3442 ( .A0(n3), .A1(cddip2_out_ia_rdata[16]), .Z(_zy_simnet_tvar_271[15]));
Q_AN02 U3443 ( .A0(n3), .A1(cddip2_out_ia_rdata[17]), .Z(_zy_simnet_tvar_271[14]));
Q_AN02 U3444 ( .A0(n3), .A1(cddip2_out_ia_rdata[18]), .Z(_zy_simnet_tvar_271[13]));
Q_AN02 U3445 ( .A0(n3), .A1(cddip2_out_ia_rdata[19]), .Z(_zy_simnet_tvar_271[12]));
Q_AN02 U3446 ( .A0(n3), .A1(cddip2_out_ia_rdata[20]), .Z(_zy_simnet_tvar_271[11]));
Q_AN02 U3447 ( .A0(n3), .A1(cddip2_out_ia_rdata[21]), .Z(_zy_simnet_tvar_271[10]));
Q_AN02 U3448 ( .A0(n3), .A1(cddip2_out_ia_rdata[22]), .Z(_zy_simnet_tvar_271[9]));
Q_AN02 U3449 ( .A0(n3), .A1(cddip2_out_ia_rdata[23]), .Z(_zy_simnet_tvar_271[8]));
Q_AN02 U3450 ( .A0(n3), .A1(cddip2_out_ia_rdata[24]), .Z(_zy_simnet_tvar_271[7]));
Q_AN02 U3451 ( .A0(n3), .A1(cddip2_out_ia_rdata[25]), .Z(_zy_simnet_tvar_271[6]));
Q_AN02 U3452 ( .A0(n3), .A1(cddip2_out_ia_rdata[26]), .Z(_zy_simnet_tvar_271[5]));
Q_AN02 U3453 ( .A0(n3), .A1(cddip2_out_ia_rdata[27]), .Z(_zy_simnet_tvar_271[4]));
Q_AN02 U3454 ( .A0(n3), .A1(cddip2_out_ia_rdata[28]), .Z(_zy_simnet_tvar_271[3]));
Q_AN02 U3455 ( .A0(n3), .A1(cddip2_out_ia_rdata[29]), .Z(_zy_simnet_tvar_271[2]));
Q_AN02 U3456 ( .A0(n3), .A1(cddip2_out_ia_rdata[30]), .Z(_zy_simnet_tvar_271[1]));
Q_AN02 U3457 ( .A0(n3), .A1(cddip2_out_ia_rdata[31]), .Z(_zy_simnet_tvar_271[0]));
Q_AN02 U3458 ( .A0(n3), .A1(cddip2_out_ia_rdata[32]), .Z(_zy_simnet_tvar_272[31]));
Q_AN02 U3459 ( .A0(n3), .A1(cddip2_out_ia_rdata[33]), .Z(_zy_simnet_tvar_272[30]));
Q_AN02 U3460 ( .A0(n3), .A1(cddip2_out_ia_rdata[34]), .Z(_zy_simnet_tvar_272[29]));
Q_AN02 U3461 ( .A0(n3), .A1(cddip2_out_ia_rdata[35]), .Z(_zy_simnet_tvar_272[28]));
Q_AN02 U3462 ( .A0(n3), .A1(cddip2_out_ia_rdata[36]), .Z(_zy_simnet_tvar_272[27]));
Q_AN02 U3463 ( .A0(n3), .A1(cddip2_out_ia_rdata[37]), .Z(_zy_simnet_tvar_272[26]));
Q_AN02 U3464 ( .A0(n3), .A1(cddip2_out_ia_rdata[38]), .Z(_zy_simnet_tvar_272[25]));
Q_AN02 U3465 ( .A0(n3), .A1(cddip2_out_ia_rdata[39]), .Z(_zy_simnet_tvar_272[24]));
Q_AN02 U3466 ( .A0(n3), .A1(cddip2_out_ia_rdata[40]), .Z(_zy_simnet_tvar_272[23]));
Q_AN02 U3467 ( .A0(n3), .A1(cddip2_out_ia_rdata[41]), .Z(_zy_simnet_tvar_272[22]));
Q_AN02 U3468 ( .A0(n3), .A1(cddip2_out_ia_rdata[42]), .Z(_zy_simnet_tvar_272[21]));
Q_AN02 U3469 ( .A0(n3), .A1(cddip2_out_ia_rdata[43]), .Z(_zy_simnet_tvar_272[20]));
Q_AN02 U3470 ( .A0(n3), .A1(cddip2_out_ia_rdata[44]), .Z(_zy_simnet_tvar_272[19]));
Q_AN02 U3471 ( .A0(n3), .A1(cddip2_out_ia_rdata[45]), .Z(_zy_simnet_tvar_272[18]));
Q_AN02 U3472 ( .A0(n3), .A1(cddip2_out_ia_rdata[46]), .Z(_zy_simnet_tvar_272[17]));
Q_AN02 U3473 ( .A0(n3), .A1(cddip2_out_ia_rdata[47]), .Z(_zy_simnet_tvar_272[16]));
Q_AN02 U3474 ( .A0(n3), .A1(cddip2_out_ia_rdata[48]), .Z(_zy_simnet_tvar_272[15]));
Q_AN02 U3475 ( .A0(n3), .A1(cddip2_out_ia_rdata[49]), .Z(_zy_simnet_tvar_272[14]));
Q_AN02 U3476 ( .A0(n3), .A1(cddip2_out_ia_rdata[50]), .Z(_zy_simnet_tvar_272[13]));
Q_AN02 U3477 ( .A0(n3), .A1(cddip2_out_ia_rdata[51]), .Z(_zy_simnet_tvar_272[12]));
Q_AN02 U3478 ( .A0(n3), .A1(cddip2_out_ia_rdata[52]), .Z(_zy_simnet_tvar_272[11]));
Q_AN02 U3479 ( .A0(n3), .A1(cddip2_out_ia_rdata[53]), .Z(_zy_simnet_tvar_272[10]));
Q_AN02 U3480 ( .A0(n3), .A1(cddip2_out_ia_rdata[54]), .Z(_zy_simnet_tvar_272[9]));
Q_AN02 U3481 ( .A0(n3), .A1(cddip2_out_ia_rdata[55]), .Z(_zy_simnet_tvar_272[8]));
Q_AN02 U3482 ( .A0(n3), .A1(cddip2_out_ia_rdata[56]), .Z(_zy_simnet_tvar_272[7]));
Q_AN02 U3483 ( .A0(n3), .A1(cddip2_out_ia_rdata[57]), .Z(_zy_simnet_tvar_272[6]));
Q_AN02 U3484 ( .A0(n3), .A1(cddip2_out_ia_rdata[58]), .Z(_zy_simnet_tvar_272[5]));
Q_AN02 U3485 ( .A0(n3), .A1(cddip2_out_ia_rdata[59]), .Z(_zy_simnet_tvar_272[4]));
Q_AN02 U3486 ( .A0(n3), .A1(cddip2_out_ia_rdata[60]), .Z(_zy_simnet_tvar_272[3]));
Q_AN02 U3487 ( .A0(n3), .A1(cddip2_out_ia_rdata[61]), .Z(_zy_simnet_tvar_272[2]));
Q_AN02 U3488 ( .A0(n3), .A1(cddip2_out_ia_rdata[62]), .Z(_zy_simnet_tvar_272[1]));
Q_AN02 U3489 ( .A0(n3), .A1(cddip2_out_ia_rdata[63]), .Z(_zy_simnet_tvar_272[0]));
Q_AN02 U3490 ( .A0(n3), .A1(cddip2_out_ia_rdata[64]), .Z(_zy_simnet_tvar_273[31]));
Q_AN02 U3491 ( .A0(n3), .A1(cddip2_out_ia_rdata[65]), .Z(_zy_simnet_tvar_273[30]));
Q_AN02 U3492 ( .A0(n3), .A1(cddip2_out_ia_rdata[66]), .Z(_zy_simnet_tvar_273[29]));
Q_AN02 U3493 ( .A0(n3), .A1(cddip2_out_ia_rdata[67]), .Z(_zy_simnet_tvar_273[28]));
Q_AN02 U3494 ( .A0(n3), .A1(cddip2_out_ia_rdata[68]), .Z(_zy_simnet_tvar_273[27]));
Q_AN02 U3495 ( .A0(n3), .A1(cddip2_out_ia_rdata[69]), .Z(_zy_simnet_tvar_273[26]));
Q_AN02 U3496 ( .A0(n3), .A1(cddip2_out_ia_rdata[70]), .Z(_zy_simnet_tvar_273[25]));
Q_AN02 U3497 ( .A0(n3), .A1(cddip2_out_ia_rdata[71]), .Z(_zy_simnet_tvar_273[24]));
Q_AN02 U3498 ( .A0(n3), .A1(cddip2_out_ia_rdata[72]), .Z(_zy_simnet_tvar_273[23]));
Q_AN02 U3499 ( .A0(n3), .A1(cddip2_out_ia_rdata[73]), .Z(_zy_simnet_tvar_273[22]));
Q_AN02 U3500 ( .A0(n3), .A1(cddip2_out_ia_rdata[74]), .Z(_zy_simnet_tvar_273[21]));
Q_AN02 U3501 ( .A0(n3), .A1(cddip2_out_ia_rdata[75]), .Z(_zy_simnet_tvar_273[20]));
Q_AN02 U3502 ( .A0(n3), .A1(cddip2_out_ia_rdata[76]), .Z(_zy_simnet_tvar_273[19]));
Q_AN02 U3503 ( .A0(n3), .A1(cddip2_out_ia_rdata[77]), .Z(_zy_simnet_tvar_273[18]));
Q_AN02 U3504 ( .A0(n3), .A1(cddip2_out_ia_rdata[78]), .Z(_zy_simnet_tvar_273[17]));
Q_AN02 U3505 ( .A0(n3), .A1(cddip2_out_ia_rdata[79]), .Z(_zy_simnet_tvar_273[16]));
Q_AN02 U3506 ( .A0(n3), .A1(cddip2_out_ia_rdata[80]), .Z(_zy_simnet_tvar_273[15]));
Q_AN02 U3507 ( .A0(n3), .A1(cddip2_out_ia_rdata[81]), .Z(_zy_simnet_tvar_273[14]));
Q_AN02 U3508 ( .A0(n3), .A1(cddip2_out_ia_rdata[82]), .Z(_zy_simnet_tvar_273[13]));
Q_AN02 U3509 ( .A0(n3), .A1(cddip2_out_ia_rdata[83]), .Z(_zy_simnet_tvar_273[12]));
Q_AN02 U3510 ( .A0(n3), .A1(cddip2_out_ia_rdata[84]), .Z(_zy_simnet_tvar_273[11]));
Q_AN02 U3511 ( .A0(n3), .A1(cddip2_out_ia_rdata[85]), .Z(_zy_simnet_tvar_273[10]));
Q_AN02 U3512 ( .A0(n3), .A1(cddip2_out_ia_rdata[86]), .Z(_zy_simnet_tvar_273[9]));
Q_AN02 U3513 ( .A0(n3), .A1(cddip2_out_ia_rdata[87]), .Z(_zy_simnet_tvar_273[8]));
Q_AN02 U3514 ( .A0(n3), .A1(cddip2_out_ia_rdata[88]), .Z(_zy_simnet_tvar_273[7]));
Q_AN02 U3515 ( .A0(n3), .A1(cddip2_out_ia_rdata[89]), .Z(_zy_simnet_tvar_273[6]));
Q_AN02 U3516 ( .A0(n3), .A1(cddip2_out_ia_rdata[90]), .Z(_zy_simnet_tvar_273[5]));
Q_AN02 U3517 ( .A0(n3), .A1(cddip2_out_ia_rdata[91]), .Z(_zy_simnet_tvar_273[4]));
Q_AN02 U3518 ( .A0(n3), .A1(cddip2_out_ia_rdata[92]), .Z(_zy_simnet_tvar_273[3]));
Q_AN02 U3519 ( .A0(n3), .A1(cddip2_out_ia_rdata[93]), .Z(_zy_simnet_tvar_273[2]));
Q_AN02 U3520 ( .A0(n3), .A1(cddip2_out_ia_rdata[94]), .Z(_zy_simnet_tvar_273[1]));
Q_AN02 U3521 ( .A0(n3), .A1(cddip2_out_ia_rdata[95]), .Z(_zy_simnet_tvar_273[0]));
Q_AN02 U3522 ( .A0(n3), .A1(cddip3_out_ia_rdata[0]), .Z(_zy_simnet_tvar_278[31]));
Q_AN02 U3523 ( .A0(n3), .A1(cddip3_out_ia_rdata[1]), .Z(_zy_simnet_tvar_278[30]));
Q_AN02 U3524 ( .A0(n3), .A1(cddip3_out_ia_rdata[2]), .Z(_zy_simnet_tvar_278[29]));
Q_AN02 U3525 ( .A0(n3), .A1(cddip3_out_ia_rdata[3]), .Z(_zy_simnet_tvar_278[28]));
Q_AN02 U3526 ( .A0(n3), .A1(cddip3_out_ia_rdata[4]), .Z(_zy_simnet_tvar_278[27]));
Q_AN02 U3527 ( .A0(n3), .A1(cddip3_out_ia_rdata[5]), .Z(_zy_simnet_tvar_278[26]));
Q_AN02 U3528 ( .A0(n3), .A1(cddip3_out_ia_rdata[6]), .Z(_zy_simnet_tvar_278[25]));
Q_AN02 U3529 ( .A0(n3), .A1(cddip3_out_ia_rdata[7]), .Z(_zy_simnet_tvar_278[24]));
Q_AN02 U3530 ( .A0(n3), .A1(cddip3_out_ia_rdata[8]), .Z(_zy_simnet_tvar_278[23]));
Q_AN02 U3531 ( .A0(n3), .A1(cddip3_out_ia_rdata[9]), .Z(_zy_simnet_tvar_278[22]));
Q_AN02 U3532 ( .A0(n3), .A1(cddip3_out_ia_rdata[10]), .Z(_zy_simnet_tvar_278[21]));
Q_AN02 U3533 ( .A0(n3), .A1(cddip3_out_ia_rdata[11]), .Z(_zy_simnet_tvar_278[20]));
Q_AN02 U3534 ( .A0(n3), .A1(cddip3_out_ia_rdata[12]), .Z(_zy_simnet_tvar_278[19]));
Q_AN02 U3535 ( .A0(n3), .A1(cddip3_out_ia_rdata[13]), .Z(_zy_simnet_tvar_278[18]));
Q_AN02 U3536 ( .A0(n3), .A1(cddip3_out_ia_rdata[14]), .Z(_zy_simnet_tvar_278[17]));
Q_AN02 U3537 ( .A0(n3), .A1(cddip3_out_ia_rdata[15]), .Z(_zy_simnet_tvar_278[16]));
Q_AN02 U3538 ( .A0(n3), .A1(cddip3_out_ia_rdata[16]), .Z(_zy_simnet_tvar_278[15]));
Q_AN02 U3539 ( .A0(n3), .A1(cddip3_out_ia_rdata[17]), .Z(_zy_simnet_tvar_278[14]));
Q_AN02 U3540 ( .A0(n3), .A1(cddip3_out_ia_rdata[18]), .Z(_zy_simnet_tvar_278[13]));
Q_AN02 U3541 ( .A0(n3), .A1(cddip3_out_ia_rdata[19]), .Z(_zy_simnet_tvar_278[12]));
Q_AN02 U3542 ( .A0(n3), .A1(cddip3_out_ia_rdata[20]), .Z(_zy_simnet_tvar_278[11]));
Q_AN02 U3543 ( .A0(n3), .A1(cddip3_out_ia_rdata[21]), .Z(_zy_simnet_tvar_278[10]));
Q_AN02 U3544 ( .A0(n3), .A1(cddip3_out_ia_rdata[22]), .Z(_zy_simnet_tvar_278[9]));
Q_AN02 U3545 ( .A0(n3), .A1(cddip3_out_ia_rdata[23]), .Z(_zy_simnet_tvar_278[8]));
Q_AN02 U3546 ( .A0(n3), .A1(cddip3_out_ia_rdata[24]), .Z(_zy_simnet_tvar_278[7]));
Q_AN02 U3547 ( .A0(n3), .A1(cddip3_out_ia_rdata[25]), .Z(_zy_simnet_tvar_278[6]));
Q_AN02 U3548 ( .A0(n3), .A1(cddip3_out_ia_rdata[26]), .Z(_zy_simnet_tvar_278[5]));
Q_AN02 U3549 ( .A0(n3), .A1(cddip3_out_ia_rdata[27]), .Z(_zy_simnet_tvar_278[4]));
Q_AN02 U3550 ( .A0(n3), .A1(cddip3_out_ia_rdata[28]), .Z(_zy_simnet_tvar_278[3]));
Q_AN02 U3551 ( .A0(n3), .A1(cddip3_out_ia_rdata[29]), .Z(_zy_simnet_tvar_278[2]));
Q_AN02 U3552 ( .A0(n3), .A1(cddip3_out_ia_rdata[30]), .Z(_zy_simnet_tvar_278[1]));
Q_AN02 U3553 ( .A0(n3), .A1(cddip3_out_ia_rdata[31]), .Z(_zy_simnet_tvar_278[0]));
Q_AN02 U3554 ( .A0(n3), .A1(cddip3_out_ia_rdata[32]), .Z(_zy_simnet_tvar_279[31]));
Q_AN02 U3555 ( .A0(n3), .A1(cddip3_out_ia_rdata[33]), .Z(_zy_simnet_tvar_279[30]));
Q_AN02 U3556 ( .A0(n3), .A1(cddip3_out_ia_rdata[34]), .Z(_zy_simnet_tvar_279[29]));
Q_AN02 U3557 ( .A0(n3), .A1(cddip3_out_ia_rdata[35]), .Z(_zy_simnet_tvar_279[28]));
Q_AN02 U3558 ( .A0(n3), .A1(cddip3_out_ia_rdata[36]), .Z(_zy_simnet_tvar_279[27]));
Q_AN02 U3559 ( .A0(n3), .A1(cddip3_out_ia_rdata[37]), .Z(_zy_simnet_tvar_279[26]));
Q_AN02 U3560 ( .A0(n3), .A1(cddip3_out_ia_rdata[38]), .Z(_zy_simnet_tvar_279[25]));
Q_AN02 U3561 ( .A0(n3), .A1(cddip3_out_ia_rdata[39]), .Z(_zy_simnet_tvar_279[24]));
Q_AN02 U3562 ( .A0(n3), .A1(cddip3_out_ia_rdata[40]), .Z(_zy_simnet_tvar_279[23]));
Q_AN02 U3563 ( .A0(n3), .A1(cddip3_out_ia_rdata[41]), .Z(_zy_simnet_tvar_279[22]));
Q_AN02 U3564 ( .A0(n3), .A1(cddip3_out_ia_rdata[42]), .Z(_zy_simnet_tvar_279[21]));
Q_AN02 U3565 ( .A0(n3), .A1(cddip3_out_ia_rdata[43]), .Z(_zy_simnet_tvar_279[20]));
Q_AN02 U3566 ( .A0(n3), .A1(cddip3_out_ia_rdata[44]), .Z(_zy_simnet_tvar_279[19]));
Q_AN02 U3567 ( .A0(n3), .A1(cddip3_out_ia_rdata[45]), .Z(_zy_simnet_tvar_279[18]));
Q_AN02 U3568 ( .A0(n3), .A1(cddip3_out_ia_rdata[46]), .Z(_zy_simnet_tvar_279[17]));
Q_AN02 U3569 ( .A0(n3), .A1(cddip3_out_ia_rdata[47]), .Z(_zy_simnet_tvar_279[16]));
Q_AN02 U3570 ( .A0(n3), .A1(cddip3_out_ia_rdata[48]), .Z(_zy_simnet_tvar_279[15]));
Q_AN02 U3571 ( .A0(n3), .A1(cddip3_out_ia_rdata[49]), .Z(_zy_simnet_tvar_279[14]));
Q_AN02 U3572 ( .A0(n3), .A1(cddip3_out_ia_rdata[50]), .Z(_zy_simnet_tvar_279[13]));
Q_AN02 U3573 ( .A0(n3), .A1(cddip3_out_ia_rdata[51]), .Z(_zy_simnet_tvar_279[12]));
Q_AN02 U3574 ( .A0(n3), .A1(cddip3_out_ia_rdata[52]), .Z(_zy_simnet_tvar_279[11]));
Q_AN02 U3575 ( .A0(n3), .A1(cddip3_out_ia_rdata[53]), .Z(_zy_simnet_tvar_279[10]));
Q_AN02 U3576 ( .A0(n3), .A1(cddip3_out_ia_rdata[54]), .Z(_zy_simnet_tvar_279[9]));
Q_AN02 U3577 ( .A0(n3), .A1(cddip3_out_ia_rdata[55]), .Z(_zy_simnet_tvar_279[8]));
Q_AN02 U3578 ( .A0(n3), .A1(cddip3_out_ia_rdata[56]), .Z(_zy_simnet_tvar_279[7]));
Q_AN02 U3579 ( .A0(n3), .A1(cddip3_out_ia_rdata[57]), .Z(_zy_simnet_tvar_279[6]));
Q_AN02 U3580 ( .A0(n3), .A1(cddip3_out_ia_rdata[58]), .Z(_zy_simnet_tvar_279[5]));
Q_AN02 U3581 ( .A0(n3), .A1(cddip3_out_ia_rdata[59]), .Z(_zy_simnet_tvar_279[4]));
Q_AN02 U3582 ( .A0(n3), .A1(cddip3_out_ia_rdata[60]), .Z(_zy_simnet_tvar_279[3]));
Q_AN02 U3583 ( .A0(n3), .A1(cddip3_out_ia_rdata[61]), .Z(_zy_simnet_tvar_279[2]));
Q_AN02 U3584 ( .A0(n3), .A1(cddip3_out_ia_rdata[62]), .Z(_zy_simnet_tvar_279[1]));
Q_AN02 U3585 ( .A0(n3), .A1(cddip3_out_ia_rdata[63]), .Z(_zy_simnet_tvar_279[0]));
Q_AN02 U3586 ( .A0(n3), .A1(cddip3_out_ia_rdata[64]), .Z(_zy_simnet_tvar_280[31]));
Q_AN02 U3587 ( .A0(n3), .A1(cddip3_out_ia_rdata[65]), .Z(_zy_simnet_tvar_280[30]));
Q_AN02 U3588 ( .A0(n3), .A1(cddip3_out_ia_rdata[66]), .Z(_zy_simnet_tvar_280[29]));
Q_AN02 U3589 ( .A0(n3), .A1(cddip3_out_ia_rdata[67]), .Z(_zy_simnet_tvar_280[28]));
Q_AN02 U3590 ( .A0(n3), .A1(cddip3_out_ia_rdata[68]), .Z(_zy_simnet_tvar_280[27]));
Q_AN02 U3591 ( .A0(n3), .A1(cddip3_out_ia_rdata[69]), .Z(_zy_simnet_tvar_280[26]));
Q_AN02 U3592 ( .A0(n3), .A1(cddip3_out_ia_rdata[70]), .Z(_zy_simnet_tvar_280[25]));
Q_AN02 U3593 ( .A0(n3), .A1(cddip3_out_ia_rdata[71]), .Z(_zy_simnet_tvar_280[24]));
Q_AN02 U3594 ( .A0(n3), .A1(cddip3_out_ia_rdata[72]), .Z(_zy_simnet_tvar_280[23]));
Q_AN02 U3595 ( .A0(n3), .A1(cddip3_out_ia_rdata[73]), .Z(_zy_simnet_tvar_280[22]));
Q_AN02 U3596 ( .A0(n3), .A1(cddip3_out_ia_rdata[74]), .Z(_zy_simnet_tvar_280[21]));
Q_AN02 U3597 ( .A0(n3), .A1(cddip3_out_ia_rdata[75]), .Z(_zy_simnet_tvar_280[20]));
Q_AN02 U3598 ( .A0(n3), .A1(cddip3_out_ia_rdata[76]), .Z(_zy_simnet_tvar_280[19]));
Q_AN02 U3599 ( .A0(n3), .A1(cddip3_out_ia_rdata[77]), .Z(_zy_simnet_tvar_280[18]));
Q_AN02 U3600 ( .A0(n3), .A1(cddip3_out_ia_rdata[78]), .Z(_zy_simnet_tvar_280[17]));
Q_AN02 U3601 ( .A0(n3), .A1(cddip3_out_ia_rdata[79]), .Z(_zy_simnet_tvar_280[16]));
Q_AN02 U3602 ( .A0(n3), .A1(cddip3_out_ia_rdata[80]), .Z(_zy_simnet_tvar_280[15]));
Q_AN02 U3603 ( .A0(n3), .A1(cddip3_out_ia_rdata[81]), .Z(_zy_simnet_tvar_280[14]));
Q_AN02 U3604 ( .A0(n3), .A1(cddip3_out_ia_rdata[82]), .Z(_zy_simnet_tvar_280[13]));
Q_AN02 U3605 ( .A0(n3), .A1(cddip3_out_ia_rdata[83]), .Z(_zy_simnet_tvar_280[12]));
Q_AN02 U3606 ( .A0(n3), .A1(cddip3_out_ia_rdata[84]), .Z(_zy_simnet_tvar_280[11]));
Q_AN02 U3607 ( .A0(n3), .A1(cddip3_out_ia_rdata[85]), .Z(_zy_simnet_tvar_280[10]));
Q_AN02 U3608 ( .A0(n3), .A1(cddip3_out_ia_rdata[86]), .Z(_zy_simnet_tvar_280[9]));
Q_AN02 U3609 ( .A0(n3), .A1(cddip3_out_ia_rdata[87]), .Z(_zy_simnet_tvar_280[8]));
Q_AN02 U3610 ( .A0(n3), .A1(cddip3_out_ia_rdata[88]), .Z(_zy_simnet_tvar_280[7]));
Q_AN02 U3611 ( .A0(n3), .A1(cddip3_out_ia_rdata[89]), .Z(_zy_simnet_tvar_280[6]));
Q_AN02 U3612 ( .A0(n3), .A1(cddip3_out_ia_rdata[90]), .Z(_zy_simnet_tvar_280[5]));
Q_AN02 U3613 ( .A0(n3), .A1(cddip3_out_ia_rdata[91]), .Z(_zy_simnet_tvar_280[4]));
Q_AN02 U3614 ( .A0(n3), .A1(cddip3_out_ia_rdata[92]), .Z(_zy_simnet_tvar_280[3]));
Q_AN02 U3615 ( .A0(n3), .A1(cddip3_out_ia_rdata[93]), .Z(_zy_simnet_tvar_280[2]));
Q_AN02 U3616 ( .A0(n3), .A1(cddip3_out_ia_rdata[94]), .Z(_zy_simnet_tvar_280[1]));
Q_AN02 U3617 ( .A0(n3), .A1(cddip3_out_ia_rdata[95]), .Z(_zy_simnet_tvar_280[0]));
Q_MX02 U3618 ( .S(tready_override[0]), .A0(kme_cceip0_ob_in[0]), .A1(o_tready_override_val), .Z(_zy_simnet_tvar_351));
Q_MX02 U3619 ( .S(tready_override[1]), .A0(kme_cceip1_ob_in[0]), .A1(o_tready_override_val), .Z(_zy_simnet_tvar_356));
Q_MX02 U3620 ( .S(tready_override[2]), .A0(kme_cceip2_ob_in[0]), .A1(o_tready_override_val), .Z(_zy_simnet_tvar_361));
Q_MX02 U3621 ( .S(tready_override[3]), .A0(kme_cceip3_ob_in[0]), .A1(o_tready_override_val), .Z(_zy_simnet_tvar_366));
Q_MX02 U3622 ( .S(tready_override[4]), .A0(kme_cddip0_ob_in[0]), .A1(o_tready_override_val), .Z(_zy_simnet_tvar_371));
Q_MX02 U3623 ( .S(tready_override[5]), .A0(kme_cddip1_ob_in[0]), .A1(o_tready_override_val), .Z(_zy_simnet_tvar_376));
Q_MX02 U3624 ( .S(tready_override[6]), .A0(kme_cddip2_ob_in[0]), .A1(o_tready_override_val), .Z(_zy_simnet_tvar_381));
Q_MX02 U3625 ( .S(tready_override[7]), .A0(kme_cddip3_ob_in[0]), .A1(o_tready_override_val), .Z(_zy_simnet_tvar_386));
Q_INV U3626 ( .A(reg_addr[0]), .Z(n4));
Q_INV U3627 ( .A(reg_addr[1]), .Z(n5));
Q_INV U3628 ( .A(reg_addr[2]), .Z(n6));
Q_INV U3629 ( .A(reg_addr[3]), .Z(n7));
Q_INV U3630 ( .A(reg_addr[10]), .Z(n8));
Q_AN03 U3631 ( .A0(n8), .A1(reg_addr[9]), .A2(reg_addr[8]), .Z(n9));
Q_AN03 U3632 ( .A0(reg_addr[7]), .A1(reg_addr[6]), .A2(reg_addr[5]), .Z(n10));
Q_AN03 U3633 ( .A0(reg_addr[4]), .A1(n7), .A2(n6), .Z(n11));
Q_AN03 U3634 ( .A0(n5), .A1(n4), .A2(n9), .Z(n12));
Q_AN03 U3635 ( .A0(n10), .A1(n11), .A2(n12), .Z(n13));
Q_AN02 U3636 ( .A0(wr_stb), .A1(n13), .Z(n30));
Q_FDP1 \im_consumed_kme_cceip0_REG[1] ( .CK(clk), .R(rst_n), .D(n29), .Q(im_consumed_kme_cceip0[1]), .QN( ));
Q_FDP1 \im_consumed_kme_cceip0_REG[0] ( .CK(clk), .R(rst_n), .D(n28), .Q(im_consumed_kme_cceip0[0]), .QN( ));
Q_FDP1 \im_consumed_kme_cddip0_REG[1] ( .CK(clk), .R(rst_n), .D(n27), .Q(im_consumed_kme_cddip0[1]), .QN( ));
Q_FDP1 \im_consumed_kme_cddip0_REG[0] ( .CK(clk), .R(rst_n), .D(n26), .Q(im_consumed_kme_cddip0[0]), .QN( ));
Q_FDP1 \im_consumed_kme_cceip1_REG[1] ( .CK(clk), .R(rst_n), .D(n25), .Q(im_consumed_kme_cceip1[1]), .QN( ));
Q_FDP1 \im_consumed_kme_cceip1_REG[0] ( .CK(clk), .R(rst_n), .D(n24), .Q(im_consumed_kme_cceip1[0]), .QN( ));
Q_FDP1 \im_consumed_kme_cddip1_REG[1] ( .CK(clk), .R(rst_n), .D(n23), .Q(im_consumed_kme_cddip1[1]), .QN( ));
Q_FDP1 \im_consumed_kme_cddip1_REG[0] ( .CK(clk), .R(rst_n), .D(n22), .Q(im_consumed_kme_cddip1[0]), .QN( ));
Q_FDP1 \im_consumed_kme_cceip2_REG[1] ( .CK(clk), .R(rst_n), .D(n21), .Q(im_consumed_kme_cceip2[1]), .QN( ));
Q_FDP1 \im_consumed_kme_cceip2_REG[0] ( .CK(clk), .R(rst_n), .D(n20), .Q(im_consumed_kme_cceip2[0]), .QN( ));
Q_FDP1 \im_consumed_kme_cddip2_REG[1] ( .CK(clk), .R(rst_n), .D(n19), .Q(im_consumed_kme_cddip2[1]), .QN( ));
Q_FDP1 \im_consumed_kme_cddip2_REG[0] ( .CK(clk), .R(rst_n), .D(n18), .Q(im_consumed_kme_cddip2[0]), .QN( ));
Q_FDP1 \im_consumed_kme_cceip3_REG[1] ( .CK(clk), .R(rst_n), .D(n17), .Q(im_consumed_kme_cceip3[1]), .QN( ));
Q_FDP1 \im_consumed_kme_cceip3_REG[0] ( .CK(clk), .R(rst_n), .D(n16), .Q(im_consumed_kme_cceip3[0]), .QN( ));
Q_FDP1 \im_consumed_kme_cddip3_REG[1] ( .CK(clk), .R(rst_n), .D(n15), .Q(im_consumed_kme_cddip3[1]), .QN( ));
Q_FDP1 \im_consumed_kme_cddip3_REG[0] ( .CK(clk), .R(rst_n), .D(n14), .Q(im_consumed_kme_cddip3[0]), .QN( ));
Q_AN02 U3653 ( .A0(n30), .A1(wr_data[14]), .Z(n14));
Q_AN02 U3654 ( .A0(n30), .A1(wr_data[15]), .Z(n15));
Q_AN02 U3655 ( .A0(n30), .A1(wr_data[6]), .Z(n16));
Q_AN02 U3656 ( .A0(n30), .A1(wr_data[7]), .Z(n17));
Q_AN02 U3657 ( .A0(n30), .A1(wr_data[12]), .Z(n18));
Q_AN02 U3658 ( .A0(n30), .A1(wr_data[13]), .Z(n19));
Q_AN02 U3659 ( .A0(n30), .A1(wr_data[4]), .Z(n20));
Q_AN02 U3660 ( .A0(n30), .A1(wr_data[5]), .Z(n21));
Q_AN02 U3661 ( .A0(n30), .A1(wr_data[10]), .Z(n22));
Q_AN02 U3662 ( .A0(n30), .A1(wr_data[11]), .Z(n23));
Q_AN02 U3663 ( .A0(n30), .A1(wr_data[2]), .Z(n24));
Q_AN02 U3664 ( .A0(n30), .A1(wr_data[3]), .Z(n25));
Q_AN02 U3665 ( .A0(n30), .A1(wr_data[8]), .Z(n26));
Q_AN02 U3666 ( .A0(n30), .A1(wr_data[9]), .Z(n27));
Q_AN02 U3667 ( .A0(n30), .A1(wr_data[0]), .Z(n28));
Q_AN02 U3668 ( .A0(n30), .A1(wr_data[1]), .Z(n29));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "labels (2,0) 1 271 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m2 "sa_ctrl 1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m3 "sa_ctrl_rst_dat 1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "3"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\rbus_ring_o.addr  (1,0) 1 15 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\rbus_ring_o.wr_data  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\rbus_ring_o.rd_data  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\kme_cceip0_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\kme_cceip0_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\kme_cceip0_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\kme_cceip0_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\kme_cceip1_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\kme_cceip1_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\kme_cceip1_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\kme_cceip1_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\kme_cceip2_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\kme_cceip2_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\kme_cceip2_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\kme_cceip2_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\kme_cceip3_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\kme_cceip3_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\kme_cceip3_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\kme_cceip3_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\kme_cddip0_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\kme_cddip0_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\kme_cddip0_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\kme_cddip0_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\kme_cddip1_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\kme_cddip1_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\kme_cddip1_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\kme_cddip1_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\kme_cddip2_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\kme_cddip2_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\kme_cddip2_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\kme_cddip2_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\kme_cddip3_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\kme_cddip3_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\kme_cddip3_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\kme_cddip3_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\kim_dout.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\kim_dout.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\kim_dout.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m39 "\kim_dout.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m40 "\kim_dout.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m41 "\kim_dout.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m42 "\kim_dout.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m43 "\labels%s.guid_size  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m44 "\labels%s.label_size  1 5 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m45 "\labels%s.label  1 255 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m46 "\labels%s.delimiter_valid  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m47 "\labels%s.delimiter  1 7 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m48 "\tready_override.r.part0  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m49 "\cceip_encrypt_kop_fifo_override.r.part0  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m50 "\cceip_validate_kop_fifo_override.r.part0  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m51 "\cddip_decrypt_kop_fifo_override.r.part0  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m52 "\sa_global_ctrl.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m53 "\sa_global_ctrl.f.spare  (1,0) 1 29 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m54 "\sa_ctrl%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m55 "\sa_ctrl%s.f.spare  1 26 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m56 "\sa_ctrl%s.f.sa_event_sel  1 4 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m57 "\rbus_ring_i.addr  (1,0) 1 15 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m58 "\rbus_ring_i.wr_data  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m59 "\rbus_ring_i.rd_data  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m60 "\kme_cceip0_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m61 "\kme_cceip0_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m62 "\kme_cceip0_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m63 "\kme_cceip0_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m64 "\kme_cceip1_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m65 "\kme_cceip1_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m66 "\kme_cceip1_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m67 "\kme_cceip1_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m68 "\kme_cceip2_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m69 "\kme_cceip2_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m70 "\kme_cceip2_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m71 "\kme_cceip2_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m72 "\kme_cceip3_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m73 "\kme_cceip3_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m74 "\kme_cceip3_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m75 "\kme_cceip3_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m76 "\kme_cddip0_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m77 "\kme_cddip0_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m78 "\kme_cddip0_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m79 "\kme_cddip0_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m80 "\kme_cddip1_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m81 "\kme_cddip1_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m82 "\kme_cddip1_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m83 "\kme_cddip1_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m84 "\kme_cddip2_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m85 "\kme_cddip2_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m86 "\kme_cddip2_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m87 "\kme_cddip2_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m88 "\kme_cddip3_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m89 "\kme_cddip3_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m90 "\kme_cddip3_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m91 "\kme_cddip3_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m92 "\idle_components.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m93 "\idle_components.f.num_key_tlvs_in_flight  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m94 "\sa_snapshot%s.r.part1  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m95 "\sa_snapshot%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m96 "\sa_snapshot%s.f.unused  1 13 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m97 "\sa_snapshot%s.f.upper  1 17 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m98 "\sa_snapshot%s.f.lower  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m99 "sa_snapshot 1 63 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m100 "\sa_count%s.r.part1  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m101 "\sa_count%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m102 "\sa_count%s.f.unused  1 13 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m103 "\sa_count%s.f.upper  1 17 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m104 "\sa_count%s.f.lower  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m105 "sa_count 1 63 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m106 "\ckv_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m107 "\ckv_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m108 "\ckv_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m109 "\ckv_ia_status.r.part0  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m110 "\ckv_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m111 "\ckv_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m112 "\ckv_ia_status.f.addr  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m113 "\kim_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m114 "\kim_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m115 "\kim_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m116 "\kim_ia_status.r.part0  (1,0) 1 21 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m117 "\kim_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m118 "\kim_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m119 "\kim_ia_status.f.addr  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m120 "\spare.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m121 "\spare.f.spare  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m122 "\cceip0_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m123 "\cceip0_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m124 "\cceip0_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m125 "\cceip0_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m126 "\cceip0_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m127 "\cceip0_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m128 "\cceip0_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m129 "\cceip0_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m130 "\cceip0_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m131 "\cceip0_out_ia_config.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m132 "\cceip0_out_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m133 "\cceip0_out_ia_config.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m134 "\cceip0_out_ia_rdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m135 "\cceip0_out_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m136 "\cceip0_out_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m137 "\cceip0_out_ia_rdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m138 "\cceip0_out_ia_rdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m139 "\cceip0_out_ia_rdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m140 "\cceip0_out_ia_rdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m141 "\cceip0_out_ia_rdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m142 "\cceip0_out_ia_rdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m143 "\cceip0_out_ia_status.r.part0  (1,0) 1 16 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m144 "\cceip0_out_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m145 "\cceip0_out_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m146 "\cceip0_out_ia_status.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m147 "\cceip0_out_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m148 "\cceip0_out_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m149 "\cceip0_out_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m150 "\cceip0_out_im_status.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m151 "\cceip0_out_im_status.f.wr_pointer  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m152 "\cceip0_out_im_config.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m153 "\cceip0_out_im_config.f.mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m154 "\cceip0_out_im_config.f.wr_credit_config  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m155 "\cddip0_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m156 "\cddip0_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m157 "\cddip0_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m158 "\cddip0_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m159 "\cddip0_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m160 "\cddip0_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m161 "\cddip0_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m162 "\cddip0_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m163 "\cddip0_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m164 "\cddip0_out_ia_config.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m165 "\cddip0_out_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m166 "\cddip0_out_ia_config.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m167 "\cddip0_out_ia_rdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m168 "\cddip0_out_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m169 "\cddip0_out_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m170 "\cddip0_out_ia_rdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m171 "\cddip0_out_ia_rdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m172 "\cddip0_out_ia_rdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m173 "\cddip0_out_ia_rdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m174 "\cddip0_out_ia_rdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m175 "\cddip0_out_ia_rdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m176 "\cddip0_out_ia_status.r.part0  (1,0) 1 16 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m177 "\cddip0_out_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m178 "\cddip0_out_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m179 "\cddip0_out_ia_status.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m180 "\cddip0_out_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m181 "\cddip0_out_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m182 "\cddip0_out_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m183 "\cddip0_out_im_status.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m184 "\cddip0_out_im_status.f.wr_pointer  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m185 "\cddip0_out_im_config.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m186 "\cddip0_out_im_config.f.mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m187 "\cddip0_out_im_config.f.wr_credit_config  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m188 "\cceip1_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m189 "\cceip1_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m190 "\cceip1_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m191 "\cceip1_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m192 "\cceip1_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m193 "\cceip1_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m194 "\cceip1_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m195 "\cceip1_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m196 "\cceip1_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m197 "\cceip1_out_ia_config.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m198 "\cceip1_out_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m199 "\cceip1_out_ia_config.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m200 "\cceip1_out_ia_rdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m201 "\cceip1_out_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m202 "\cceip1_out_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m203 "\cceip1_out_ia_rdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m204 "\cceip1_out_ia_rdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m205 "\cceip1_out_ia_rdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m206 "\cceip1_out_ia_rdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m207 "\cceip1_out_ia_rdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m208 "\cceip1_out_ia_rdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m209 "\cceip1_out_ia_status.r.part0  (1,0) 1 16 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m210 "\cceip1_out_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m211 "\cceip1_out_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m212 "\cceip1_out_ia_status.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m213 "\cceip1_out_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m214 "\cceip1_out_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m215 "\cceip1_out_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m216 "\cceip1_out_im_status.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m217 "\cceip1_out_im_status.f.wr_pointer  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m218 "\cceip1_out_im_config.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m219 "\cceip1_out_im_config.f.mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m220 "\cceip1_out_im_config.f.wr_credit_config  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m221 "\cddip1_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m222 "\cddip1_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m223 "\cddip1_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m224 "\cddip1_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m225 "\cddip1_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m226 "\cddip1_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m227 "\cddip1_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m228 "\cddip1_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m229 "\cddip1_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m230 "\cddip1_out_ia_config.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m231 "\cddip1_out_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m232 "\cddip1_out_ia_config.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m233 "\cddip1_out_ia_rdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m234 "\cddip1_out_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m235 "\cddip1_out_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m236 "\cddip1_out_ia_rdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m237 "\cddip1_out_ia_rdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m238 "\cddip1_out_ia_rdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m239 "\cddip1_out_ia_rdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m240 "\cddip1_out_ia_rdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m241 "\cddip1_out_ia_rdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m242 "\cddip1_out_ia_status.r.part0  (1,0) 1 16 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m243 "\cddip1_out_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m244 "\cddip1_out_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m245 "\cddip1_out_ia_status.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m246 "\cddip1_out_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m247 "\cddip1_out_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m248 "\cddip1_out_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m249 "\cddip1_out_im_status.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m250 "\cddip1_out_im_status.f.wr_pointer  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m251 "\cddip1_out_im_config.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m252 "\cddip1_out_im_config.f.mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m253 "\cddip1_out_im_config.f.wr_credit_config  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m254 "\cceip2_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m255 "\cceip2_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m256 "\cceip2_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m257 "\cceip2_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m258 "\cceip2_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m259 "\cceip2_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m260 "\cceip2_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m261 "\cceip2_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m262 "\cceip2_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m263 "\cceip2_out_ia_config.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m264 "\cceip2_out_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m265 "\cceip2_out_ia_config.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m266 "\cceip2_out_ia_rdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m267 "\cceip2_out_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m268 "\cceip2_out_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m269 "\cceip2_out_ia_rdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m270 "\cceip2_out_ia_rdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m271 "\cceip2_out_ia_rdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m272 "\cceip2_out_ia_rdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m273 "\cceip2_out_ia_rdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m274 "\cceip2_out_ia_rdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m275 "\cceip2_out_ia_status.r.part0  (1,0) 1 16 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m276 "\cceip2_out_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m277 "\cceip2_out_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m278 "\cceip2_out_ia_status.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m279 "\cceip2_out_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m280 "\cceip2_out_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m281 "\cceip2_out_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m282 "\cceip2_out_im_status.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m283 "\cceip2_out_im_status.f.wr_pointer  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m284 "\cceip2_out_im_config.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m285 "\cceip2_out_im_config.f.mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m286 "\cceip2_out_im_config.f.wr_credit_config  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m287 "\cddip2_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m288 "\cddip2_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m289 "\cddip2_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m290 "\cddip2_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m291 "\cddip2_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m292 "\cddip2_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m293 "\cddip2_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m294 "\cddip2_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m295 "\cddip2_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m296 "\cddip2_out_ia_config.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m297 "\cddip2_out_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m298 "\cddip2_out_ia_config.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m299 "\cddip2_out_ia_rdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m300 "\cddip2_out_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m301 "\cddip2_out_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m302 "\cddip2_out_ia_rdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m303 "\cddip2_out_ia_rdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m304 "\cddip2_out_ia_rdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m305 "\cddip2_out_ia_rdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m306 "\cddip2_out_ia_rdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m307 "\cddip2_out_ia_rdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m308 "\cddip2_out_ia_status.r.part0  (1,0) 1 16 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m309 "\cddip2_out_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m310 "\cddip2_out_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m311 "\cddip2_out_ia_status.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m312 "\cddip2_out_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m313 "\cddip2_out_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m314 "\cddip2_out_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m315 "\cddip2_out_im_status.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m316 "\cddip2_out_im_status.f.wr_pointer  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m317 "\cddip2_out_im_config.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m318 "\cddip2_out_im_config.f.mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m319 "\cddip2_out_im_config.f.wr_credit_config  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m320 "\cceip3_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m321 "\cceip3_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m322 "\cceip3_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m323 "\cceip3_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m324 "\cceip3_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m325 "\cceip3_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m326 "\cceip3_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m327 "\cceip3_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m328 "\cceip3_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m329 "\cceip3_out_ia_config.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m330 "\cceip3_out_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m331 "\cceip3_out_ia_config.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m332 "\cceip3_out_ia_rdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m333 "\cceip3_out_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m334 "\cceip3_out_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m335 "\cceip3_out_ia_rdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m336 "\cceip3_out_ia_rdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m337 "\cceip3_out_ia_rdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m338 "\cceip3_out_ia_rdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m339 "\cceip3_out_ia_rdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m340 "\cceip3_out_ia_rdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m341 "\cceip3_out_ia_status.r.part0  (1,0) 1 16 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m342 "\cceip3_out_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m343 "\cceip3_out_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m344 "\cceip3_out_ia_status.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m345 "\cceip3_out_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m346 "\cceip3_out_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m347 "\cceip3_out_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m348 "\cceip3_out_im_status.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m349 "\cceip3_out_im_status.f.wr_pointer  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m350 "\cceip3_out_im_config.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m351 "\cceip3_out_im_config.f.mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m352 "\cceip3_out_im_config.f.wr_credit_config  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m353 "\cddip3_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m354 "\cddip3_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m355 "\cddip3_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m356 "\cddip3_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m357 "\cddip3_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m358 "\cddip3_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m359 "\cddip3_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m360 "\cddip3_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m361 "\cddip3_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m362 "\cddip3_out_ia_config.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m363 "\cddip3_out_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m364 "\cddip3_out_ia_config.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m365 "\cddip3_out_ia_rdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m366 "\cddip3_out_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m367 "\cddip3_out_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m368 "\cddip3_out_ia_rdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m369 "\cddip3_out_ia_rdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m370 "\cddip3_out_ia_rdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m371 "\cddip3_out_ia_rdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m372 "\cddip3_out_ia_rdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m373 "\cddip3_out_ia_rdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m374 "\cddip3_out_ia_status.r.part0  (1,0) 1 16 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m375 "\cddip3_out_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m376 "\cddip3_out_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m377 "\cddip3_out_ia_status.f.addr  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m378 "\cddip3_out_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m379 "\cddip3_out_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m380 "\cddip3_out_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m381 "\cddip3_out_im_status.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m382 "\cddip3_out_im_status.f.wr_pointer  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m383 "\cddip3_out_im_config.r.part0  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m384 "\cddip3_out_im_config.f.mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m385 "\cddip3_out_im_config.f.wr_credit_config  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m386 "\sa_snapshot_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m387 "\sa_snapshot_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m388 "\sa_snapshot_ia_wdata.f.unused  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m389 "\sa_snapshot_ia_wdata.f.upper  (1,0) 1 17 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m390 "\sa_snapshot_ia_wdata.f.lower  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m391 "\sa_snapshot_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m392 "\sa_snapshot_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m393 "\sa_snapshot_ia_rdata.f.unused  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m394 "\sa_snapshot_ia_rdata.f.upper  (1,0) 1 17 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m395 "\sa_snapshot_ia_rdata.f.lower  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m396 "\sa_snapshot_ia_config.r.part0  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m397 "\sa_snapshot_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m398 "\sa_snapshot_ia_config.f.addr  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m399 "\sa_snapshot_ia_status.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m400 "\sa_snapshot_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m401 "\sa_snapshot_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m402 "\sa_snapshot_ia_status.f.addr  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m403 "\sa_snapshot_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m404 "\sa_snapshot_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m405 "\sa_snapshot_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m406 "\sa_count_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m407 "\sa_count_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m408 "\sa_count_ia_wdata.f.unused  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m409 "\sa_count_ia_wdata.f.upper  (1,0) 1 17 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m410 "\sa_count_ia_wdata.f.lower  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m411 "\sa_count_ia_rdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m412 "\sa_count_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m413 "\sa_count_ia_rdata.f.unused  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m414 "\sa_count_ia_rdata.f.upper  (1,0) 1 17 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m415 "\sa_count_ia_rdata.f.lower  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m416 "\sa_count_ia_config.r.part0  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m417 "\sa_count_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m418 "\sa_count_ia_config.f.addr  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m419 "\sa_count_ia_status.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m420 "\sa_count_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m421 "\sa_count_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m422 "\sa_count_ia_status.f.addr  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m423 "\sa_count_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m424 "\sa_count_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m425 "\sa_count_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m426 "\sa_ctrl_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m427 "\sa_ctrl_ia_wdata.f.spare  (1,0) 1 26 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m428 "\sa_ctrl_ia_wdata.f.sa_event_sel  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m429 "\sa_ctrl_ia_rdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m430 "\sa_ctrl_ia_rdata.f.spare  (1,0) 1 26 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m431 "\sa_ctrl_ia_rdata.f.sa_event_sel  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m432 "\sa_ctrl_ia_config.r.part0  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m433 "\sa_ctrl_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m434 "\sa_ctrl_ia_config.f.addr  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m435 "\sa_ctrl_ia_status.r.part0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m436 "\sa_ctrl_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m437 "\sa_ctrl_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m438 "\sa_ctrl_ia_status.f.addr  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m439 "\sa_ctrl_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m440 "\sa_ctrl_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m441 "\sa_ctrl_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m442 "\sa_ctrl_rst_dat%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m443 "\sa_ctrl_rst_dat%s.f.spare  1 26 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m444 "\sa_ctrl_rst_dat%s.f.sa_event_sel  1 4 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m445 "\cceip0_im_din.data.data  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m446 "\cceip0_im_din.desc.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m447 "\cceip0_im_din.desc.im_meta  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m448 "\cddip0_im_din.data.data  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m449 "\cddip0_im_din.desc.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m450 "\cddip0_im_din.desc.im_meta  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m451 "\cceip1_im_din.data.data  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m452 "\cceip1_im_din.desc.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m453 "\cceip1_im_din.desc.im_meta  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m454 "\cddip1_im_din.data.data  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m455 "\cddip1_im_din.desc.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m456 "\cddip1_im_din.desc.im_meta  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m457 "\cceip2_im_din.data.data  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m458 "\cceip2_im_din.desc.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m459 "\cceip2_im_din.desc.im_meta  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m460 "\cddip2_im_din.data.data  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m461 "\cddip2_im_din.desc.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m462 "\cddip2_im_din.desc.im_meta  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m463 "\cceip3_im_din.data.data  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m464 "\cceip3_im_din.desc.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m465 "\cceip3_im_din.desc.im_meta  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m466 "\cddip3_im_din.data.data  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m467 "\cddip3_im_din.desc.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m468 "\cddip3_im_din.desc.im_meta  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m469 "\kme_cceip0_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m470 "\kme_cceip0_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m471 "\kme_cceip0_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m472 "\kme_cceip0_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m473 "\kme_cceip1_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m474 "\kme_cceip1_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m475 "\kme_cceip1_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m476 "\kme_cceip1_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m477 "\kme_cceip2_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m478 "\kme_cceip2_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m479 "\kme_cceip2_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m480 "\kme_cceip2_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m481 "\kme_cceip3_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m482 "\kme_cceip3_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m483 "\kme_cceip3_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m484 "\kme_cceip3_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m485 "\kme_cddip0_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m486 "\kme_cddip0_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m487 "\kme_cddip0_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m488 "\kme_cddip0_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m489 "\kme_cddip1_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m490 "\kme_cddip1_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m491 "\kme_cddip1_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m492 "\kme_cddip1_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m493 "\kme_cddip2_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m494 "\kme_cddip2_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m495 "\kme_cddip2_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m496 "\kme_cddip2_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m497 "\kme_cddip3_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m498 "\kme_cddip3_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m499 "\kme_cddip3_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m500 "\kme_cddip3_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m501 "\revid_wire.r.part0  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m502 "\revid_wire.f.revid  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "502"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "rbus_ring_o 7 \rbus_ring_o.addr  \rbus_ring_o.wr_strb  \rbus_ring_o.wr_data  \rbus_ring_o.rd_strb  \rbus_ring_o.rd_data  \rbus_ring_o.ack  \rbus_ring_o.err_ack "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "kme_cceip0_ob_out 6 \kme_cceip0_ob_out.tvalid  \kme_cceip0_ob_out.tlast  \kme_cceip0_ob_out.tid  \kme_cceip0_ob_out.tstrb  \kme_cceip0_ob_out.tuser  \kme_cceip0_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "kme_cceip0_ob_in_mod 1 \kme_cceip0_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "kme_cceip1_ob_out 6 \kme_cceip1_ob_out.tvalid  \kme_cceip1_ob_out.tlast  \kme_cceip1_ob_out.tid  \kme_cceip1_ob_out.tstrb  \kme_cceip1_ob_out.tuser  \kme_cceip1_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "kme_cceip1_ob_in_mod 1 \kme_cceip1_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "kme_cceip2_ob_out 6 \kme_cceip2_ob_out.tvalid  \kme_cceip2_ob_out.tlast  \kme_cceip2_ob_out.tid  \kme_cceip2_ob_out.tstrb  \kme_cceip2_ob_out.tuser  \kme_cceip2_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "kme_cceip2_ob_in_mod 1 \kme_cceip2_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r8 "kme_cceip3_ob_out 6 \kme_cceip3_ob_out.tvalid  \kme_cceip3_ob_out.tlast  \kme_cceip3_ob_out.tid  \kme_cceip3_ob_out.tstrb  \kme_cceip3_ob_out.tuser  \kme_cceip3_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r9 "kme_cceip3_ob_in_mod 1 \kme_cceip3_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r10 "kme_cddip0_ob_out 6 \kme_cddip0_ob_out.tvalid  \kme_cddip0_ob_out.tlast  \kme_cddip0_ob_out.tid  \kme_cddip0_ob_out.tstrb  \kme_cddip0_ob_out.tuser  \kme_cddip0_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r11 "kme_cddip0_ob_in_mod 1 \kme_cddip0_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r12 "kme_cddip1_ob_out 6 \kme_cddip1_ob_out.tvalid  \kme_cddip1_ob_out.tlast  \kme_cddip1_ob_out.tid  \kme_cddip1_ob_out.tstrb  \kme_cddip1_ob_out.tuser  \kme_cddip1_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r13 "kme_cddip1_ob_in_mod 1 \kme_cddip1_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r14 "kme_cddip2_ob_out 6 \kme_cddip2_ob_out.tvalid  \kme_cddip2_ob_out.tlast  \kme_cddip2_ob_out.tid  \kme_cddip2_ob_out.tstrb  \kme_cddip2_ob_out.tuser  \kme_cddip2_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r15 "kme_cddip2_ob_in_mod 1 \kme_cddip2_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r16 "kme_cddip3_ob_out 6 \kme_cddip3_ob_out.tvalid  \kme_cddip3_ob_out.tlast  \kme_cddip3_ob_out.tid  \kme_cddip3_ob_out.tstrb  \kme_cddip3_ob_out.tuser  \kme_cddip3_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r17 "kme_cddip3_ob_in_mod 1 \kme_cddip3_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r18 "kim_dout 7 \kim_dout.valid  \kim_dout.label_index  \kim_dout.ckv_length  \kim_dout.ckv_pointer  \kim_dout.pf_num  \kim_dout.vf_num  \kim_dout.vf_valid "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r19 "labels%s 5 \labels%s.guid_size  \labels%s.label_size  \labels%s.label  \labels%s.delimiter_valid  \labels%s.delimiter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r1 "tready_override 2 \tready_override.r  { \tready_override.r.part0  } \tready_override.f  { \tready_override.f.txc_tready_override  \tready_override.f.engine_7_tready_override  \tready_override.f.engine_6_tready_override  \tready_override.f.engine_5_tready_override  \tready_override.f.engine_4_tready_override  \tready_override.f.engine_3_tready_override  \tready_override.f.engine_2_tready_override  \tready_override.f.engine_1_tready_override  \tready_override.f.engine_0_tready_override  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r2 "cceip_encrypt_kop_fifo_override 2 \cceip_encrypt_kop_fifo_override.r  { \cceip_encrypt_kop_fifo_override.r.part0  } \cceip_encrypt_kop_fifo_override.f  { \cceip_encrypt_kop_fifo_override.f.gcm_status_data_fifo  \cceip_encrypt_kop_fifo_override.f.tlv_sb_data_fifo  \cceip_encrypt_kop_fifo_override.f.kdf_cmd_fifo  \cceip_encrypt_kop_fifo_override.f.kdfstream_cmd_fifo  \cceip_encrypt_kop_fifo_override.f.keyfilter_cmd_fifo  \cceip_encrypt_kop_fifo_override.f.gcm_tag_data_fifo  \cceip_encrypt_kop_fifo_override.f.gcm_cmd_fifo  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r3 "cceip_validate_kop_fifo_override 2 \cceip_validate_kop_fifo_override.r  { \cceip_validate_kop_fifo_override.r.part0  } \cceip_validate_kop_fifo_override.f  { \cceip_validate_kop_fifo_override.f.gcm_status_data_fifo  \cceip_validate_kop_fifo_override.f.tlv_sb_data_fifo  \cceip_validate_kop_fifo_override.f.kdf_cmd_fifo  \cceip_validate_kop_fifo_override.f.kdfstream_cmd_fifo  \cceip_validate_kop_fifo_override.f.keyfilter_cmd_fifo  \cceip_validate_kop_fifo_override.f.gcm_tag_data_fifo  \cceip_validate_kop_fifo_override.f.gcm_cmd_fifo  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r4 "cddip_decrypt_kop_fifo_override 2 \cddip_decrypt_kop_fifo_override.r  { \cddip_decrypt_kop_fifo_override.r.part0  } \cddip_decrypt_kop_fifo_override.f  { \cddip_decrypt_kop_fifo_override.f.gcm_status_data_fifo  \cddip_decrypt_kop_fifo_override.f.tlv_sb_data_fifo  \cddip_decrypt_kop_fifo_override.f.kdf_cmd_fifo  \cddip_decrypt_kop_fifo_override.f.kdfstream_cmd_fifo  \cddip_decrypt_kop_fifo_override.f.keyfilter_cmd_fifo  \cddip_decrypt_kop_fifo_override.f.gcm_tag_data_fifo  \cddip_decrypt_kop_fifo_override.f.gcm_cmd_fifo  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r5 "sa_global_ctrl 2 \sa_global_ctrl.r  { \sa_global_ctrl.r.part0  } \sa_global_ctrl.f  { \sa_global_ctrl.f.spare  \sa_global_ctrl.f.sa_snap  \sa_global_ctrl.f.sa_clear_live  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r6 "sa_ctrl%s 2 \sa_ctrl%s.r  { \sa_ctrl%s.r.part0  } \sa_ctrl%s.f  { \sa_ctrl%s.f.spare  \sa_ctrl%s.f.sa_event_sel  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r20 "rbus_ring_i 7 \rbus_ring_i.addr  \rbus_ring_i.wr_strb  \rbus_ring_i.wr_data  \rbus_ring_i.rd_strb  \rbus_ring_i.rd_data  \rbus_ring_i.ack  \rbus_ring_i.err_ack "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r21 "kme_cceip0_ob_out_pre 6 \kme_cceip0_ob_out_pre.tvalid  \kme_cceip0_ob_out_pre.tlast  \kme_cceip0_ob_out_pre.tid  \kme_cceip0_ob_out_pre.tstrb  \kme_cceip0_ob_out_pre.tuser  \kme_cceip0_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r22 "kme_cceip0_ob_in 1 \kme_cceip0_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r23 "kme_cceip1_ob_out_pre 6 \kme_cceip1_ob_out_pre.tvalid  \kme_cceip1_ob_out_pre.tlast  \kme_cceip1_ob_out_pre.tid  \kme_cceip1_ob_out_pre.tstrb  \kme_cceip1_ob_out_pre.tuser  \kme_cceip1_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r24 "kme_cceip1_ob_in 1 \kme_cceip1_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r25 "kme_cceip2_ob_out_pre 6 \kme_cceip2_ob_out_pre.tvalid  \kme_cceip2_ob_out_pre.tlast  \kme_cceip2_ob_out_pre.tid  \kme_cceip2_ob_out_pre.tstrb  \kme_cceip2_ob_out_pre.tuser  \kme_cceip2_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r26 "kme_cceip2_ob_in 1 \kme_cceip2_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r27 "kme_cceip3_ob_out_pre 6 \kme_cceip3_ob_out_pre.tvalid  \kme_cceip3_ob_out_pre.tlast  \kme_cceip3_ob_out_pre.tid  \kme_cceip3_ob_out_pre.tstrb  \kme_cceip3_ob_out_pre.tuser  \kme_cceip3_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r28 "kme_cceip3_ob_in 1 \kme_cceip3_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r29 "kme_cddip0_ob_out_pre 6 \kme_cddip0_ob_out_pre.tvalid  \kme_cddip0_ob_out_pre.tlast  \kme_cddip0_ob_out_pre.tid  \kme_cddip0_ob_out_pre.tstrb  \kme_cddip0_ob_out_pre.tuser  \kme_cddip0_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r30 "kme_cddip0_ob_in 1 \kme_cddip0_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r31 "kme_cddip1_ob_out_pre 6 \kme_cddip1_ob_out_pre.tvalid  \kme_cddip1_ob_out_pre.tlast  \kme_cddip1_ob_out_pre.tid  \kme_cddip1_ob_out_pre.tstrb  \kme_cddip1_ob_out_pre.tuser  \kme_cddip1_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r32 "kme_cddip1_ob_in 1 \kme_cddip1_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r33 "kme_cddip2_ob_out_pre 6 \kme_cddip2_ob_out_pre.tvalid  \kme_cddip2_ob_out_pre.tlast  \kme_cddip2_ob_out_pre.tid  \kme_cddip2_ob_out_pre.tstrb  \kme_cddip2_ob_out_pre.tuser  \kme_cddip2_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r34 "kme_cddip2_ob_in 1 \kme_cddip2_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r35 "kme_cddip3_ob_out_pre 6 \kme_cddip3_ob_out_pre.tvalid  \kme_cddip3_ob_out_pre.tlast  \kme_cddip3_ob_out_pre.tid  \kme_cddip3_ob_out_pre.tstrb  \kme_cddip3_ob_out_pre.tuser  \kme_cddip3_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r36 "kme_cddip3_ob_in 1 \kme_cddip3_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r7 "idle_components 2 \idle_components.r  { \idle_components.r.part0  } \idle_components.f  { \idle_components.f.num_key_tlvs_in_flight  \idle_components.f.cddip0_key_tlv_rsm_idle  \idle_components.f.cddip1_key_tlv_rsm_idle  \idle_components.f.cddip2_key_tlv_rsm_idle  \idle_components.f.cddip3_key_tlv_rsm_idle  \idle_components.f.cceip0_key_tlv_rsm_idle  \idle_components.f.cceip1_key_tlv_rsm_idle  \idle_components.f.cceip2_key_tlv_rsm_idle  \idle_components.f.cceip3_key_tlv_rsm_idle  \idle_components.f.no_key_tlv_in_flight  \idle_components.f.tlv_parser_idle  \idle_components.f.drng_idle  \idle_components.f.kme_slv_empty  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r8 "sa_snapshot%s 2 \sa_snapshot%s.r  { \sa_snapshot%s.r.part1  \sa_snapshot%s.r.part0  } \sa_snapshot%s.f  { \sa_snapshot%s.f.unused  \sa_snapshot%s.f.upper  \sa_snapshot%s.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r9 "sa_count%s 2 \sa_count%s.r  { \sa_count%s.r.part1  \sa_count%s.r.part0  } \sa_count%s.f  { \sa_count%s.f.unused  \sa_count%s.f.upper  \sa_count%s.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r10 "ckv_ia_capability 2 \ckv_ia_capability.r  { \ckv_ia_capability.r.part0  } \ckv_ia_capability.f  { \ckv_ia_capability.f.mem_type  \ckv_ia_capability.f.ack_error  \ckv_ia_capability.f.sim_tmo  \ckv_ia_capability.f.reserved_op  \ckv_ia_capability.f.compare  \ckv_ia_capability.f.set_init_start  \ckv_ia_capability.f.initialize_inc  \ckv_ia_capability.f.initialize  \ckv_ia_capability.f.reset  \ckv_ia_capability.f.disabled  \ckv_ia_capability.f.enable  \ckv_ia_capability.f.write  \ckv_ia_capability.f.read  \ckv_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r11 "ckv_ia_status 2 \ckv_ia_status.r  { \ckv_ia_status.r.part0  } \ckv_ia_status.f  { \ckv_ia_status.f.code  \ckv_ia_status.f.datawords  \ckv_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r12 "kim_ia_capability 2 \kim_ia_capability.r  { \kim_ia_capability.r.part0  } \kim_ia_capability.f  { \kim_ia_capability.f.mem_type  \kim_ia_capability.f.ack_error  \kim_ia_capability.f.sim_tmo  \kim_ia_capability.f.reserved_op  \kim_ia_capability.f.compare  \kim_ia_capability.f.set_init_start  \kim_ia_capability.f.initialize_inc  \kim_ia_capability.f.initialize  \kim_ia_capability.f.reset  \kim_ia_capability.f.disabled  \kim_ia_capability.f.enable  \kim_ia_capability.f.write  \kim_ia_capability.f.read  \kim_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r13 "kim_ia_status 2 \kim_ia_status.r  { \kim_ia_status.r.part0  } \kim_ia_status.f  { \kim_ia_status.f.code  \kim_ia_status.f.datawords  \kim_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r14 "spare 2 \spare.r  { \spare.r.part0  } \spare.f  { \spare.f.spare  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r15 "cceip0_out_ia_wdata 2 \cceip0_out_ia_wdata.r  { \cceip0_out_ia_wdata.r.part2  \cceip0_out_ia_wdata.r.part1  \cceip0_out_ia_wdata.r.part0  } \cceip0_out_ia_wdata.f  { \cceip0_out_ia_wdata.f.tdata_hi  \cceip0_out_ia_wdata.f.tdata_lo  \cceip0_out_ia_wdata.f.eob  \cceip0_out_ia_wdata.f.bytes_vld  \cceip0_out_ia_wdata.f.unused1  \cceip0_out_ia_wdata.f.tid  \cceip0_out_ia_wdata.f.tuser  \cceip0_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r16 "cceip0_out_ia_config 2 \cceip0_out_ia_config.r  { \cceip0_out_ia_config.r.part0  } \cceip0_out_ia_config.f  { \cceip0_out_ia_config.f.op  \cceip0_out_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r17 "cceip0_out_ia_rdata 2 \cceip0_out_ia_rdata.r  { \cceip0_out_ia_rdata.r.part2  \cceip0_out_ia_rdata.r.part1  \cceip0_out_ia_rdata.r.part0  } \cceip0_out_ia_rdata.f  { \cceip0_out_ia_rdata.f.tdata_hi  \cceip0_out_ia_rdata.f.tdata_lo  \cceip0_out_ia_rdata.f.eob  \cceip0_out_ia_rdata.f.bytes_vld  \cceip0_out_ia_rdata.f.unused1  \cceip0_out_ia_rdata.f.tid  \cceip0_out_ia_rdata.f.tuser  \cceip0_out_ia_rdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r18 "cceip0_out_ia_status 2 \cceip0_out_ia_status.r  { \cceip0_out_ia_status.r.part0  } \cceip0_out_ia_status.f  { \cceip0_out_ia_status.f.code  \cceip0_out_ia_status.f.datawords  \cceip0_out_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r19 "cceip0_out_ia_capability 2 \cceip0_out_ia_capability.r  { \cceip0_out_ia_capability.r.part0  } \cceip0_out_ia_capability.f  { \cceip0_out_ia_capability.f.mem_type  \cceip0_out_ia_capability.f.ack_error  \cceip0_out_ia_capability.f.sim_tmo  \cceip0_out_ia_capability.f.reserved_op  \cceip0_out_ia_capability.f.compare  \cceip0_out_ia_capability.f.set_init_start  \cceip0_out_ia_capability.f.initialize_inc  \cceip0_out_ia_capability.f.initialize  \cceip0_out_ia_capability.f.reset  \cceip0_out_ia_capability.f.disabled  \cceip0_out_ia_capability.f.enable  \cceip0_out_ia_capability.f.write  \cceip0_out_ia_capability.f.read  \cceip0_out_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r20 "cceip0_out_im_status 2 \cceip0_out_im_status.r  { \cceip0_out_im_status.r.part0  } \cceip0_out_im_status.f  { \cceip0_out_im_status.f.bank_hi  \cceip0_out_im_status.f.bank_lo  \cceip0_out_im_status.f.overflow  \cceip0_out_im_status.f.wr_pointer  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r21 "cceip0_out_im_config 2 \cceip0_out_im_config.r  { \cceip0_out_im_config.r.part0  } \cceip0_out_im_config.f  { \cceip0_out_im_config.f.mode  \cceip0_out_im_config.f.wr_credit_config  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r22 "cddip0_out_ia_wdata 2 \cddip0_out_ia_wdata.r  { \cddip0_out_ia_wdata.r.part2  \cddip0_out_ia_wdata.r.part1  \cddip0_out_ia_wdata.r.part0  } \cddip0_out_ia_wdata.f  { \cddip0_out_ia_wdata.f.tdata_hi  \cddip0_out_ia_wdata.f.tdata_lo  \cddip0_out_ia_wdata.f.eob  \cddip0_out_ia_wdata.f.bytes_vld  \cddip0_out_ia_wdata.f.unused1  \cddip0_out_ia_wdata.f.tid  \cddip0_out_ia_wdata.f.tuser  \cddip0_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r23 "cddip0_out_ia_config 2 \cddip0_out_ia_config.r  { \cddip0_out_ia_config.r.part0  } \cddip0_out_ia_config.f  { \cddip0_out_ia_config.f.op  \cddip0_out_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r24 "cddip0_out_ia_rdata 2 \cddip0_out_ia_rdata.r  { \cddip0_out_ia_rdata.r.part2  \cddip0_out_ia_rdata.r.part1  \cddip0_out_ia_rdata.r.part0  } \cddip0_out_ia_rdata.f  { \cddip0_out_ia_rdata.f.tdata_hi  \cddip0_out_ia_rdata.f.tdata_lo  \cddip0_out_ia_rdata.f.eob  \cddip0_out_ia_rdata.f.bytes_vld  \cddip0_out_ia_rdata.f.unused1  \cddip0_out_ia_rdata.f.tid  \cddip0_out_ia_rdata.f.tuser  \cddip0_out_ia_rdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r25 "cddip0_out_ia_status 2 \cddip0_out_ia_status.r  { \cddip0_out_ia_status.r.part0  } \cddip0_out_ia_status.f  { \cddip0_out_ia_status.f.code  \cddip0_out_ia_status.f.datawords  \cddip0_out_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r26 "cddip0_out_ia_capability 2 \cddip0_out_ia_capability.r  { \cddip0_out_ia_capability.r.part0  } \cddip0_out_ia_capability.f  { \cddip0_out_ia_capability.f.mem_type  \cddip0_out_ia_capability.f.ack_error  \cddip0_out_ia_capability.f.sim_tmo  \cddip0_out_ia_capability.f.reserved_op  \cddip0_out_ia_capability.f.compare  \cddip0_out_ia_capability.f.set_init_start  \cddip0_out_ia_capability.f.initialize_inc  \cddip0_out_ia_capability.f.initialize  \cddip0_out_ia_capability.f.reset  \cddip0_out_ia_capability.f.disabled  \cddip0_out_ia_capability.f.enable  \cddip0_out_ia_capability.f.write  \cddip0_out_ia_capability.f.read  \cddip0_out_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r27 "cddip0_out_im_status 2 \cddip0_out_im_status.r  { \cddip0_out_im_status.r.part0  } \cddip0_out_im_status.f  { \cddip0_out_im_status.f.bank_hi  \cddip0_out_im_status.f.bank_lo  \cddip0_out_im_status.f.overflow  \cddip0_out_im_status.f.wr_pointer  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r28 "cddip0_out_im_config 2 \cddip0_out_im_config.r  { \cddip0_out_im_config.r.part0  } \cddip0_out_im_config.f  { \cddip0_out_im_config.f.mode  \cddip0_out_im_config.f.wr_credit_config  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r29 "cceip1_out_ia_wdata 2 \cceip1_out_ia_wdata.r  { \cceip1_out_ia_wdata.r.part2  \cceip1_out_ia_wdata.r.part1  \cceip1_out_ia_wdata.r.part0  } \cceip1_out_ia_wdata.f  { \cceip1_out_ia_wdata.f.tdata_hi  \cceip1_out_ia_wdata.f.tdata_lo  \cceip1_out_ia_wdata.f.eob  \cceip1_out_ia_wdata.f.bytes_vld  \cceip1_out_ia_wdata.f.unused1  \cceip1_out_ia_wdata.f.tid  \cceip1_out_ia_wdata.f.tuser  \cceip1_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r30 "cceip1_out_ia_config 2 \cceip1_out_ia_config.r  { \cceip1_out_ia_config.r.part0  } \cceip1_out_ia_config.f  { \cceip1_out_ia_config.f.op  \cceip1_out_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r31 "cceip1_out_ia_rdata 2 \cceip1_out_ia_rdata.r  { \cceip1_out_ia_rdata.r.part2  \cceip1_out_ia_rdata.r.part1  \cceip1_out_ia_rdata.r.part0  } \cceip1_out_ia_rdata.f  { \cceip1_out_ia_rdata.f.tdata_hi  \cceip1_out_ia_rdata.f.tdata_lo  \cceip1_out_ia_rdata.f.eob  \cceip1_out_ia_rdata.f.bytes_vld  \cceip1_out_ia_rdata.f.unused1  \cceip1_out_ia_rdata.f.tid  \cceip1_out_ia_rdata.f.tuser  \cceip1_out_ia_rdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r32 "cceip1_out_ia_status 2 \cceip1_out_ia_status.r  { \cceip1_out_ia_status.r.part0  } \cceip1_out_ia_status.f  { \cceip1_out_ia_status.f.code  \cceip1_out_ia_status.f.datawords  \cceip1_out_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r33 "cceip1_out_ia_capability 2 \cceip1_out_ia_capability.r  { \cceip1_out_ia_capability.r.part0  } \cceip1_out_ia_capability.f  { \cceip1_out_ia_capability.f.mem_type  \cceip1_out_ia_capability.f.ack_error  \cceip1_out_ia_capability.f.sim_tmo  \cceip1_out_ia_capability.f.reserved_op  \cceip1_out_ia_capability.f.compare  \cceip1_out_ia_capability.f.set_init_start  \cceip1_out_ia_capability.f.initialize_inc  \cceip1_out_ia_capability.f.initialize  \cceip1_out_ia_capability.f.reset  \cceip1_out_ia_capability.f.disabled  \cceip1_out_ia_capability.f.enable  \cceip1_out_ia_capability.f.write  \cceip1_out_ia_capability.f.read  \cceip1_out_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r34 "cceip1_out_im_status 2 \cceip1_out_im_status.r  { \cceip1_out_im_status.r.part0  } \cceip1_out_im_status.f  { \cceip1_out_im_status.f.bank_hi  \cceip1_out_im_status.f.bank_lo  \cceip1_out_im_status.f.overflow  \cceip1_out_im_status.f.wr_pointer  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r35 "cceip1_out_im_config 2 \cceip1_out_im_config.r  { \cceip1_out_im_config.r.part0  } \cceip1_out_im_config.f  { \cceip1_out_im_config.f.mode  \cceip1_out_im_config.f.wr_credit_config  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r36 "cddip1_out_ia_wdata 2 \cddip1_out_ia_wdata.r  { \cddip1_out_ia_wdata.r.part2  \cddip1_out_ia_wdata.r.part1  \cddip1_out_ia_wdata.r.part0  } \cddip1_out_ia_wdata.f  { \cddip1_out_ia_wdata.f.tdata_hi  \cddip1_out_ia_wdata.f.tdata_lo  \cddip1_out_ia_wdata.f.eob  \cddip1_out_ia_wdata.f.bytes_vld  \cddip1_out_ia_wdata.f.unused1  \cddip1_out_ia_wdata.f.tid  \cddip1_out_ia_wdata.f.tuser  \cddip1_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r37 "cddip1_out_ia_config 2 \cddip1_out_ia_config.r  { \cddip1_out_ia_config.r.part0  } \cddip1_out_ia_config.f  { \cddip1_out_ia_config.f.op  \cddip1_out_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r38 "cddip1_out_ia_rdata 2 \cddip1_out_ia_rdata.r  { \cddip1_out_ia_rdata.r.part2  \cddip1_out_ia_rdata.r.part1  \cddip1_out_ia_rdata.r.part0  } \cddip1_out_ia_rdata.f  { \cddip1_out_ia_rdata.f.tdata_hi  \cddip1_out_ia_rdata.f.tdata_lo  \cddip1_out_ia_rdata.f.eob  \cddip1_out_ia_rdata.f.bytes_vld  \cddip1_out_ia_rdata.f.unused1  \cddip1_out_ia_rdata.f.tid  \cddip1_out_ia_rdata.f.tuser  \cddip1_out_ia_rdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r39 "cddip1_out_ia_status 2 \cddip1_out_ia_status.r  { \cddip1_out_ia_status.r.part0  } \cddip1_out_ia_status.f  { \cddip1_out_ia_status.f.code  \cddip1_out_ia_status.f.datawords  \cddip1_out_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r40 "cddip1_out_ia_capability 2 \cddip1_out_ia_capability.r  { \cddip1_out_ia_capability.r.part0  } \cddip1_out_ia_capability.f  { \cddip1_out_ia_capability.f.mem_type  \cddip1_out_ia_capability.f.ack_error  \cddip1_out_ia_capability.f.sim_tmo  \cddip1_out_ia_capability.f.reserved_op  \cddip1_out_ia_capability.f.compare  \cddip1_out_ia_capability.f.set_init_start  \cddip1_out_ia_capability.f.initialize_inc  \cddip1_out_ia_capability.f.initialize  \cddip1_out_ia_capability.f.reset  \cddip1_out_ia_capability.f.disabled  \cddip1_out_ia_capability.f.enable  \cddip1_out_ia_capability.f.write  \cddip1_out_ia_capability.f.read  \cddip1_out_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r41 "cddip1_out_im_status 2 \cddip1_out_im_status.r  { \cddip1_out_im_status.r.part0  } \cddip1_out_im_status.f  { \cddip1_out_im_status.f.bank_hi  \cddip1_out_im_status.f.bank_lo  \cddip1_out_im_status.f.overflow  \cddip1_out_im_status.f.wr_pointer  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r42 "cddip1_out_im_config 2 \cddip1_out_im_config.r  { \cddip1_out_im_config.r.part0  } \cddip1_out_im_config.f  { \cddip1_out_im_config.f.mode  \cddip1_out_im_config.f.wr_credit_config  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r43 "cceip2_out_ia_wdata 2 \cceip2_out_ia_wdata.r  { \cceip2_out_ia_wdata.r.part2  \cceip2_out_ia_wdata.r.part1  \cceip2_out_ia_wdata.r.part0  } \cceip2_out_ia_wdata.f  { \cceip2_out_ia_wdata.f.tdata_hi  \cceip2_out_ia_wdata.f.tdata_lo  \cceip2_out_ia_wdata.f.eob  \cceip2_out_ia_wdata.f.bytes_vld  \cceip2_out_ia_wdata.f.unused1  \cceip2_out_ia_wdata.f.tid  \cceip2_out_ia_wdata.f.tuser  \cceip2_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r44 "cceip2_out_ia_config 2 \cceip2_out_ia_config.r  { \cceip2_out_ia_config.r.part0  } \cceip2_out_ia_config.f  { \cceip2_out_ia_config.f.op  \cceip2_out_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r45 "cceip2_out_ia_rdata 2 \cceip2_out_ia_rdata.r  { \cceip2_out_ia_rdata.r.part2  \cceip2_out_ia_rdata.r.part1  \cceip2_out_ia_rdata.r.part0  } \cceip2_out_ia_rdata.f  { \cceip2_out_ia_rdata.f.tdata_hi  \cceip2_out_ia_rdata.f.tdata_lo  \cceip2_out_ia_rdata.f.eob  \cceip2_out_ia_rdata.f.bytes_vld  \cceip2_out_ia_rdata.f.unused1  \cceip2_out_ia_rdata.f.tid  \cceip2_out_ia_rdata.f.tuser  \cceip2_out_ia_rdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r46 "cceip2_out_ia_status 2 \cceip2_out_ia_status.r  { \cceip2_out_ia_status.r.part0  } \cceip2_out_ia_status.f  { \cceip2_out_ia_status.f.code  \cceip2_out_ia_status.f.datawords  \cceip2_out_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r47 "cceip2_out_ia_capability 2 \cceip2_out_ia_capability.r  { \cceip2_out_ia_capability.r.part0  } \cceip2_out_ia_capability.f  { \cceip2_out_ia_capability.f.mem_type  \cceip2_out_ia_capability.f.ack_error  \cceip2_out_ia_capability.f.sim_tmo  \cceip2_out_ia_capability.f.reserved_op  \cceip2_out_ia_capability.f.compare  \cceip2_out_ia_capability.f.set_init_start  \cceip2_out_ia_capability.f.initialize_inc  \cceip2_out_ia_capability.f.initialize  \cceip2_out_ia_capability.f.reset  \cceip2_out_ia_capability.f.disabled  \cceip2_out_ia_capability.f.enable  \cceip2_out_ia_capability.f.write  \cceip2_out_ia_capability.f.read  \cceip2_out_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r48 "cceip2_out_im_status 2 \cceip2_out_im_status.r  { \cceip2_out_im_status.r.part0  } \cceip2_out_im_status.f  { \cceip2_out_im_status.f.bank_hi  \cceip2_out_im_status.f.bank_lo  \cceip2_out_im_status.f.overflow  \cceip2_out_im_status.f.wr_pointer  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r49 "cceip2_out_im_config 2 \cceip2_out_im_config.r  { \cceip2_out_im_config.r.part0  } \cceip2_out_im_config.f  { \cceip2_out_im_config.f.mode  \cceip2_out_im_config.f.wr_credit_config  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r50 "cddip2_out_ia_wdata 2 \cddip2_out_ia_wdata.r  { \cddip2_out_ia_wdata.r.part2  \cddip2_out_ia_wdata.r.part1  \cddip2_out_ia_wdata.r.part0  } \cddip2_out_ia_wdata.f  { \cddip2_out_ia_wdata.f.tdata_hi  \cddip2_out_ia_wdata.f.tdata_lo  \cddip2_out_ia_wdata.f.eob  \cddip2_out_ia_wdata.f.bytes_vld  \cddip2_out_ia_wdata.f.unused1  \cddip2_out_ia_wdata.f.tid  \cddip2_out_ia_wdata.f.tuser  \cddip2_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r51 "cddip2_out_ia_config 2 \cddip2_out_ia_config.r  { \cddip2_out_ia_config.r.part0  } \cddip2_out_ia_config.f  { \cddip2_out_ia_config.f.op  \cddip2_out_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r52 "cddip2_out_ia_rdata 2 \cddip2_out_ia_rdata.r  { \cddip2_out_ia_rdata.r.part2  \cddip2_out_ia_rdata.r.part1  \cddip2_out_ia_rdata.r.part0  } \cddip2_out_ia_rdata.f  { \cddip2_out_ia_rdata.f.tdata_hi  \cddip2_out_ia_rdata.f.tdata_lo  \cddip2_out_ia_rdata.f.eob  \cddip2_out_ia_rdata.f.bytes_vld  \cddip2_out_ia_rdata.f.unused1  \cddip2_out_ia_rdata.f.tid  \cddip2_out_ia_rdata.f.tuser  \cddip2_out_ia_rdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r53 "cddip2_out_ia_status 2 \cddip2_out_ia_status.r  { \cddip2_out_ia_status.r.part0  } \cddip2_out_ia_status.f  { \cddip2_out_ia_status.f.code  \cddip2_out_ia_status.f.datawords  \cddip2_out_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r54 "cddip2_out_ia_capability 2 \cddip2_out_ia_capability.r  { \cddip2_out_ia_capability.r.part0  } \cddip2_out_ia_capability.f  { \cddip2_out_ia_capability.f.mem_type  \cddip2_out_ia_capability.f.ack_error  \cddip2_out_ia_capability.f.sim_tmo  \cddip2_out_ia_capability.f.reserved_op  \cddip2_out_ia_capability.f.compare  \cddip2_out_ia_capability.f.set_init_start  \cddip2_out_ia_capability.f.initialize_inc  \cddip2_out_ia_capability.f.initialize  \cddip2_out_ia_capability.f.reset  \cddip2_out_ia_capability.f.disabled  \cddip2_out_ia_capability.f.enable  \cddip2_out_ia_capability.f.write  \cddip2_out_ia_capability.f.read  \cddip2_out_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r55 "cddip2_out_im_status 2 \cddip2_out_im_status.r  { \cddip2_out_im_status.r.part0  } \cddip2_out_im_status.f  { \cddip2_out_im_status.f.bank_hi  \cddip2_out_im_status.f.bank_lo  \cddip2_out_im_status.f.overflow  \cddip2_out_im_status.f.wr_pointer  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r56 "cddip2_out_im_config 2 \cddip2_out_im_config.r  { \cddip2_out_im_config.r.part0  } \cddip2_out_im_config.f  { \cddip2_out_im_config.f.mode  \cddip2_out_im_config.f.wr_credit_config  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r57 "cceip3_out_ia_wdata 2 \cceip3_out_ia_wdata.r  { \cceip3_out_ia_wdata.r.part2  \cceip3_out_ia_wdata.r.part1  \cceip3_out_ia_wdata.r.part0  } \cceip3_out_ia_wdata.f  { \cceip3_out_ia_wdata.f.tdata_hi  \cceip3_out_ia_wdata.f.tdata_lo  \cceip3_out_ia_wdata.f.eob  \cceip3_out_ia_wdata.f.bytes_vld  \cceip3_out_ia_wdata.f.unused1  \cceip3_out_ia_wdata.f.tid  \cceip3_out_ia_wdata.f.tuser  \cceip3_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r58 "cceip3_out_ia_config 2 \cceip3_out_ia_config.r  { \cceip3_out_ia_config.r.part0  } \cceip3_out_ia_config.f  { \cceip3_out_ia_config.f.op  \cceip3_out_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r59 "cceip3_out_ia_rdata 2 \cceip3_out_ia_rdata.r  { \cceip3_out_ia_rdata.r.part2  \cceip3_out_ia_rdata.r.part1  \cceip3_out_ia_rdata.r.part0  } \cceip3_out_ia_rdata.f  { \cceip3_out_ia_rdata.f.tdata_hi  \cceip3_out_ia_rdata.f.tdata_lo  \cceip3_out_ia_rdata.f.eob  \cceip3_out_ia_rdata.f.bytes_vld  \cceip3_out_ia_rdata.f.unused1  \cceip3_out_ia_rdata.f.tid  \cceip3_out_ia_rdata.f.tuser  \cceip3_out_ia_rdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r60 "cceip3_out_ia_status 2 \cceip3_out_ia_status.r  { \cceip3_out_ia_status.r.part0  } \cceip3_out_ia_status.f  { \cceip3_out_ia_status.f.code  \cceip3_out_ia_status.f.datawords  \cceip3_out_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r61 "cceip3_out_ia_capability 2 \cceip3_out_ia_capability.r  { \cceip3_out_ia_capability.r.part0  } \cceip3_out_ia_capability.f  { \cceip3_out_ia_capability.f.mem_type  \cceip3_out_ia_capability.f.ack_error  \cceip3_out_ia_capability.f.sim_tmo  \cceip3_out_ia_capability.f.reserved_op  \cceip3_out_ia_capability.f.compare  \cceip3_out_ia_capability.f.set_init_start  \cceip3_out_ia_capability.f.initialize_inc  \cceip3_out_ia_capability.f.initialize  \cceip3_out_ia_capability.f.reset  \cceip3_out_ia_capability.f.disabled  \cceip3_out_ia_capability.f.enable  \cceip3_out_ia_capability.f.write  \cceip3_out_ia_capability.f.read  \cceip3_out_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r62 "cceip3_out_im_status 2 \cceip3_out_im_status.r  { \cceip3_out_im_status.r.part0  } \cceip3_out_im_status.f  { \cceip3_out_im_status.f.bank_hi  \cceip3_out_im_status.f.bank_lo  \cceip3_out_im_status.f.overflow  \cceip3_out_im_status.f.wr_pointer  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r63 "cceip3_out_im_config 2 \cceip3_out_im_config.r  { \cceip3_out_im_config.r.part0  } \cceip3_out_im_config.f  { \cceip3_out_im_config.f.mode  \cceip3_out_im_config.f.wr_credit_config  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r64 "cddip3_out_ia_wdata 2 \cddip3_out_ia_wdata.r  { \cddip3_out_ia_wdata.r.part2  \cddip3_out_ia_wdata.r.part1  \cddip3_out_ia_wdata.r.part0  } \cddip3_out_ia_wdata.f  { \cddip3_out_ia_wdata.f.tdata_hi  \cddip3_out_ia_wdata.f.tdata_lo  \cddip3_out_ia_wdata.f.eob  \cddip3_out_ia_wdata.f.bytes_vld  \cddip3_out_ia_wdata.f.unused1  \cddip3_out_ia_wdata.f.tid  \cddip3_out_ia_wdata.f.tuser  \cddip3_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r65 "cddip3_out_ia_config 2 \cddip3_out_ia_config.r  { \cddip3_out_ia_config.r.part0  } \cddip3_out_ia_config.f  { \cddip3_out_ia_config.f.op  \cddip3_out_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r66 "cddip3_out_ia_rdata 2 \cddip3_out_ia_rdata.r  { \cddip3_out_ia_rdata.r.part2  \cddip3_out_ia_rdata.r.part1  \cddip3_out_ia_rdata.r.part0  } \cddip3_out_ia_rdata.f  { \cddip3_out_ia_rdata.f.tdata_hi  \cddip3_out_ia_rdata.f.tdata_lo  \cddip3_out_ia_rdata.f.eob  \cddip3_out_ia_rdata.f.bytes_vld  \cddip3_out_ia_rdata.f.unused1  \cddip3_out_ia_rdata.f.tid  \cddip3_out_ia_rdata.f.tuser  \cddip3_out_ia_rdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r67 "cddip3_out_ia_status 2 \cddip3_out_ia_status.r  { \cddip3_out_ia_status.r.part0  } \cddip3_out_ia_status.f  { \cddip3_out_ia_status.f.code  \cddip3_out_ia_status.f.datawords  \cddip3_out_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r68 "cddip3_out_ia_capability 2 \cddip3_out_ia_capability.r  { \cddip3_out_ia_capability.r.part0  } \cddip3_out_ia_capability.f  { \cddip3_out_ia_capability.f.mem_type  \cddip3_out_ia_capability.f.ack_error  \cddip3_out_ia_capability.f.sim_tmo  \cddip3_out_ia_capability.f.reserved_op  \cddip3_out_ia_capability.f.compare  \cddip3_out_ia_capability.f.set_init_start  \cddip3_out_ia_capability.f.initialize_inc  \cddip3_out_ia_capability.f.initialize  \cddip3_out_ia_capability.f.reset  \cddip3_out_ia_capability.f.disabled  \cddip3_out_ia_capability.f.enable  \cddip3_out_ia_capability.f.write  \cddip3_out_ia_capability.f.read  \cddip3_out_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r69 "cddip3_out_im_status 2 \cddip3_out_im_status.r  { \cddip3_out_im_status.r.part0  } \cddip3_out_im_status.f  { \cddip3_out_im_status.f.bank_hi  \cddip3_out_im_status.f.bank_lo  \cddip3_out_im_status.f.overflow  \cddip3_out_im_status.f.wr_pointer  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r70 "cddip3_out_im_config 2 \cddip3_out_im_config.r  { \cddip3_out_im_config.r.part0  } \cddip3_out_im_config.f  { \cddip3_out_im_config.f.mode  \cddip3_out_im_config.f.wr_credit_config  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r71 "sa_snapshot_ia_wdata 2 \sa_snapshot_ia_wdata.r  { \sa_snapshot_ia_wdata.r.part1  \sa_snapshot_ia_wdata.r.part0  } \sa_snapshot_ia_wdata.f  { \sa_snapshot_ia_wdata.f.unused  \sa_snapshot_ia_wdata.f.upper  \sa_snapshot_ia_wdata.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r72 "sa_snapshot_ia_rdata 2 \sa_snapshot_ia_rdata.r  { \sa_snapshot_ia_rdata.r.part1  \sa_snapshot_ia_rdata.r.part0  } \sa_snapshot_ia_rdata.f  { \sa_snapshot_ia_rdata.f.unused  \sa_snapshot_ia_rdata.f.upper  \sa_snapshot_ia_rdata.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r73 "sa_snapshot_ia_config 2 \sa_snapshot_ia_config.r  { \sa_snapshot_ia_config.r.part0  } \sa_snapshot_ia_config.f  { \sa_snapshot_ia_config.f.op  \sa_snapshot_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r74 "sa_snapshot_ia_status 2 \sa_snapshot_ia_status.r  { \sa_snapshot_ia_status.r.part0  } \sa_snapshot_ia_status.f  { \sa_snapshot_ia_status.f.code  \sa_snapshot_ia_status.f.datawords  \sa_snapshot_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r75 "sa_snapshot_ia_capability 2 \sa_snapshot_ia_capability.r  { \sa_snapshot_ia_capability.r.part0  } \sa_snapshot_ia_capability.f  { \sa_snapshot_ia_capability.f.mem_type  \sa_snapshot_ia_capability.f.ack_error  \sa_snapshot_ia_capability.f.sim_tmo  \sa_snapshot_ia_capability.f.reserved_op  \sa_snapshot_ia_capability.f.compare  \sa_snapshot_ia_capability.f.set_init_start  \sa_snapshot_ia_capability.f.initialize_inc  \sa_snapshot_ia_capability.f.initialize  \sa_snapshot_ia_capability.f.reset  \sa_snapshot_ia_capability.f.disabled  \sa_snapshot_ia_capability.f.enable  \sa_snapshot_ia_capability.f.write  \sa_snapshot_ia_capability.f.read  \sa_snapshot_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r76 "sa_count_ia_wdata 2 \sa_count_ia_wdata.r  { \sa_count_ia_wdata.r.part1  \sa_count_ia_wdata.r.part0  } \sa_count_ia_wdata.f  { \sa_count_ia_wdata.f.unused  \sa_count_ia_wdata.f.upper  \sa_count_ia_wdata.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r77 "sa_count_ia_rdata 2 \sa_count_ia_rdata.r  { \sa_count_ia_rdata.r.part1  \sa_count_ia_rdata.r.part0  } \sa_count_ia_rdata.f  { \sa_count_ia_rdata.f.unused  \sa_count_ia_rdata.f.upper  \sa_count_ia_rdata.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r78 "sa_count_ia_config 2 \sa_count_ia_config.r  { \sa_count_ia_config.r.part0  } \sa_count_ia_config.f  { \sa_count_ia_config.f.op  \sa_count_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r79 "sa_count_ia_status 2 \sa_count_ia_status.r  { \sa_count_ia_status.r.part0  } \sa_count_ia_status.f  { \sa_count_ia_status.f.code  \sa_count_ia_status.f.datawords  \sa_count_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r80 "sa_count_ia_capability 2 \sa_count_ia_capability.r  { \sa_count_ia_capability.r.part0  } \sa_count_ia_capability.f  { \sa_count_ia_capability.f.mem_type  \sa_count_ia_capability.f.ack_error  \sa_count_ia_capability.f.sim_tmo  \sa_count_ia_capability.f.reserved_op  \sa_count_ia_capability.f.compare  \sa_count_ia_capability.f.set_init_start  \sa_count_ia_capability.f.initialize_inc  \sa_count_ia_capability.f.initialize  \sa_count_ia_capability.f.reset  \sa_count_ia_capability.f.disabled  \sa_count_ia_capability.f.enable  \sa_count_ia_capability.f.write  \sa_count_ia_capability.f.read  \sa_count_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r81 "sa_ctrl_ia_wdata 2 \sa_ctrl_ia_wdata.r  { \sa_ctrl_ia_wdata.r.part0  } \sa_ctrl_ia_wdata.f  { \sa_ctrl_ia_wdata.f.spare  \sa_ctrl_ia_wdata.f.sa_event_sel  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r82 "sa_ctrl_ia_rdata 2 \sa_ctrl_ia_rdata.r  { \sa_ctrl_ia_rdata.r.part0  } \sa_ctrl_ia_rdata.f  { \sa_ctrl_ia_rdata.f.spare  \sa_ctrl_ia_rdata.f.sa_event_sel  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r83 "sa_ctrl_ia_config 2 \sa_ctrl_ia_config.r  { \sa_ctrl_ia_config.r.part0  } \sa_ctrl_ia_config.f  { \sa_ctrl_ia_config.f.op  \sa_ctrl_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r84 "sa_ctrl_ia_status 2 \sa_ctrl_ia_status.r  { \sa_ctrl_ia_status.r.part0  } \sa_ctrl_ia_status.f  { \sa_ctrl_ia_status.f.code  \sa_ctrl_ia_status.f.datawords  \sa_ctrl_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r85 "sa_ctrl_ia_capability 2 \sa_ctrl_ia_capability.r  { \sa_ctrl_ia_capability.r.part0  } \sa_ctrl_ia_capability.f  { \sa_ctrl_ia_capability.f.mem_type  \sa_ctrl_ia_capability.f.ack_error  \sa_ctrl_ia_capability.f.sim_tmo  \sa_ctrl_ia_capability.f.reserved_op  \sa_ctrl_ia_capability.f.compare  \sa_ctrl_ia_capability.f.set_init_start  \sa_ctrl_ia_capability.f.initialize_inc  \sa_ctrl_ia_capability.f.initialize  \sa_ctrl_ia_capability.f.reset  \sa_ctrl_ia_capability.f.disabled  \sa_ctrl_ia_capability.f.enable  \sa_ctrl_ia_capability.f.write  \sa_ctrl_ia_capability.f.read  \sa_ctrl_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r86 "sa_ctrl_rst_dat%s 2 \sa_ctrl_rst_dat%s.r  { \sa_ctrl_rst_dat%s.r.part0  } \sa_ctrl_rst_dat%s.f  { \sa_ctrl_rst_dat%s.f.spare  \sa_ctrl_rst_dat%s.f.sa_event_sel  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r37 "cceip0_im_din 2 \cceip0_im_din.data  { \cceip0_im_din.data.data  } \cceip0_im_din.desc  { \cceip0_im_din.desc.eob  \cceip0_im_din.desc.bytes_vld  \cceip0_im_din.desc.im_meta  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r38 "cddip0_im_din 2 \cddip0_im_din.data  { \cddip0_im_din.data.data  } \cddip0_im_din.desc  { \cddip0_im_din.desc.eob  \cddip0_im_din.desc.bytes_vld  \cddip0_im_din.desc.im_meta  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r39 "cceip1_im_din 2 \cceip1_im_din.data  { \cceip1_im_din.data.data  } \cceip1_im_din.desc  { \cceip1_im_din.desc.eob  \cceip1_im_din.desc.bytes_vld  \cceip1_im_din.desc.im_meta  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r40 "cddip1_im_din 2 \cddip1_im_din.data  { \cddip1_im_din.data.data  } \cddip1_im_din.desc  { \cddip1_im_din.desc.eob  \cddip1_im_din.desc.bytes_vld  \cddip1_im_din.desc.im_meta  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r41 "cceip2_im_din 2 \cceip2_im_din.data  { \cceip2_im_din.data.data  } \cceip2_im_din.desc  { \cceip2_im_din.desc.eob  \cceip2_im_din.desc.bytes_vld  \cceip2_im_din.desc.im_meta  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r42 "cddip2_im_din 2 \cddip2_im_din.data  { \cddip2_im_din.data.data  } \cddip2_im_din.desc  { \cddip2_im_din.desc.eob  \cddip2_im_din.desc.bytes_vld  \cddip2_im_din.desc.im_meta  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r43 "cceip3_im_din 2 \cceip3_im_din.data  { \cceip3_im_din.data.data  } \cceip3_im_din.desc  { \cceip3_im_din.desc.eob  \cceip3_im_din.desc.bytes_vld  \cceip3_im_din.desc.im_meta  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r44 "cddip3_im_din 2 \cddip3_im_din.data  { \cddip3_im_din.data.data  } \cddip3_im_din.desc  { \cddip3_im_din.desc.eob  \cddip3_im_din.desc.bytes_vld  \cddip3_im_din.desc.im_meta  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r45 "im_consumed_kme_cceip0 2 \im_consumed_kme_cceip0.bank_hi  \im_consumed_kme_cceip0.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r46 "im_available_kme_cceip0 2 \im_available_kme_cceip0.bank_hi  \im_available_kme_cceip0.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r47 "im_consumed_kme_cddip0 2 \im_consumed_kme_cddip0.bank_hi  \im_consumed_kme_cddip0.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r48 "im_available_kme_cddip0 2 \im_available_kme_cddip0.bank_hi  \im_available_kme_cddip0.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r49 "im_consumed_kme_cceip1 2 \im_consumed_kme_cceip1.bank_hi  \im_consumed_kme_cceip1.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r50 "im_available_kme_cceip1 2 \im_available_kme_cceip1.bank_hi  \im_available_kme_cceip1.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r51 "im_consumed_kme_cddip1 2 \im_consumed_kme_cddip1.bank_hi  \im_consumed_kme_cddip1.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r52 "im_available_kme_cddip1 2 \im_available_kme_cddip1.bank_hi  \im_available_kme_cddip1.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r53 "im_consumed_kme_cceip2 2 \im_consumed_kme_cceip2.bank_hi  \im_consumed_kme_cceip2.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r54 "im_available_kme_cceip2 2 \im_available_kme_cceip2.bank_hi  \im_available_kme_cceip2.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r55 "im_consumed_kme_cddip2 2 \im_consumed_kme_cddip2.bank_hi  \im_consumed_kme_cddip2.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r56 "im_available_kme_cddip2 2 \im_available_kme_cddip2.bank_hi  \im_available_kme_cddip2.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r57 "im_consumed_kme_cceip3 2 \im_consumed_kme_cceip3.bank_hi  \im_consumed_kme_cceip3.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r58 "im_available_kme_cceip3 2 \im_available_kme_cceip3.bank_hi  \im_available_kme_cceip3.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r59 "im_consumed_kme_cddip3 2 \im_consumed_kme_cddip3.bank_hi  \im_consumed_kme_cddip3.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r60 "im_available_kme_cddip3 2 \im_available_kme_cddip3.bank_hi  \im_available_kme_cddip3.bank_lo "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r61 "kme_cceip0_ob_out_post 6 \kme_cceip0_ob_out_post.tvalid  \kme_cceip0_ob_out_post.tlast  \kme_cceip0_ob_out_post.tid  \kme_cceip0_ob_out_post.tstrb  \kme_cceip0_ob_out_post.tuser  \kme_cceip0_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r62 "kme_cceip1_ob_out_post 6 \kme_cceip1_ob_out_post.tvalid  \kme_cceip1_ob_out_post.tlast  \kme_cceip1_ob_out_post.tid  \kme_cceip1_ob_out_post.tstrb  \kme_cceip1_ob_out_post.tuser  \kme_cceip1_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r63 "kme_cceip2_ob_out_post 6 \kme_cceip2_ob_out_post.tvalid  \kme_cceip2_ob_out_post.tlast  \kme_cceip2_ob_out_post.tid  \kme_cceip2_ob_out_post.tstrb  \kme_cceip2_ob_out_post.tuser  \kme_cceip2_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r64 "kme_cceip3_ob_out_post 6 \kme_cceip3_ob_out_post.tvalid  \kme_cceip3_ob_out_post.tlast  \kme_cceip3_ob_out_post.tid  \kme_cceip3_ob_out_post.tstrb  \kme_cceip3_ob_out_post.tuser  \kme_cceip3_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r65 "kme_cddip0_ob_out_post 6 \kme_cddip0_ob_out_post.tvalid  \kme_cddip0_ob_out_post.tlast  \kme_cddip0_ob_out_post.tid  \kme_cddip0_ob_out_post.tstrb  \kme_cddip0_ob_out_post.tuser  \kme_cddip0_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r66 "kme_cddip1_ob_out_post 6 \kme_cddip1_ob_out_post.tvalid  \kme_cddip1_ob_out_post.tlast  \kme_cddip1_ob_out_post.tid  \kme_cddip1_ob_out_post.tstrb  \kme_cddip1_ob_out_post.tuser  \kme_cddip1_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r67 "kme_cddip2_ob_out_post 6 \kme_cddip2_ob_out_post.tvalid  \kme_cddip2_ob_out_post.tlast  \kme_cddip2_ob_out_post.tid  \kme_cddip2_ob_out_post.tstrb  \kme_cddip2_ob_out_post.tuser  \kme_cddip2_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r68 "kme_cddip3_ob_out_post 6 \kme_cddip3_ob_out_post.tvalid  \kme_cddip3_ob_out_post.tlast  \kme_cddip3_ob_out_post.tid  \kme_cddip3_ob_out_post.tstrb  \kme_cddip3_ob_out_post.tuser  \kme_cddip3_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r87 "revid_wire 2 \revid_wire.r  { \revid_wire.r.part0  } \revid_wire.f  { \revid_wire.f.revid  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "68"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_NUM "87"
endmodule
