library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity bimc_master is
  generic (
    MSB : integer := 71;
    BIMC_FLENGTH : integer := 72;
    NOP : std_logic_vector := std_logic_vector'("00000000");
    RD_REG : std_logic_vector := std_logic_vector'("00000001");
    WR_ID : std_logic_vector := std_logic_vector'("00000010");
    POLL_ERR : std_logic_vector := std_logic_vector'("00000011");
    WR_ECTRL : std_logic_vector := std_logic_vector'("00001010");
    WR_ECCP : std_logic_vector := std_logic_vector'("00001011");
    WR_ECCCNT : std_logic_vector := std_logic_vector'("00001100");
    WR_ECCIN : std_logic_vector := std_logic_vector'("00010000");
    WR_ECCOUT : std_logic_vector := std_logic_vector'("00010001");
    WR_TM : std_logic_vector := std_logic_vector'("00011110");
    WR_LVM : std_logic_vector := std_logic_vector'("00011111");
    WR_MLVM : std_logic_vector := std_logic_vector'("00100000");
    WR_MRDTEN : std_logic_vector := std_logic_vector'("00100001");
    WR_RDT : std_logic_vector := std_logic_vector'("00100010");
    WR_WBT : std_logic_vector := std_logic_vector'("00100011");
    WR_WMS : std_logic_vector := std_logic_vector'("00100100");
    MEM_INIT : std_logic_vector := std_logic_vector'("11111111");
    RESET : std_logic_vector := std_logic_vector'("0000");
    AUTOID : std_logic_vector := std_logic_vector'("1011");
    CPU : std_logic_vector := std_logic_vector'("0001");
    IDLE : std_logic_vector := std_logic_vector'("0010");
    AUTOPOLL : std_logic_vector := std_logic_vector'("0111");
    MEMWRINIT : std_logic_vector := std_logic_vector'("1000");
    PICK_NXT : std_logic_vector := std_logic_vector'("0011");
    ECCPAR_DEBUG : std_logic_vector := std_logic_vector'("0101");
    COMMAND : std_logic_vector := std_logic_vector'("0001");
    CMD_DONE : std_logic_vector := std_logic_vector'("0000");
    RESPONSE_CMD : std_logic_vector := std_logic_vector'("0011");
    RESPONSE_IDLE : std_logic_vector := std_logic_vector'("0100");
    RESPONSE_MEM : std_logic_vector := std_logic_vector'("0101");
    RSP_DONE : std_logic_vector := std_logic_vector'("0110");
    POLL_ERR_CMD : std_logic_vector := std_logic_vector'("0111");
    POLL_ERR_IDLE : std_logic_vector := std_logic_vector'("1000");
    POLL_ERR_MEM : std_logic_vector := std_logic_vector'("1001");
    POLL_ERR_DONE : std_logic_vector := std_logic_vector'("1010")
  ) ;
  port (
    bimc_ecc_error : out std_logic ;
    bimc_interrupt : out std_logic ;
    bimc_odat : out std_logic ;
    bimc_osync : out std_logic ;
    bimc_rst_n : out std_logic ;
    clk : in std_logic ;
    rst_n : in std_logic ;
    bimc_idat : in std_logic ;
    bimc_isync : in std_logic ;
    o_bimc_monitor_mask : in std_logic_vector(6 downto 0) ;
    o_bimc_ecc_uncorrectable_error_cnt : in std_logic_vector(31 downto 0) ;
    o_bimc_ecc_correctable_error_cnt : in std_logic_vector(31 downto 0) ;
    o_bimc_parity_error_cnt : in std_logic_vector(31 downto 0) ;
    o_bimc_global_config : in std_logic_vector(31 downto 0) ;
    o_bimc_eccpar_debug : in std_logic_vector(28 downto 0) ;
    o_bimc_cmd2 : in std_logic_vector(10 downto 0) ;
    o_bimc_cmd1 : in std_logic_vector(31 downto 0) ;
    o_bimc_cmd0 : in std_logic_vector(31 downto 0) ;
    o_bimc_rxcmd2 : in std_logic_vector(9 downto 0) ;
    o_bimc_rxrsp2 : in std_logic_vector(9 downto 0) ;
    o_bimc_pollrsp2 : in std_logic_vector(9 downto 0) ;
    o_bimc_dbgcmd2 : in std_logic_vector(9 downto 0) ;
    i_bimc_monitor : out std_logic_vector(6 downto 0) ;
    i_bimc_ecc_uncorrectable_error_cnt : out std_logic_vector(31 downto 0) ;
    i_bimc_ecc_correctable_error_cnt : out std_logic_vector(31 downto 0) ;
    i_bimc_parity_error_cnt : out std_logic_vector(31 downto 0) ;
    i_bimc_global_config : out std_logic_vector(31 downto 0) ;
    i_bimc_memid : out std_logic_vector(11 downto 0) ;
    i_bimc_eccpar_debug : out std_logic_vector(28 downto 0) ;
    i_bimc_cmd2 : out std_logic_vector(10 downto 0) ;
    i_bimc_rxcmd2 : out std_logic_vector(9 downto 0) ;
    i_bimc_rxcmd1 : out std_logic_vector(31 downto 0) ;
    i_bimc_rxcmd0 : out std_logic_vector(31 downto 0) ;
    i_bimc_rxrsp2 : out std_logic_vector(9 downto 0) ;
    i_bimc_rxrsp1 : out std_logic_vector(31 downto 0) ;
    i_bimc_rxrsp0 : out std_logic_vector(31 downto 0) ;
    i_bimc_pollrsp2 : out std_logic_vector(9 downto 0) ;
    i_bimc_pollrsp1 : out std_logic_vector(31 downto 0) ;
    i_bimc_pollrsp0 : out std_logic_vector(31 downto 0) ;
    i_bimc_dbgcmd2 : out std_logic_vector(9 downto 0) ;
    i_bimc_dbgcmd1 : out std_logic_vector(31 downto 0) ;
  i_bimc_dbgcmd0 : out std_logic_vector(31 downto 0) ) ;
  attribute _2_state_: integer;
  attribute celldefine : integer;
  attribute celldefine of bimc_master: entity is 1 ;
end bimc_master ;
