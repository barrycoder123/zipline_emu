
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme ( kme_interrupt, kme_ib_tready, kme_cceip0_ob_tvalid, 
	kme_cceip0_ob_tlast, kme_cceip0_ob_tid, kme_cceip0_ob_tstrb, 
	kme_cceip0_ob_tuser, kme_cceip0_ob_tdata, apb_prdata, apb_pready, 
	apb_pslverr, kme_idle, clk, rst_n, scan_en, scan_mode, scan_rst_n, 
	ovstb, lvm, mlvm, disable_debug_cmd, disable_unencrypted_keys, 
	kme_ib_tvalid, kme_ib_tlast, kme_ib_tid, kme_ib_tstrb, kme_ib_tuser, 
	kme_ib_tdata, kme_cceip0_ob_tready, apb_paddr, apb_psel, apb_penable, 
	apb_pwrite, apb_pwdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output kme_interrupt;
output kme_ib_tready;
output kme_cceip0_ob_tvalid;
output kme_cceip0_ob_tlast;
output [0:0] kme_cceip0_ob_tid;
output [7:0] kme_cceip0_ob_tstrb;
output [7:0] kme_cceip0_ob_tuser;
output [63:0] kme_cceip0_ob_tdata;
output [31:0] apb_prdata;
output apb_pready;
output apb_pslverr;
output kme_idle;
input clk;
input rst_n;
input scan_en;
input scan_mode;
input scan_rst_n;
input ovstb;
input lvm;
input mlvm;
input disable_debug_cmd;
input disable_unencrypted_keys;
input kme_ib_tvalid;
input kme_ib_tlast;
input [0:0] kme_ib_tid;
input [7:0] kme_ib_tstrb;
input [7:0] kme_ib_tuser;
input [63:0] kme_ib_tdata;
input kme_cceip0_ob_tready;
input [15:0] apb_paddr;
input apb_psel;
input apb_penable;
input apb_pwrite;
input [31:0] apb_pwdata;
wire debug_kme_ib_tready;
wire always_validate_kim_ref;
wire axi_bimc_idat;
wire axi_bimc_isync;
wire axi_bimc_odat;
wire axi_bimc_osync;
wire axi_mbe;
wire bimc_rst_n;
wire cceip_encrypt_bimc_idat;
wire cceip_encrypt_bimc_isync;
wire cceip_encrypt_bimc_odat;
wire cceip_encrypt_bimc_osync;
wire cceip_encrypt_mbe;
wire cceip_validate_bimc_idat;
wire cceip_validate_bimc_isync;
wire cceip_validate_bimc_odat;
wire cceip_validate_bimc_osync;
wire cceip_validate_mbe;
wire cddip_decrypt_bimc_idat;
wire cddip_decrypt_bimc_isync;
wire cddip_decrypt_bimc_odat;
wire cddip_decrypt_bimc_osync;
wire cddip_decrypt_mbe;
wire [14:0] ckv_addr;
wire [63:0] ckv_dout;
wire ckv_mbe;
wire ckv_rd;
wire [63:0] debug_kme_ib_tdata;
wire [0:0] debug_kme_ib_tid;
wire debug_kme_ib_tlast;
wire [7:0] debug_kme_ib_tstrb;
wire [7:0] debug_kme_ib_tuser;
wire debug_kme_ib_tvalid;
wire [31:0] kdf_test_key_size;
wire kdf_test_mode_en;
wire [13:0] kim_addr;
wire kim_mbe;
wire kim_rd;
wire manual_txc;
wire rst_sync_n;
wire [255:0] seed0_internal_state_key;
wire [127:0] seed0_internal_state_value;
wire seed0_invalidate;
wire [47:0] seed0_reseed_interval;
wire seed0_valid;
wire [255:0] seed1_internal_state_key;
wire [127:0] seed1_internal_state_value;
wire seed1_invalidate;
wire [47:0] seed1_reseed_interval;
wire seed1_valid;
wire set_gcm_tag_fail_int;
wire set_key_tlv_miscmp_int;
wire [7:0] set_rsm_is_backpressuring;
wire set_tlv_bip2_error_int;
wire set_txc_bp_int;
wire suppress_key_tlvs;
wire clock;
wire clock_1;
wire kme_cceip1_ob_tready;
wire kme_cceip2_ob_tready;
wire kme_cceip3_ob_tready;
wire kme_cddip0_ob_tready;
wire kme_cddip1_ob_tready;
wire kme_cddip2_ob_tready;
wire kme_cddip3_ob_tready;
wire _zy_simnet_kme_ib_out_0_w$;
wire [0:82] _zy_simnet_kme_cceip0_ob_out_pre_1_w$;
wire [0:82] _zy_simnet_kme_cceip1_ob_out_pre_2_w$;
wire [0:82] _zy_simnet_kme_cceip2_ob_out_pre_3_w$;
wire [0:82] _zy_simnet_kme_cceip3_ob_out_pre_4_w$;
wire [0:82] _zy_simnet_kme_cddip0_ob_out_pre_5_w$;
wire [0:82] _zy_simnet_kme_cddip1_ob_out_pre_6_w$;
wire [0:82] _zy_simnet_kme_cddip2_ob_out_pre_7_w$;
wire [0:82] _zy_simnet_kme_cddip3_ob_out_pre_8_w$;
wire [0:31] _zy_simnet_idle_components_9_w$;
wire [0:82] _zy_simnet_kme_ib_in_10_w$;
wire _zy_simnet_kme_cceip0_ob_in_mod_11_w$;
wire _zy_simnet_kme_cceip1_ob_in_mod_12_w$;
wire _zy_simnet_kme_cceip2_ob_in_mod_13_w$;
wire _zy_simnet_kme_cceip3_ob_in_mod_14_w$;
wire _zy_simnet_kme_cddip0_ob_in_mod_15_w$;
wire _zy_simnet_kme_cddip1_ob_in_mod_16_w$;
wire _zy_simnet_kme_cddip2_ob_in_mod_17_w$;
wire _zy_simnet_kme_cddip3_ob_in_mod_18_w$;
wire [0:37] _zy_simnet_kim_dout_19_w$;
wire [0:8] _zy_simnet_tready_override_21_w$;
wire [0:6] _zy_simnet_cceip_encrypt_kop_fifo_override_22_w$;
wire [0:6] _zy_simnet_cceip_validate_kop_fifo_override_23_w$;
wire [0:6] _zy_simnet_cddip_decrypt_kop_fifo_override_24_w$;
wire [0:31] _zy_simnet_sa_global_ctrl_25_w$;
wire [0:15] _zy_simnet_rbus_ring_i_26_w$;
wire _zy_simnet_rbus_ring_i_27_w$;
wire [0:31] _zy_simnet_rbus_ring_i_28_w$;
wire _zy_simnet_rbus_ring_i_29_w$;
wire [0:31] _zy_simnet_rbus_ring_o_30_w$;
wire _zy_simnet_rbus_ring_o_31_w$;
wire _zy_simnet_rbus_ring_o_32_w$;
wire _zy_simnet_rbus_ring_o_33_w$;
wire _zy_simnet_rbus_ring_o_34_w$;
wire [0:83] _zy_simnet_rbus_ring_o_35_w$;
wire [0:82] _zy_simnet_kme_cceip0_ob_out_36_w$;
wire _zy_simnet_kme_cceip0_ob_in_mod_37_w$;
wire [0:82] _zy_simnet_kme_cceip1_ob_out_38_w$;
wire _zy_simnet_kme_cceip1_ob_in_mod_39_w$;
wire [0:82] _zy_simnet_kme_cceip2_ob_out_40_w$;
wire _zy_simnet_kme_cceip2_ob_in_mod_41_w$;
wire [0:82] _zy_simnet_kme_cceip3_ob_out_42_w$;
wire _zy_simnet_kme_cceip3_ob_in_mod_43_w$;
wire [0:82] _zy_simnet_kme_cddip0_ob_out_44_w$;
wire _zy_simnet_kme_cddip0_ob_in_mod_45_w$;
wire [0:82] _zy_simnet_kme_cddip1_ob_out_46_w$;
wire _zy_simnet_kme_cddip1_ob_in_mod_47_w$;
wire [0:82] _zy_simnet_kme_cddip2_ob_out_48_w$;
wire _zy_simnet_kme_cddip2_ob_in_mod_49_w$;
wire [0:82] _zy_simnet_kme_cddip3_ob_out_50_w$;
wire _zy_simnet_kme_cddip3_ob_in_mod_51_w$;
wire [0:37] _zy_simnet_kim_dout_52_w$;
wire [0:8] _zy_simnet_tready_override_54_w$;
wire [0:6] _zy_simnet_cceip_encrypt_kop_fifo_override_55_w$;
wire [0:6] _zy_simnet_cceip_validate_kop_fifo_override_56_w$;
wire [0:6] _zy_simnet_cddip_decrypt_kop_fifo_override_57_w$;
wire [0:31] _zy_simnet_sa_global_ctrl_58_w$;
wire [0:83] _zy_simnet_rbus_ring_i_59_w$;
wire [0:15] _zy_simnet_cio_60;
wire [0:15] _zy_simnet_cio_61;
wire [0:82] _zy_simnet_kme_cceip0_ob_out_pre_62_w$;
wire _zy_simnet_kme_cceip0_ob_in_63_w$;
wire [0:82] _zy_simnet_kme_cceip1_ob_out_pre_64_w$;
wire _zy_simnet_kme_cceip1_ob_in_65_w$;
wire [0:82] _zy_simnet_kme_cceip2_ob_out_pre_66_w$;
wire _zy_simnet_kme_cceip2_ob_in_67_w$;
wire [0:82] _zy_simnet_kme_cceip3_ob_out_pre_68_w$;
wire _zy_simnet_kme_cceip3_ob_in_69_w$;
wire [0:82] _zy_simnet_kme_cddip0_ob_out_pre_70_w$;
wire _zy_simnet_kme_cddip0_ob_in_71_w$;
wire [0:82] _zy_simnet_kme_cddip1_ob_out_pre_72_w$;
wire _zy_simnet_kme_cddip1_ob_in_73_w$;
wire [0:82] _zy_simnet_kme_cddip2_ob_out_pre_74_w$;
wire _zy_simnet_kme_cddip2_ob_in_75_w$;
wire [0:82] _zy_simnet_kme_cddip3_ob_out_pre_76_w$;
wire _zy_simnet_kme_cddip3_ob_in_77_w$;
wire [0:31] _zy_simnet_idle_components_78_w$;
wire _zyclock_1_x$tbc;
wire [83:0] rbus_ring_i;
wire [83:0] rbus_ring_o;
wire [82:0] kme_ib_in;
wire [0:0] kme_ib_out;
wire [82:0] kme_cceip0_ob_out;
wire [82:0] kme_cceip1_ob_out;
wire [82:0] kme_cceip2_ob_out;
wire [82:0] kme_cceip3_ob_out;
wire [0:0] kme_cceip0_ob_in;
wire [0:0] kme_cceip1_ob_in;
wire [0:0] kme_cceip2_ob_in;
wire [0:0] kme_cceip3_ob_in;
wire [82:0] kme_cddip0_ob_out;
wire [82:0] kme_cddip1_ob_out;
wire [82:0] kme_cddip2_ob_out;
wire [82:0] kme_cddip3_ob_out;
wire [0:0] kme_cddip0_ob_in;
wire [0:0] kme_cddip1_ob_in;
wire [0:0] kme_cddip2_ob_in;
wire [0:0] kme_cddip3_ob_in;
wire [6:0] cceip_encrypt_kop_fifo_override;
wire [6:0] cceip_validate_kop_fifo_override;
wire [6:0] cddip_decrypt_kop_fifo_override;
wire [31:0] idle_components;
wire [37:0] kim_dout;
wire [0:0] kme_cceip0_ob_in_mod;
wire [82:0] kme_cceip0_ob_out_pre;
wire [0:0] kme_cceip1_ob_in_mod;
wire [82:0] kme_cceip1_ob_out_pre;
wire [0:0] kme_cceip2_ob_in_mod;
wire [82:0] kme_cceip2_ob_out_pre;
wire [0:0] kme_cceip3_ob_in_mod;
wire [82:0] kme_cceip3_ob_out_pre;
wire [0:0] kme_cddip0_ob_in_mod;
wire [82:0] kme_cddip0_ob_out_pre;
wire [0:0] kme_cddip1_ob_in_mod;
wire [82:0] kme_cddip1_ob_out_pre;
wire [0:0] kme_cddip2_ob_in_mod;
wire [82:0] kme_cddip2_ob_out_pre;
wire [0:0] kme_cddip3_ob_in_mod;
wire [82:0] kme_cddip3_ob_out_pre;
wire [31:0] sa_global_ctrl;
wire [8:0] tready_override;
supply0 n1;
supply1 n2;
wire [15:0] \rbus_ring_i.addr ;
wire \rbus_ring_i.wr_strb ;
wire [31:0] \rbus_ring_i.wr_data ;
wire \rbus_ring_i.rd_strb ;
wire [31:0] \rbus_ring_i.rd_data ;
wire \rbus_ring_i.ack ;
wire \rbus_ring_i.err_ack ;
wire [15:0] \rbus_ring_o.addr ;
wire \rbus_ring_o.wr_strb ;
wire [31:0] \rbus_ring_o.wr_data ;
wire \rbus_ring_o.rd_strb ;
wire [31:0] \rbus_ring_o.rd_data ;
wire \rbus_ring_o.ack ;
wire \rbus_ring_o.err_ack ;
wire \kme_ib_in.tvalid ;
wire \kme_ib_in.tlast ;
wire [0:0] \kme_ib_in.tid ;
wire [7:0] \kme_ib_in.tstrb ;
wire [7:0] \kme_ib_in.tuser ;
wire [63:0] \kme_ib_in.tdata ;
wire \kme_ib_out.tready ;
wire \kme_cceip0_ob_out.tvalid ;
wire \kme_cceip0_ob_out.tlast ;
wire [0:0] \kme_cceip0_ob_out.tid ;
wire [7:0] \kme_cceip0_ob_out.tstrb ;
wire [7:0] \kme_cceip0_ob_out.tuser ;
wire [63:0] \kme_cceip0_ob_out.tdata ;
wire \kme_cceip1_ob_out.tvalid ;
wire \kme_cceip1_ob_out.tlast ;
wire [0:0] \kme_cceip1_ob_out.tid ;
wire [7:0] \kme_cceip1_ob_out.tstrb ;
wire [7:0] \kme_cceip1_ob_out.tuser ;
wire [63:0] \kme_cceip1_ob_out.tdata ;
wire \kme_cceip2_ob_out.tvalid ;
wire \kme_cceip2_ob_out.tlast ;
wire [0:0] \kme_cceip2_ob_out.tid ;
wire [7:0] \kme_cceip2_ob_out.tstrb ;
wire [7:0] \kme_cceip2_ob_out.tuser ;
wire [63:0] \kme_cceip2_ob_out.tdata ;
wire \kme_cceip3_ob_out.tvalid ;
wire \kme_cceip3_ob_out.tlast ;
wire [0:0] \kme_cceip3_ob_out.tid ;
wire [7:0] \kme_cceip3_ob_out.tstrb ;
wire [7:0] \kme_cceip3_ob_out.tuser ;
wire [63:0] \kme_cceip3_ob_out.tdata ;
wire \kme_cceip0_ob_in.tready ;
wire \kme_cceip1_ob_in.tready ;
wire \kme_cceip2_ob_in.tready ;
wire \kme_cceip3_ob_in.tready ;
wire \kme_cddip0_ob_out.tvalid ;
wire \kme_cddip0_ob_out.tlast ;
wire [0:0] \kme_cddip0_ob_out.tid ;
wire [7:0] \kme_cddip0_ob_out.tstrb ;
wire [7:0] \kme_cddip0_ob_out.tuser ;
wire [63:0] \kme_cddip0_ob_out.tdata ;
wire \kme_cddip1_ob_out.tvalid ;
wire \kme_cddip1_ob_out.tlast ;
wire [0:0] \kme_cddip1_ob_out.tid ;
wire [7:0] \kme_cddip1_ob_out.tstrb ;
wire [7:0] \kme_cddip1_ob_out.tuser ;
wire [63:0] \kme_cddip1_ob_out.tdata ;
wire \kme_cddip2_ob_out.tvalid ;
wire \kme_cddip2_ob_out.tlast ;
wire [0:0] \kme_cddip2_ob_out.tid ;
wire [7:0] \kme_cddip2_ob_out.tstrb ;
wire [7:0] \kme_cddip2_ob_out.tuser ;
wire [63:0] \kme_cddip2_ob_out.tdata ;
wire \kme_cddip3_ob_out.tvalid ;
wire \kme_cddip3_ob_out.tlast ;
wire [0:0] \kme_cddip3_ob_out.tid ;
wire [7:0] \kme_cddip3_ob_out.tstrb ;
wire [7:0] \kme_cddip3_ob_out.tuser ;
wire [63:0] \kme_cddip3_ob_out.tdata ;
wire \kme_cddip0_ob_in.tready ;
wire \kme_cddip1_ob_in.tready ;
wire \kme_cddip2_ob_in.tready ;
wire \kme_cddip3_ob_in.tready ;
wire [6:0] \cceip_encrypt_kop_fifo_override.r.part0 ;
wire \cceip_encrypt_kop_fifo_override.f.gcm_status_data_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.tlv_sb_data_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.kdf_cmd_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.kdfstream_cmd_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.keyfilter_cmd_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.gcm_tag_data_fifo ;
wire \cceip_encrypt_kop_fifo_override.f.gcm_cmd_fifo ;
wire [6:0] \cceip_validate_kop_fifo_override.r.part0 ;
wire \cceip_validate_kop_fifo_override.f.gcm_status_data_fifo ;
wire \cceip_validate_kop_fifo_override.f.tlv_sb_data_fifo ;
wire \cceip_validate_kop_fifo_override.f.kdf_cmd_fifo ;
wire \cceip_validate_kop_fifo_override.f.kdfstream_cmd_fifo ;
wire \cceip_validate_kop_fifo_override.f.keyfilter_cmd_fifo ;
wire \cceip_validate_kop_fifo_override.f.gcm_tag_data_fifo ;
wire \cceip_validate_kop_fifo_override.f.gcm_cmd_fifo ;
wire [6:0] \cddip_decrypt_kop_fifo_override.r.part0 ;
wire \cddip_decrypt_kop_fifo_override.f.gcm_status_data_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.tlv_sb_data_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.kdf_cmd_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.kdfstream_cmd_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.keyfilter_cmd_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.gcm_tag_data_fifo ;
wire \cddip_decrypt_kop_fifo_override.f.gcm_cmd_fifo ;
wire [31:0] \idle_components.r.part0 ;
wire [19:0] \idle_components.f.num_key_tlvs_in_flight ;
wire \idle_components.f.cddip0_key_tlv_rsm_idle ;
wire \idle_components.f.cddip1_key_tlv_rsm_idle ;
wire \idle_components.f.cddip2_key_tlv_rsm_idle ;
wire \idle_components.f.cddip3_key_tlv_rsm_idle ;
wire \idle_components.f.cceip0_key_tlv_rsm_idle ;
wire \idle_components.f.cceip1_key_tlv_rsm_idle ;
wire \idle_components.f.cceip2_key_tlv_rsm_idle ;
wire \idle_components.f.cceip3_key_tlv_rsm_idle ;
wire \idle_components.f.no_key_tlv_in_flight ;
wire \idle_components.f.tlv_parser_idle ;
wire \idle_components.f.drng_idle ;
wire \idle_components.f.kme_slv_empty ;
wire [0:0] \kim_dout.valid ;
wire [2:0] \kim_dout.label_index ;
wire [1:0] \kim_dout.ckv_length ;
wire [14:0] \kim_dout.ckv_pointer ;
wire [3:0] \kim_dout.pf_num ;
wire [11:0] \kim_dout.vf_num ;
wire [0:0] \kim_dout.vf_valid ;
wire \kme_cceip0_ob_in_mod.tready ;
wire \kme_cceip0_ob_out_pre.tvalid ;
wire \kme_cceip0_ob_out_pre.tlast ;
wire [0:0] \kme_cceip0_ob_out_pre.tid ;
wire [7:0] \kme_cceip0_ob_out_pre.tstrb ;
wire [7:0] \kme_cceip0_ob_out_pre.tuser ;
wire [63:0] \kme_cceip0_ob_out_pre.tdata ;
wire \kme_cceip1_ob_in_mod.tready ;
wire \kme_cceip1_ob_out_pre.tvalid ;
wire \kme_cceip1_ob_out_pre.tlast ;
wire [0:0] \kme_cceip1_ob_out_pre.tid ;
wire [7:0] \kme_cceip1_ob_out_pre.tstrb ;
wire [7:0] \kme_cceip1_ob_out_pre.tuser ;
wire [63:0] \kme_cceip1_ob_out_pre.tdata ;
wire \kme_cceip2_ob_in_mod.tready ;
wire \kme_cceip2_ob_out_pre.tvalid ;
wire \kme_cceip2_ob_out_pre.tlast ;
wire [0:0] \kme_cceip2_ob_out_pre.tid ;
wire [7:0] \kme_cceip2_ob_out_pre.tstrb ;
wire [7:0] \kme_cceip2_ob_out_pre.tuser ;
wire [63:0] \kme_cceip2_ob_out_pre.tdata ;
wire \kme_cceip3_ob_in_mod.tready ;
wire \kme_cceip3_ob_out_pre.tvalid ;
wire \kme_cceip3_ob_out_pre.tlast ;
wire [0:0] \kme_cceip3_ob_out_pre.tid ;
wire [7:0] \kme_cceip3_ob_out_pre.tstrb ;
wire [7:0] \kme_cceip3_ob_out_pre.tuser ;
wire [63:0] \kme_cceip3_ob_out_pre.tdata ;
wire \kme_cddip0_ob_in_mod.tready ;
wire \kme_cddip0_ob_out_pre.tvalid ;
wire \kme_cddip0_ob_out_pre.tlast ;
wire [0:0] \kme_cddip0_ob_out_pre.tid ;
wire [7:0] \kme_cddip0_ob_out_pre.tstrb ;
wire [7:0] \kme_cddip0_ob_out_pre.tuser ;
wire [63:0] \kme_cddip0_ob_out_pre.tdata ;
wire \kme_cddip1_ob_in_mod.tready ;
wire \kme_cddip1_ob_out_pre.tvalid ;
wire \kme_cddip1_ob_out_pre.tlast ;
wire [0:0] \kme_cddip1_ob_out_pre.tid ;
wire [7:0] \kme_cddip1_ob_out_pre.tstrb ;
wire [7:0] \kme_cddip1_ob_out_pre.tuser ;
wire [63:0] \kme_cddip1_ob_out_pre.tdata ;
wire \kme_cddip2_ob_in_mod.tready ;
wire \kme_cddip2_ob_out_pre.tvalid ;
wire \kme_cddip2_ob_out_pre.tlast ;
wire [0:0] \kme_cddip2_ob_out_pre.tid ;
wire [7:0] \kme_cddip2_ob_out_pre.tstrb ;
wire [7:0] \kme_cddip2_ob_out_pre.tuser ;
wire [63:0] \kme_cddip2_ob_out_pre.tdata ;
wire \kme_cddip3_ob_in_mod.tready ;
wire \kme_cddip3_ob_out_pre.tvalid ;
wire \kme_cddip3_ob_out_pre.tlast ;
wire [0:0] \kme_cddip3_ob_out_pre.tid ;
wire [7:0] \kme_cddip3_ob_out_pre.tstrb ;
wire [7:0] \kme_cddip3_ob_out_pre.tuser ;
wire [63:0] \kme_cddip3_ob_out_pre.tdata ;
wire [31:0] \sa_global_ctrl.r.part0 ;
wire [29:0] \sa_global_ctrl.f.spare ;
wire \sa_global_ctrl.f.sa_snap ;
wire \sa_global_ctrl.f.sa_clear_live ;
wire [8:0] \tready_override.r.part0 ;
wire \tready_override.f.txc_tready_override ;
wire \tready_override.f.engine_7_tready_override ;
wire \tready_override.f.engine_6_tready_override ;
wire \tready_override.f.engine_5_tready_override ;
wire \tready_override.f.engine_4_tready_override ;
wire \tready_override.f.engine_3_tready_override ;
wire \tready_override.f.engine_2_tready_override ;
wire \tready_override.f.engine_1_tready_override ;
wire \tready_override.f.engine_0_tready_override ;
tran (kme_ib_in[82], \kme_ib_in.tvalid );
tran (kme_ib_in[81], \kme_ib_in.tlast );
tran (kme_ib_in[80], \kme_ib_in.tid [0]);
tran (kme_ib_in[79], \kme_ib_in.tstrb [7]);
tran (kme_ib_in[78], \kme_ib_in.tstrb [6]);
tran (kme_ib_in[77], \kme_ib_in.tstrb [5]);
tran (kme_ib_in[76], \kme_ib_in.tstrb [4]);
tran (kme_ib_in[75], \kme_ib_in.tstrb [3]);
tran (kme_ib_in[74], \kme_ib_in.tstrb [2]);
tran (kme_ib_in[73], \kme_ib_in.tstrb [1]);
tran (kme_ib_in[72], \kme_ib_in.tstrb [0]);
tran (kme_ib_in[71], \kme_ib_in.tuser [7]);
tran (kme_ib_in[70], \kme_ib_in.tuser [6]);
tran (kme_ib_in[69], \kme_ib_in.tuser [5]);
tran (kme_ib_in[68], \kme_ib_in.tuser [4]);
tran (kme_ib_in[67], \kme_ib_in.tuser [3]);
tran (kme_ib_in[66], \kme_ib_in.tuser [2]);
tran (kme_ib_in[65], \kme_ib_in.tuser [1]);
tran (kme_ib_in[64], \kme_ib_in.tuser [0]);
tran (kme_ib_in[63], \kme_ib_in.tdata [63]);
tran (kme_ib_in[62], \kme_ib_in.tdata [62]);
tran (kme_ib_in[61], \kme_ib_in.tdata [61]);
tran (kme_ib_in[60], \kme_ib_in.tdata [60]);
tran (kme_ib_in[59], \kme_ib_in.tdata [59]);
tran (kme_ib_in[58], \kme_ib_in.tdata [58]);
tran (kme_ib_in[57], \kme_ib_in.tdata [57]);
tran (kme_ib_in[56], \kme_ib_in.tdata [56]);
tran (kme_ib_in[55], \kme_ib_in.tdata [55]);
tran (kme_ib_in[54], \kme_ib_in.tdata [54]);
tran (kme_ib_in[53], \kme_ib_in.tdata [53]);
tran (kme_ib_in[52], \kme_ib_in.tdata [52]);
tran (kme_ib_in[51], \kme_ib_in.tdata [51]);
tran (kme_ib_in[50], \kme_ib_in.tdata [50]);
tran (kme_ib_in[49], \kme_ib_in.tdata [49]);
tran (kme_ib_in[48], \kme_ib_in.tdata [48]);
tran (kme_ib_in[47], \kme_ib_in.tdata [47]);
tran (kme_ib_in[46], \kme_ib_in.tdata [46]);
tran (kme_ib_in[45], \kme_ib_in.tdata [45]);
tran (kme_ib_in[44], \kme_ib_in.tdata [44]);
tran (kme_ib_in[43], \kme_ib_in.tdata [43]);
tran (kme_ib_in[42], \kme_ib_in.tdata [42]);
tran (kme_ib_in[41], \kme_ib_in.tdata [41]);
tran (kme_ib_in[40], \kme_ib_in.tdata [40]);
tran (kme_ib_in[39], \kme_ib_in.tdata [39]);
tran (kme_ib_in[38], \kme_ib_in.tdata [38]);
tran (kme_ib_in[37], \kme_ib_in.tdata [37]);
tran (kme_ib_in[36], \kme_ib_in.tdata [36]);
tran (kme_ib_in[35], \kme_ib_in.tdata [35]);
tran (kme_ib_in[34], \kme_ib_in.tdata [34]);
tran (kme_ib_in[33], \kme_ib_in.tdata [33]);
tran (kme_ib_in[32], \kme_ib_in.tdata [32]);
tran (kme_ib_in[31], \kme_ib_in.tdata [31]);
tran (kme_ib_in[30], \kme_ib_in.tdata [30]);
tran (kme_ib_in[29], \kme_ib_in.tdata [29]);
tran (kme_ib_in[28], \kme_ib_in.tdata [28]);
tran (kme_ib_in[27], \kme_ib_in.tdata [27]);
tran (kme_ib_in[26], \kme_ib_in.tdata [26]);
tran (kme_ib_in[25], \kme_ib_in.tdata [25]);
tran (kme_ib_in[24], \kme_ib_in.tdata [24]);
tran (kme_ib_in[23], \kme_ib_in.tdata [23]);
tran (kme_ib_in[22], \kme_ib_in.tdata [22]);
tran (kme_ib_in[21], \kme_ib_in.tdata [21]);
tran (kme_ib_in[20], \kme_ib_in.tdata [20]);
tran (kme_ib_in[19], \kme_ib_in.tdata [19]);
tran (kme_ib_in[18], \kme_ib_in.tdata [18]);
tran (kme_ib_in[17], \kme_ib_in.tdata [17]);
tran (kme_ib_in[16], \kme_ib_in.tdata [16]);
tran (kme_ib_in[15], \kme_ib_in.tdata [15]);
tran (kme_ib_in[14], \kme_ib_in.tdata [14]);
tran (kme_ib_in[13], \kme_ib_in.tdata [13]);
tran (kme_ib_in[12], \kme_ib_in.tdata [12]);
tran (kme_ib_in[11], \kme_ib_in.tdata [11]);
tran (kme_ib_in[10], \kme_ib_in.tdata [10]);
tran (kme_ib_in[9], \kme_ib_in.tdata [9]);
tran (kme_ib_in[8], \kme_ib_in.tdata [8]);
tran (kme_ib_in[7], \kme_ib_in.tdata [7]);
tran (kme_ib_in[6], \kme_ib_in.tdata [6]);
tran (kme_ib_in[5], \kme_ib_in.tdata [5]);
tran (kme_ib_in[4], \kme_ib_in.tdata [4]);
tran (kme_ib_in[3], \kme_ib_in.tdata [3]);
tran (kme_ib_in[2], \kme_ib_in.tdata [2]);
tran (kme_ib_in[1], \kme_ib_in.tdata [1]);
tran (kme_ib_in[0], \kme_ib_in.tdata [0]);
tran (kme_cceip0_ob_in[0], \kme_cceip0_ob_in.tready );
tran (kme_ib_out[0], \kme_ib_out.tready );
tran (kme_cceip0_ob_out_pre[82], \kme_cceip0_ob_out_pre.tvalid );
tran (kme_cceip0_ob_out_pre[81], \kme_cceip0_ob_out_pre.tlast );
tran (kme_cceip0_ob_out_pre[80], \kme_cceip0_ob_out_pre.tid [0]);
tran (kme_cceip0_ob_out_pre[79], \kme_cceip0_ob_out_pre.tstrb [7]);
tran (kme_cceip0_ob_out_pre[78], \kme_cceip0_ob_out_pre.tstrb [6]);
tran (kme_cceip0_ob_out_pre[77], \kme_cceip0_ob_out_pre.tstrb [5]);
tran (kme_cceip0_ob_out_pre[76], \kme_cceip0_ob_out_pre.tstrb [4]);
tran (kme_cceip0_ob_out_pre[75], \kme_cceip0_ob_out_pre.tstrb [3]);
tran (kme_cceip0_ob_out_pre[74], \kme_cceip0_ob_out_pre.tstrb [2]);
tran (kme_cceip0_ob_out_pre[73], \kme_cceip0_ob_out_pre.tstrb [1]);
tran (kme_cceip0_ob_out_pre[72], \kme_cceip0_ob_out_pre.tstrb [0]);
tran (kme_cceip0_ob_out_pre[71], \kme_cceip0_ob_out_pre.tuser [7]);
tran (kme_cceip0_ob_out_pre[70], \kme_cceip0_ob_out_pre.tuser [6]);
tran (kme_cceip0_ob_out_pre[69], \kme_cceip0_ob_out_pre.tuser [5]);
tran (kme_cceip0_ob_out_pre[68], \kme_cceip0_ob_out_pre.tuser [4]);
tran (kme_cceip0_ob_out_pre[67], \kme_cceip0_ob_out_pre.tuser [3]);
tran (kme_cceip0_ob_out_pre[66], \kme_cceip0_ob_out_pre.tuser [2]);
tran (kme_cceip0_ob_out_pre[65], \kme_cceip0_ob_out_pre.tuser [1]);
tran (kme_cceip0_ob_out_pre[64], \kme_cceip0_ob_out_pre.tuser [0]);
tran (kme_cceip0_ob_out_pre[63], \kme_cceip0_ob_out_pre.tdata [63]);
tran (kme_cceip0_ob_out_pre[62], \kme_cceip0_ob_out_pre.tdata [62]);
tran (kme_cceip0_ob_out_pre[61], \kme_cceip0_ob_out_pre.tdata [61]);
tran (kme_cceip0_ob_out_pre[60], \kme_cceip0_ob_out_pre.tdata [60]);
tran (kme_cceip0_ob_out_pre[59], \kme_cceip0_ob_out_pre.tdata [59]);
tran (kme_cceip0_ob_out_pre[58], \kme_cceip0_ob_out_pre.tdata [58]);
tran (kme_cceip0_ob_out_pre[57], \kme_cceip0_ob_out_pre.tdata [57]);
tran (kme_cceip0_ob_out_pre[56], \kme_cceip0_ob_out_pre.tdata [56]);
tran (kme_cceip0_ob_out_pre[55], \kme_cceip0_ob_out_pre.tdata [55]);
tran (kme_cceip0_ob_out_pre[54], \kme_cceip0_ob_out_pre.tdata [54]);
tran (kme_cceip0_ob_out_pre[53], \kme_cceip0_ob_out_pre.tdata [53]);
tran (kme_cceip0_ob_out_pre[52], \kme_cceip0_ob_out_pre.tdata [52]);
tran (kme_cceip0_ob_out_pre[51], \kme_cceip0_ob_out_pre.tdata [51]);
tran (kme_cceip0_ob_out_pre[50], \kme_cceip0_ob_out_pre.tdata [50]);
tran (kme_cceip0_ob_out_pre[49], \kme_cceip0_ob_out_pre.tdata [49]);
tran (kme_cceip0_ob_out_pre[48], \kme_cceip0_ob_out_pre.tdata [48]);
tran (kme_cceip0_ob_out_pre[47], \kme_cceip0_ob_out_pre.tdata [47]);
tran (kme_cceip0_ob_out_pre[46], \kme_cceip0_ob_out_pre.tdata [46]);
tran (kme_cceip0_ob_out_pre[45], \kme_cceip0_ob_out_pre.tdata [45]);
tran (kme_cceip0_ob_out_pre[44], \kme_cceip0_ob_out_pre.tdata [44]);
tran (kme_cceip0_ob_out_pre[43], \kme_cceip0_ob_out_pre.tdata [43]);
tran (kme_cceip0_ob_out_pre[42], \kme_cceip0_ob_out_pre.tdata [42]);
tran (kme_cceip0_ob_out_pre[41], \kme_cceip0_ob_out_pre.tdata [41]);
tran (kme_cceip0_ob_out_pre[40], \kme_cceip0_ob_out_pre.tdata [40]);
tran (kme_cceip0_ob_out_pre[39], \kme_cceip0_ob_out_pre.tdata [39]);
tran (kme_cceip0_ob_out_pre[38], \kme_cceip0_ob_out_pre.tdata [38]);
tran (kme_cceip0_ob_out_pre[37], \kme_cceip0_ob_out_pre.tdata [37]);
tran (kme_cceip0_ob_out_pre[36], \kme_cceip0_ob_out_pre.tdata [36]);
tran (kme_cceip0_ob_out_pre[35], \kme_cceip0_ob_out_pre.tdata [35]);
tran (kme_cceip0_ob_out_pre[34], \kme_cceip0_ob_out_pre.tdata [34]);
tran (kme_cceip0_ob_out_pre[33], \kme_cceip0_ob_out_pre.tdata [33]);
tran (kme_cceip0_ob_out_pre[32], \kme_cceip0_ob_out_pre.tdata [32]);
tran (kme_cceip0_ob_out_pre[31], \kme_cceip0_ob_out_pre.tdata [31]);
tran (kme_cceip0_ob_out_pre[30], \kme_cceip0_ob_out_pre.tdata [30]);
tran (kme_cceip0_ob_out_pre[29], \kme_cceip0_ob_out_pre.tdata [29]);
tran (kme_cceip0_ob_out_pre[28], \kme_cceip0_ob_out_pre.tdata [28]);
tran (kme_cceip0_ob_out_pre[27], \kme_cceip0_ob_out_pre.tdata [27]);
tran (kme_cceip0_ob_out_pre[26], \kme_cceip0_ob_out_pre.tdata [26]);
tran (kme_cceip0_ob_out_pre[25], \kme_cceip0_ob_out_pre.tdata [25]);
tran (kme_cceip0_ob_out_pre[24], \kme_cceip0_ob_out_pre.tdata [24]);
tran (kme_cceip0_ob_out_pre[23], \kme_cceip0_ob_out_pre.tdata [23]);
tran (kme_cceip0_ob_out_pre[22], \kme_cceip0_ob_out_pre.tdata [22]);
tran (kme_cceip0_ob_out_pre[21], \kme_cceip0_ob_out_pre.tdata [21]);
tran (kme_cceip0_ob_out_pre[20], \kme_cceip0_ob_out_pre.tdata [20]);
tran (kme_cceip0_ob_out_pre[19], \kme_cceip0_ob_out_pre.tdata [19]);
tran (kme_cceip0_ob_out_pre[18], \kme_cceip0_ob_out_pre.tdata [18]);
tran (kme_cceip0_ob_out_pre[17], \kme_cceip0_ob_out_pre.tdata [17]);
tran (kme_cceip0_ob_out_pre[16], \kme_cceip0_ob_out_pre.tdata [16]);
tran (kme_cceip0_ob_out_pre[15], \kme_cceip0_ob_out_pre.tdata [15]);
tran (kme_cceip0_ob_out_pre[14], \kme_cceip0_ob_out_pre.tdata [14]);
tran (kme_cceip0_ob_out_pre[13], \kme_cceip0_ob_out_pre.tdata [13]);
tran (kme_cceip0_ob_out_pre[12], \kme_cceip0_ob_out_pre.tdata [12]);
tran (kme_cceip0_ob_out_pre[11], \kme_cceip0_ob_out_pre.tdata [11]);
tran (kme_cceip0_ob_out_pre[10], \kme_cceip0_ob_out_pre.tdata [10]);
tran (kme_cceip0_ob_out_pre[9], \kme_cceip0_ob_out_pre.tdata [9]);
tran (kme_cceip0_ob_out_pre[8], \kme_cceip0_ob_out_pre.tdata [8]);
tran (kme_cceip0_ob_out_pre[7], \kme_cceip0_ob_out_pre.tdata [7]);
tran (kme_cceip0_ob_out_pre[6], \kme_cceip0_ob_out_pre.tdata [6]);
tran (kme_cceip0_ob_out_pre[5], \kme_cceip0_ob_out_pre.tdata [5]);
tran (kme_cceip0_ob_out_pre[4], \kme_cceip0_ob_out_pre.tdata [4]);
tran (kme_cceip0_ob_out_pre[3], \kme_cceip0_ob_out_pre.tdata [3]);
tran (kme_cceip0_ob_out_pre[2], \kme_cceip0_ob_out_pre.tdata [2]);
tran (kme_cceip0_ob_out_pre[1], \kme_cceip0_ob_out_pre.tdata [1]);
tran (kme_cceip0_ob_out_pre[0], \kme_cceip0_ob_out_pre.tdata [0]);
tran (kme_cceip1_ob_out_pre[82], \kme_cceip1_ob_out_pre.tvalid );
tran (kme_cceip1_ob_out_pre[81], \kme_cceip1_ob_out_pre.tlast );
tran (kme_cceip1_ob_out_pre[80], \kme_cceip1_ob_out_pre.tid [0]);
tran (kme_cceip1_ob_out_pre[79], \kme_cceip1_ob_out_pre.tstrb [7]);
tran (kme_cceip1_ob_out_pre[78], \kme_cceip1_ob_out_pre.tstrb [6]);
tran (kme_cceip1_ob_out_pre[77], \kme_cceip1_ob_out_pre.tstrb [5]);
tran (kme_cceip1_ob_out_pre[76], \kme_cceip1_ob_out_pre.tstrb [4]);
tran (kme_cceip1_ob_out_pre[75], \kme_cceip1_ob_out_pre.tstrb [3]);
tran (kme_cceip1_ob_out_pre[74], \kme_cceip1_ob_out_pre.tstrb [2]);
tran (kme_cceip1_ob_out_pre[73], \kme_cceip1_ob_out_pre.tstrb [1]);
tran (kme_cceip1_ob_out_pre[72], \kme_cceip1_ob_out_pre.tstrb [0]);
tran (kme_cceip1_ob_out_pre[71], \kme_cceip1_ob_out_pre.tuser [7]);
tran (kme_cceip1_ob_out_pre[70], \kme_cceip1_ob_out_pre.tuser [6]);
tran (kme_cceip1_ob_out_pre[69], \kme_cceip1_ob_out_pre.tuser [5]);
tran (kme_cceip1_ob_out_pre[68], \kme_cceip1_ob_out_pre.tuser [4]);
tran (kme_cceip1_ob_out_pre[67], \kme_cceip1_ob_out_pre.tuser [3]);
tran (kme_cceip1_ob_out_pre[66], \kme_cceip1_ob_out_pre.tuser [2]);
tran (kme_cceip1_ob_out_pre[65], \kme_cceip1_ob_out_pre.tuser [1]);
tran (kme_cceip1_ob_out_pre[64], \kme_cceip1_ob_out_pre.tuser [0]);
tran (kme_cceip1_ob_out_pre[63], \kme_cceip1_ob_out_pre.tdata [63]);
tran (kme_cceip1_ob_out_pre[62], \kme_cceip1_ob_out_pre.tdata [62]);
tran (kme_cceip1_ob_out_pre[61], \kme_cceip1_ob_out_pre.tdata [61]);
tran (kme_cceip1_ob_out_pre[60], \kme_cceip1_ob_out_pre.tdata [60]);
tran (kme_cceip1_ob_out_pre[59], \kme_cceip1_ob_out_pre.tdata [59]);
tran (kme_cceip1_ob_out_pre[58], \kme_cceip1_ob_out_pre.tdata [58]);
tran (kme_cceip1_ob_out_pre[57], \kme_cceip1_ob_out_pre.tdata [57]);
tran (kme_cceip1_ob_out_pre[56], \kme_cceip1_ob_out_pre.tdata [56]);
tran (kme_cceip1_ob_out_pre[55], \kme_cceip1_ob_out_pre.tdata [55]);
tran (kme_cceip1_ob_out_pre[54], \kme_cceip1_ob_out_pre.tdata [54]);
tran (kme_cceip1_ob_out_pre[53], \kme_cceip1_ob_out_pre.tdata [53]);
tran (kme_cceip1_ob_out_pre[52], \kme_cceip1_ob_out_pre.tdata [52]);
tran (kme_cceip1_ob_out_pre[51], \kme_cceip1_ob_out_pre.tdata [51]);
tran (kme_cceip1_ob_out_pre[50], \kme_cceip1_ob_out_pre.tdata [50]);
tran (kme_cceip1_ob_out_pre[49], \kme_cceip1_ob_out_pre.tdata [49]);
tran (kme_cceip1_ob_out_pre[48], \kme_cceip1_ob_out_pre.tdata [48]);
tran (kme_cceip1_ob_out_pre[47], \kme_cceip1_ob_out_pre.tdata [47]);
tran (kme_cceip1_ob_out_pre[46], \kme_cceip1_ob_out_pre.tdata [46]);
tran (kme_cceip1_ob_out_pre[45], \kme_cceip1_ob_out_pre.tdata [45]);
tran (kme_cceip1_ob_out_pre[44], \kme_cceip1_ob_out_pre.tdata [44]);
tran (kme_cceip1_ob_out_pre[43], \kme_cceip1_ob_out_pre.tdata [43]);
tran (kme_cceip1_ob_out_pre[42], \kme_cceip1_ob_out_pre.tdata [42]);
tran (kme_cceip1_ob_out_pre[41], \kme_cceip1_ob_out_pre.tdata [41]);
tran (kme_cceip1_ob_out_pre[40], \kme_cceip1_ob_out_pre.tdata [40]);
tran (kme_cceip1_ob_out_pre[39], \kme_cceip1_ob_out_pre.tdata [39]);
tran (kme_cceip1_ob_out_pre[38], \kme_cceip1_ob_out_pre.tdata [38]);
tran (kme_cceip1_ob_out_pre[37], \kme_cceip1_ob_out_pre.tdata [37]);
tran (kme_cceip1_ob_out_pre[36], \kme_cceip1_ob_out_pre.tdata [36]);
tran (kme_cceip1_ob_out_pre[35], \kme_cceip1_ob_out_pre.tdata [35]);
tran (kme_cceip1_ob_out_pre[34], \kme_cceip1_ob_out_pre.tdata [34]);
tran (kme_cceip1_ob_out_pre[33], \kme_cceip1_ob_out_pre.tdata [33]);
tran (kme_cceip1_ob_out_pre[32], \kme_cceip1_ob_out_pre.tdata [32]);
tran (kme_cceip1_ob_out_pre[31], \kme_cceip1_ob_out_pre.tdata [31]);
tran (kme_cceip1_ob_out_pre[30], \kme_cceip1_ob_out_pre.tdata [30]);
tran (kme_cceip1_ob_out_pre[29], \kme_cceip1_ob_out_pre.tdata [29]);
tran (kme_cceip1_ob_out_pre[28], \kme_cceip1_ob_out_pre.tdata [28]);
tran (kme_cceip1_ob_out_pre[27], \kme_cceip1_ob_out_pre.tdata [27]);
tran (kme_cceip1_ob_out_pre[26], \kme_cceip1_ob_out_pre.tdata [26]);
tran (kme_cceip1_ob_out_pre[25], \kme_cceip1_ob_out_pre.tdata [25]);
tran (kme_cceip1_ob_out_pre[24], \kme_cceip1_ob_out_pre.tdata [24]);
tran (kme_cceip1_ob_out_pre[23], \kme_cceip1_ob_out_pre.tdata [23]);
tran (kme_cceip1_ob_out_pre[22], \kme_cceip1_ob_out_pre.tdata [22]);
tran (kme_cceip1_ob_out_pre[21], \kme_cceip1_ob_out_pre.tdata [21]);
tran (kme_cceip1_ob_out_pre[20], \kme_cceip1_ob_out_pre.tdata [20]);
tran (kme_cceip1_ob_out_pre[19], \kme_cceip1_ob_out_pre.tdata [19]);
tran (kme_cceip1_ob_out_pre[18], \kme_cceip1_ob_out_pre.tdata [18]);
tran (kme_cceip1_ob_out_pre[17], \kme_cceip1_ob_out_pre.tdata [17]);
tran (kme_cceip1_ob_out_pre[16], \kme_cceip1_ob_out_pre.tdata [16]);
tran (kme_cceip1_ob_out_pre[15], \kme_cceip1_ob_out_pre.tdata [15]);
tran (kme_cceip1_ob_out_pre[14], \kme_cceip1_ob_out_pre.tdata [14]);
tran (kme_cceip1_ob_out_pre[13], \kme_cceip1_ob_out_pre.tdata [13]);
tran (kme_cceip1_ob_out_pre[12], \kme_cceip1_ob_out_pre.tdata [12]);
tran (kme_cceip1_ob_out_pre[11], \kme_cceip1_ob_out_pre.tdata [11]);
tran (kme_cceip1_ob_out_pre[10], \kme_cceip1_ob_out_pre.tdata [10]);
tran (kme_cceip1_ob_out_pre[9], \kme_cceip1_ob_out_pre.tdata [9]);
tran (kme_cceip1_ob_out_pre[8], \kme_cceip1_ob_out_pre.tdata [8]);
tran (kme_cceip1_ob_out_pre[7], \kme_cceip1_ob_out_pre.tdata [7]);
tran (kme_cceip1_ob_out_pre[6], \kme_cceip1_ob_out_pre.tdata [6]);
tran (kme_cceip1_ob_out_pre[5], \kme_cceip1_ob_out_pre.tdata [5]);
tran (kme_cceip1_ob_out_pre[4], \kme_cceip1_ob_out_pre.tdata [4]);
tran (kme_cceip1_ob_out_pre[3], \kme_cceip1_ob_out_pre.tdata [3]);
tran (kme_cceip1_ob_out_pre[2], \kme_cceip1_ob_out_pre.tdata [2]);
tran (kme_cceip1_ob_out_pre[1], \kme_cceip1_ob_out_pre.tdata [1]);
tran (kme_cceip1_ob_out_pre[0], \kme_cceip1_ob_out_pre.tdata [0]);
tran (kme_cceip2_ob_out_pre[82], \kme_cceip2_ob_out_pre.tvalid );
tran (kme_cceip2_ob_out_pre[81], \kme_cceip2_ob_out_pre.tlast );
tran (kme_cceip2_ob_out_pre[80], \kme_cceip2_ob_out_pre.tid [0]);
tran (kme_cceip2_ob_out_pre[79], \kme_cceip2_ob_out_pre.tstrb [7]);
tran (kme_cceip2_ob_out_pre[78], \kme_cceip2_ob_out_pre.tstrb [6]);
tran (kme_cceip2_ob_out_pre[77], \kme_cceip2_ob_out_pre.tstrb [5]);
tran (kme_cceip2_ob_out_pre[76], \kme_cceip2_ob_out_pre.tstrb [4]);
tran (kme_cceip2_ob_out_pre[75], \kme_cceip2_ob_out_pre.tstrb [3]);
tran (kme_cceip2_ob_out_pre[74], \kme_cceip2_ob_out_pre.tstrb [2]);
tran (kme_cceip2_ob_out_pre[73], \kme_cceip2_ob_out_pre.tstrb [1]);
tran (kme_cceip2_ob_out_pre[72], \kme_cceip2_ob_out_pre.tstrb [0]);
tran (kme_cceip2_ob_out_pre[71], \kme_cceip2_ob_out_pre.tuser [7]);
tran (kme_cceip2_ob_out_pre[70], \kme_cceip2_ob_out_pre.tuser [6]);
tran (kme_cceip2_ob_out_pre[69], \kme_cceip2_ob_out_pre.tuser [5]);
tran (kme_cceip2_ob_out_pre[68], \kme_cceip2_ob_out_pre.tuser [4]);
tran (kme_cceip2_ob_out_pre[67], \kme_cceip2_ob_out_pre.tuser [3]);
tran (kme_cceip2_ob_out_pre[66], \kme_cceip2_ob_out_pre.tuser [2]);
tran (kme_cceip2_ob_out_pre[65], \kme_cceip2_ob_out_pre.tuser [1]);
tran (kme_cceip2_ob_out_pre[64], \kme_cceip2_ob_out_pre.tuser [0]);
tran (kme_cceip2_ob_out_pre[63], \kme_cceip2_ob_out_pre.tdata [63]);
tran (kme_cceip2_ob_out_pre[62], \kme_cceip2_ob_out_pre.tdata [62]);
tran (kme_cceip2_ob_out_pre[61], \kme_cceip2_ob_out_pre.tdata [61]);
tran (kme_cceip2_ob_out_pre[60], \kme_cceip2_ob_out_pre.tdata [60]);
tran (kme_cceip2_ob_out_pre[59], \kme_cceip2_ob_out_pre.tdata [59]);
tran (kme_cceip2_ob_out_pre[58], \kme_cceip2_ob_out_pre.tdata [58]);
tran (kme_cceip2_ob_out_pre[57], \kme_cceip2_ob_out_pre.tdata [57]);
tran (kme_cceip2_ob_out_pre[56], \kme_cceip2_ob_out_pre.tdata [56]);
tran (kme_cceip2_ob_out_pre[55], \kme_cceip2_ob_out_pre.tdata [55]);
tran (kme_cceip2_ob_out_pre[54], \kme_cceip2_ob_out_pre.tdata [54]);
tran (kme_cceip2_ob_out_pre[53], \kme_cceip2_ob_out_pre.tdata [53]);
tran (kme_cceip2_ob_out_pre[52], \kme_cceip2_ob_out_pre.tdata [52]);
tran (kme_cceip2_ob_out_pre[51], \kme_cceip2_ob_out_pre.tdata [51]);
tran (kme_cceip2_ob_out_pre[50], \kme_cceip2_ob_out_pre.tdata [50]);
tran (kme_cceip2_ob_out_pre[49], \kme_cceip2_ob_out_pre.tdata [49]);
tran (kme_cceip2_ob_out_pre[48], \kme_cceip2_ob_out_pre.tdata [48]);
tran (kme_cceip2_ob_out_pre[47], \kme_cceip2_ob_out_pre.tdata [47]);
tran (kme_cceip2_ob_out_pre[46], \kme_cceip2_ob_out_pre.tdata [46]);
tran (kme_cceip2_ob_out_pre[45], \kme_cceip2_ob_out_pre.tdata [45]);
tran (kme_cceip2_ob_out_pre[44], \kme_cceip2_ob_out_pre.tdata [44]);
tran (kme_cceip2_ob_out_pre[43], \kme_cceip2_ob_out_pre.tdata [43]);
tran (kme_cceip2_ob_out_pre[42], \kme_cceip2_ob_out_pre.tdata [42]);
tran (kme_cceip2_ob_out_pre[41], \kme_cceip2_ob_out_pre.tdata [41]);
tran (kme_cceip2_ob_out_pre[40], \kme_cceip2_ob_out_pre.tdata [40]);
tran (kme_cceip2_ob_out_pre[39], \kme_cceip2_ob_out_pre.tdata [39]);
tran (kme_cceip2_ob_out_pre[38], \kme_cceip2_ob_out_pre.tdata [38]);
tran (kme_cceip2_ob_out_pre[37], \kme_cceip2_ob_out_pre.tdata [37]);
tran (kme_cceip2_ob_out_pre[36], \kme_cceip2_ob_out_pre.tdata [36]);
tran (kme_cceip2_ob_out_pre[35], \kme_cceip2_ob_out_pre.tdata [35]);
tran (kme_cceip2_ob_out_pre[34], \kme_cceip2_ob_out_pre.tdata [34]);
tran (kme_cceip2_ob_out_pre[33], \kme_cceip2_ob_out_pre.tdata [33]);
tran (kme_cceip2_ob_out_pre[32], \kme_cceip2_ob_out_pre.tdata [32]);
tran (kme_cceip2_ob_out_pre[31], \kme_cceip2_ob_out_pre.tdata [31]);
tran (kme_cceip2_ob_out_pre[30], \kme_cceip2_ob_out_pre.tdata [30]);
tran (kme_cceip2_ob_out_pre[29], \kme_cceip2_ob_out_pre.tdata [29]);
tran (kme_cceip2_ob_out_pre[28], \kme_cceip2_ob_out_pre.tdata [28]);
tran (kme_cceip2_ob_out_pre[27], \kme_cceip2_ob_out_pre.tdata [27]);
tran (kme_cceip2_ob_out_pre[26], \kme_cceip2_ob_out_pre.tdata [26]);
tran (kme_cceip2_ob_out_pre[25], \kme_cceip2_ob_out_pre.tdata [25]);
tran (kme_cceip2_ob_out_pre[24], \kme_cceip2_ob_out_pre.tdata [24]);
tran (kme_cceip2_ob_out_pre[23], \kme_cceip2_ob_out_pre.tdata [23]);
tran (kme_cceip2_ob_out_pre[22], \kme_cceip2_ob_out_pre.tdata [22]);
tran (kme_cceip2_ob_out_pre[21], \kme_cceip2_ob_out_pre.tdata [21]);
tran (kme_cceip2_ob_out_pre[20], \kme_cceip2_ob_out_pre.tdata [20]);
tran (kme_cceip2_ob_out_pre[19], \kme_cceip2_ob_out_pre.tdata [19]);
tran (kme_cceip2_ob_out_pre[18], \kme_cceip2_ob_out_pre.tdata [18]);
tran (kme_cceip2_ob_out_pre[17], \kme_cceip2_ob_out_pre.tdata [17]);
tran (kme_cceip2_ob_out_pre[16], \kme_cceip2_ob_out_pre.tdata [16]);
tran (kme_cceip2_ob_out_pre[15], \kme_cceip2_ob_out_pre.tdata [15]);
tran (kme_cceip2_ob_out_pre[14], \kme_cceip2_ob_out_pre.tdata [14]);
tran (kme_cceip2_ob_out_pre[13], \kme_cceip2_ob_out_pre.tdata [13]);
tran (kme_cceip2_ob_out_pre[12], \kme_cceip2_ob_out_pre.tdata [12]);
tran (kme_cceip2_ob_out_pre[11], \kme_cceip2_ob_out_pre.tdata [11]);
tran (kme_cceip2_ob_out_pre[10], \kme_cceip2_ob_out_pre.tdata [10]);
tran (kme_cceip2_ob_out_pre[9], \kme_cceip2_ob_out_pre.tdata [9]);
tran (kme_cceip2_ob_out_pre[8], \kme_cceip2_ob_out_pre.tdata [8]);
tran (kme_cceip2_ob_out_pre[7], \kme_cceip2_ob_out_pre.tdata [7]);
tran (kme_cceip2_ob_out_pre[6], \kme_cceip2_ob_out_pre.tdata [6]);
tran (kme_cceip2_ob_out_pre[5], \kme_cceip2_ob_out_pre.tdata [5]);
tran (kme_cceip2_ob_out_pre[4], \kme_cceip2_ob_out_pre.tdata [4]);
tran (kme_cceip2_ob_out_pre[3], \kme_cceip2_ob_out_pre.tdata [3]);
tran (kme_cceip2_ob_out_pre[2], \kme_cceip2_ob_out_pre.tdata [2]);
tran (kme_cceip2_ob_out_pre[1], \kme_cceip2_ob_out_pre.tdata [1]);
tran (kme_cceip2_ob_out_pre[0], \kme_cceip2_ob_out_pre.tdata [0]);
tran (kme_cceip3_ob_out_pre[82], \kme_cceip3_ob_out_pre.tvalid );
tran (kme_cceip3_ob_out_pre[81], \kme_cceip3_ob_out_pre.tlast );
tran (kme_cceip3_ob_out_pre[80], \kme_cceip3_ob_out_pre.tid [0]);
tran (kme_cceip3_ob_out_pre[79], \kme_cceip3_ob_out_pre.tstrb [7]);
tran (kme_cceip3_ob_out_pre[78], \kme_cceip3_ob_out_pre.tstrb [6]);
tran (kme_cceip3_ob_out_pre[77], \kme_cceip3_ob_out_pre.tstrb [5]);
tran (kme_cceip3_ob_out_pre[76], \kme_cceip3_ob_out_pre.tstrb [4]);
tran (kme_cceip3_ob_out_pre[75], \kme_cceip3_ob_out_pre.tstrb [3]);
tran (kme_cceip3_ob_out_pre[74], \kme_cceip3_ob_out_pre.tstrb [2]);
tran (kme_cceip3_ob_out_pre[73], \kme_cceip3_ob_out_pre.tstrb [1]);
tran (kme_cceip3_ob_out_pre[72], \kme_cceip3_ob_out_pre.tstrb [0]);
tran (kme_cceip3_ob_out_pre[71], \kme_cceip3_ob_out_pre.tuser [7]);
tran (kme_cceip3_ob_out_pre[70], \kme_cceip3_ob_out_pre.tuser [6]);
tran (kme_cceip3_ob_out_pre[69], \kme_cceip3_ob_out_pre.tuser [5]);
tran (kme_cceip3_ob_out_pre[68], \kme_cceip3_ob_out_pre.tuser [4]);
tran (kme_cceip3_ob_out_pre[67], \kme_cceip3_ob_out_pre.tuser [3]);
tran (kme_cceip3_ob_out_pre[66], \kme_cceip3_ob_out_pre.tuser [2]);
tran (kme_cceip3_ob_out_pre[65], \kme_cceip3_ob_out_pre.tuser [1]);
tran (kme_cceip3_ob_out_pre[64], \kme_cceip3_ob_out_pre.tuser [0]);
tran (kme_cceip3_ob_out_pre[63], \kme_cceip3_ob_out_pre.tdata [63]);
tran (kme_cceip3_ob_out_pre[62], \kme_cceip3_ob_out_pre.tdata [62]);
tran (kme_cceip3_ob_out_pre[61], \kme_cceip3_ob_out_pre.tdata [61]);
tran (kme_cceip3_ob_out_pre[60], \kme_cceip3_ob_out_pre.tdata [60]);
tran (kme_cceip3_ob_out_pre[59], \kme_cceip3_ob_out_pre.tdata [59]);
tran (kme_cceip3_ob_out_pre[58], \kme_cceip3_ob_out_pre.tdata [58]);
tran (kme_cceip3_ob_out_pre[57], \kme_cceip3_ob_out_pre.tdata [57]);
tran (kme_cceip3_ob_out_pre[56], \kme_cceip3_ob_out_pre.tdata [56]);
tran (kme_cceip3_ob_out_pre[55], \kme_cceip3_ob_out_pre.tdata [55]);
tran (kme_cceip3_ob_out_pre[54], \kme_cceip3_ob_out_pre.tdata [54]);
tran (kme_cceip3_ob_out_pre[53], \kme_cceip3_ob_out_pre.tdata [53]);
tran (kme_cceip3_ob_out_pre[52], \kme_cceip3_ob_out_pre.tdata [52]);
tran (kme_cceip3_ob_out_pre[51], \kme_cceip3_ob_out_pre.tdata [51]);
tran (kme_cceip3_ob_out_pre[50], \kme_cceip3_ob_out_pre.tdata [50]);
tran (kme_cceip3_ob_out_pre[49], \kme_cceip3_ob_out_pre.tdata [49]);
tran (kme_cceip3_ob_out_pre[48], \kme_cceip3_ob_out_pre.tdata [48]);
tran (kme_cceip3_ob_out_pre[47], \kme_cceip3_ob_out_pre.tdata [47]);
tran (kme_cceip3_ob_out_pre[46], \kme_cceip3_ob_out_pre.tdata [46]);
tran (kme_cceip3_ob_out_pre[45], \kme_cceip3_ob_out_pre.tdata [45]);
tran (kme_cceip3_ob_out_pre[44], \kme_cceip3_ob_out_pre.tdata [44]);
tran (kme_cceip3_ob_out_pre[43], \kme_cceip3_ob_out_pre.tdata [43]);
tran (kme_cceip3_ob_out_pre[42], \kme_cceip3_ob_out_pre.tdata [42]);
tran (kme_cceip3_ob_out_pre[41], \kme_cceip3_ob_out_pre.tdata [41]);
tran (kme_cceip3_ob_out_pre[40], \kme_cceip3_ob_out_pre.tdata [40]);
tran (kme_cceip3_ob_out_pre[39], \kme_cceip3_ob_out_pre.tdata [39]);
tran (kme_cceip3_ob_out_pre[38], \kme_cceip3_ob_out_pre.tdata [38]);
tran (kme_cceip3_ob_out_pre[37], \kme_cceip3_ob_out_pre.tdata [37]);
tran (kme_cceip3_ob_out_pre[36], \kme_cceip3_ob_out_pre.tdata [36]);
tran (kme_cceip3_ob_out_pre[35], \kme_cceip3_ob_out_pre.tdata [35]);
tran (kme_cceip3_ob_out_pre[34], \kme_cceip3_ob_out_pre.tdata [34]);
tran (kme_cceip3_ob_out_pre[33], \kme_cceip3_ob_out_pre.tdata [33]);
tran (kme_cceip3_ob_out_pre[32], \kme_cceip3_ob_out_pre.tdata [32]);
tran (kme_cceip3_ob_out_pre[31], \kme_cceip3_ob_out_pre.tdata [31]);
tran (kme_cceip3_ob_out_pre[30], \kme_cceip3_ob_out_pre.tdata [30]);
tran (kme_cceip3_ob_out_pre[29], \kme_cceip3_ob_out_pre.tdata [29]);
tran (kme_cceip3_ob_out_pre[28], \kme_cceip3_ob_out_pre.tdata [28]);
tran (kme_cceip3_ob_out_pre[27], \kme_cceip3_ob_out_pre.tdata [27]);
tran (kme_cceip3_ob_out_pre[26], \kme_cceip3_ob_out_pre.tdata [26]);
tran (kme_cceip3_ob_out_pre[25], \kme_cceip3_ob_out_pre.tdata [25]);
tran (kme_cceip3_ob_out_pre[24], \kme_cceip3_ob_out_pre.tdata [24]);
tran (kme_cceip3_ob_out_pre[23], \kme_cceip3_ob_out_pre.tdata [23]);
tran (kme_cceip3_ob_out_pre[22], \kme_cceip3_ob_out_pre.tdata [22]);
tran (kme_cceip3_ob_out_pre[21], \kme_cceip3_ob_out_pre.tdata [21]);
tran (kme_cceip3_ob_out_pre[20], \kme_cceip3_ob_out_pre.tdata [20]);
tran (kme_cceip3_ob_out_pre[19], \kme_cceip3_ob_out_pre.tdata [19]);
tran (kme_cceip3_ob_out_pre[18], \kme_cceip3_ob_out_pre.tdata [18]);
tran (kme_cceip3_ob_out_pre[17], \kme_cceip3_ob_out_pre.tdata [17]);
tran (kme_cceip3_ob_out_pre[16], \kme_cceip3_ob_out_pre.tdata [16]);
tran (kme_cceip3_ob_out_pre[15], \kme_cceip3_ob_out_pre.tdata [15]);
tran (kme_cceip3_ob_out_pre[14], \kme_cceip3_ob_out_pre.tdata [14]);
tran (kme_cceip3_ob_out_pre[13], \kme_cceip3_ob_out_pre.tdata [13]);
tran (kme_cceip3_ob_out_pre[12], \kme_cceip3_ob_out_pre.tdata [12]);
tran (kme_cceip3_ob_out_pre[11], \kme_cceip3_ob_out_pre.tdata [11]);
tran (kme_cceip3_ob_out_pre[10], \kme_cceip3_ob_out_pre.tdata [10]);
tran (kme_cceip3_ob_out_pre[9], \kme_cceip3_ob_out_pre.tdata [9]);
tran (kme_cceip3_ob_out_pre[8], \kme_cceip3_ob_out_pre.tdata [8]);
tran (kme_cceip3_ob_out_pre[7], \kme_cceip3_ob_out_pre.tdata [7]);
tran (kme_cceip3_ob_out_pre[6], \kme_cceip3_ob_out_pre.tdata [6]);
tran (kme_cceip3_ob_out_pre[5], \kme_cceip3_ob_out_pre.tdata [5]);
tran (kme_cceip3_ob_out_pre[4], \kme_cceip3_ob_out_pre.tdata [4]);
tran (kme_cceip3_ob_out_pre[3], \kme_cceip3_ob_out_pre.tdata [3]);
tran (kme_cceip3_ob_out_pre[2], \kme_cceip3_ob_out_pre.tdata [2]);
tran (kme_cceip3_ob_out_pre[1], \kme_cceip3_ob_out_pre.tdata [1]);
tran (kme_cceip3_ob_out_pre[0], \kme_cceip3_ob_out_pre.tdata [0]);
tran (kme_cddip0_ob_out_pre[82], \kme_cddip0_ob_out_pre.tvalid );
tran (kme_cddip0_ob_out_pre[81], \kme_cddip0_ob_out_pre.tlast );
tran (kme_cddip0_ob_out_pre[80], \kme_cddip0_ob_out_pre.tid [0]);
tran (kme_cddip0_ob_out_pre[79], \kme_cddip0_ob_out_pre.tstrb [7]);
tran (kme_cddip0_ob_out_pre[78], \kme_cddip0_ob_out_pre.tstrb [6]);
tran (kme_cddip0_ob_out_pre[77], \kme_cddip0_ob_out_pre.tstrb [5]);
tran (kme_cddip0_ob_out_pre[76], \kme_cddip0_ob_out_pre.tstrb [4]);
tran (kme_cddip0_ob_out_pre[75], \kme_cddip0_ob_out_pre.tstrb [3]);
tran (kme_cddip0_ob_out_pre[74], \kme_cddip0_ob_out_pre.tstrb [2]);
tran (kme_cddip0_ob_out_pre[73], \kme_cddip0_ob_out_pre.tstrb [1]);
tran (kme_cddip0_ob_out_pre[72], \kme_cddip0_ob_out_pre.tstrb [0]);
tran (kme_cddip0_ob_out_pre[71], \kme_cddip0_ob_out_pre.tuser [7]);
tran (kme_cddip0_ob_out_pre[70], \kme_cddip0_ob_out_pre.tuser [6]);
tran (kme_cddip0_ob_out_pre[69], \kme_cddip0_ob_out_pre.tuser [5]);
tran (kme_cddip0_ob_out_pre[68], \kme_cddip0_ob_out_pre.tuser [4]);
tran (kme_cddip0_ob_out_pre[67], \kme_cddip0_ob_out_pre.tuser [3]);
tran (kme_cddip0_ob_out_pre[66], \kme_cddip0_ob_out_pre.tuser [2]);
tran (kme_cddip0_ob_out_pre[65], \kme_cddip0_ob_out_pre.tuser [1]);
tran (kme_cddip0_ob_out_pre[64], \kme_cddip0_ob_out_pre.tuser [0]);
tran (kme_cddip0_ob_out_pre[63], \kme_cddip0_ob_out_pre.tdata [63]);
tran (kme_cddip0_ob_out_pre[62], \kme_cddip0_ob_out_pre.tdata [62]);
tran (kme_cddip0_ob_out_pre[61], \kme_cddip0_ob_out_pre.tdata [61]);
tran (kme_cddip0_ob_out_pre[60], \kme_cddip0_ob_out_pre.tdata [60]);
tran (kme_cddip0_ob_out_pre[59], \kme_cddip0_ob_out_pre.tdata [59]);
tran (kme_cddip0_ob_out_pre[58], \kme_cddip0_ob_out_pre.tdata [58]);
tran (kme_cddip0_ob_out_pre[57], \kme_cddip0_ob_out_pre.tdata [57]);
tran (kme_cddip0_ob_out_pre[56], \kme_cddip0_ob_out_pre.tdata [56]);
tran (kme_cddip0_ob_out_pre[55], \kme_cddip0_ob_out_pre.tdata [55]);
tran (kme_cddip0_ob_out_pre[54], \kme_cddip0_ob_out_pre.tdata [54]);
tran (kme_cddip0_ob_out_pre[53], \kme_cddip0_ob_out_pre.tdata [53]);
tran (kme_cddip0_ob_out_pre[52], \kme_cddip0_ob_out_pre.tdata [52]);
tran (kme_cddip0_ob_out_pre[51], \kme_cddip0_ob_out_pre.tdata [51]);
tran (kme_cddip0_ob_out_pre[50], \kme_cddip0_ob_out_pre.tdata [50]);
tran (kme_cddip0_ob_out_pre[49], \kme_cddip0_ob_out_pre.tdata [49]);
tran (kme_cddip0_ob_out_pre[48], \kme_cddip0_ob_out_pre.tdata [48]);
tran (kme_cddip0_ob_out_pre[47], \kme_cddip0_ob_out_pre.tdata [47]);
tran (kme_cddip0_ob_out_pre[46], \kme_cddip0_ob_out_pre.tdata [46]);
tran (kme_cddip0_ob_out_pre[45], \kme_cddip0_ob_out_pre.tdata [45]);
tran (kme_cddip0_ob_out_pre[44], \kme_cddip0_ob_out_pre.tdata [44]);
tran (kme_cddip0_ob_out_pre[43], \kme_cddip0_ob_out_pre.tdata [43]);
tran (kme_cddip0_ob_out_pre[42], \kme_cddip0_ob_out_pre.tdata [42]);
tran (kme_cddip0_ob_out_pre[41], \kme_cddip0_ob_out_pre.tdata [41]);
tran (kme_cddip0_ob_out_pre[40], \kme_cddip0_ob_out_pre.tdata [40]);
tran (kme_cddip0_ob_out_pre[39], \kme_cddip0_ob_out_pre.tdata [39]);
tran (kme_cddip0_ob_out_pre[38], \kme_cddip0_ob_out_pre.tdata [38]);
tran (kme_cddip0_ob_out_pre[37], \kme_cddip0_ob_out_pre.tdata [37]);
tran (kme_cddip0_ob_out_pre[36], \kme_cddip0_ob_out_pre.tdata [36]);
tran (kme_cddip0_ob_out_pre[35], \kme_cddip0_ob_out_pre.tdata [35]);
tran (kme_cddip0_ob_out_pre[34], \kme_cddip0_ob_out_pre.tdata [34]);
tran (kme_cddip0_ob_out_pre[33], \kme_cddip0_ob_out_pre.tdata [33]);
tran (kme_cddip0_ob_out_pre[32], \kme_cddip0_ob_out_pre.tdata [32]);
tran (kme_cddip0_ob_out_pre[31], \kme_cddip0_ob_out_pre.tdata [31]);
tran (kme_cddip0_ob_out_pre[30], \kme_cddip0_ob_out_pre.tdata [30]);
tran (kme_cddip0_ob_out_pre[29], \kme_cddip0_ob_out_pre.tdata [29]);
tran (kme_cddip0_ob_out_pre[28], \kme_cddip0_ob_out_pre.tdata [28]);
tran (kme_cddip0_ob_out_pre[27], \kme_cddip0_ob_out_pre.tdata [27]);
tran (kme_cddip0_ob_out_pre[26], \kme_cddip0_ob_out_pre.tdata [26]);
tran (kme_cddip0_ob_out_pre[25], \kme_cddip0_ob_out_pre.tdata [25]);
tran (kme_cddip0_ob_out_pre[24], \kme_cddip0_ob_out_pre.tdata [24]);
tran (kme_cddip0_ob_out_pre[23], \kme_cddip0_ob_out_pre.tdata [23]);
tran (kme_cddip0_ob_out_pre[22], \kme_cddip0_ob_out_pre.tdata [22]);
tran (kme_cddip0_ob_out_pre[21], \kme_cddip0_ob_out_pre.tdata [21]);
tran (kme_cddip0_ob_out_pre[20], \kme_cddip0_ob_out_pre.tdata [20]);
tran (kme_cddip0_ob_out_pre[19], \kme_cddip0_ob_out_pre.tdata [19]);
tran (kme_cddip0_ob_out_pre[18], \kme_cddip0_ob_out_pre.tdata [18]);
tran (kme_cddip0_ob_out_pre[17], \kme_cddip0_ob_out_pre.tdata [17]);
tran (kme_cddip0_ob_out_pre[16], \kme_cddip0_ob_out_pre.tdata [16]);
tran (kme_cddip0_ob_out_pre[15], \kme_cddip0_ob_out_pre.tdata [15]);
tran (kme_cddip0_ob_out_pre[14], \kme_cddip0_ob_out_pre.tdata [14]);
tran (kme_cddip0_ob_out_pre[13], \kme_cddip0_ob_out_pre.tdata [13]);
tran (kme_cddip0_ob_out_pre[12], \kme_cddip0_ob_out_pre.tdata [12]);
tran (kme_cddip0_ob_out_pre[11], \kme_cddip0_ob_out_pre.tdata [11]);
tran (kme_cddip0_ob_out_pre[10], \kme_cddip0_ob_out_pre.tdata [10]);
tran (kme_cddip0_ob_out_pre[9], \kme_cddip0_ob_out_pre.tdata [9]);
tran (kme_cddip0_ob_out_pre[8], \kme_cddip0_ob_out_pre.tdata [8]);
tran (kme_cddip0_ob_out_pre[7], \kme_cddip0_ob_out_pre.tdata [7]);
tran (kme_cddip0_ob_out_pre[6], \kme_cddip0_ob_out_pre.tdata [6]);
tran (kme_cddip0_ob_out_pre[5], \kme_cddip0_ob_out_pre.tdata [5]);
tran (kme_cddip0_ob_out_pre[4], \kme_cddip0_ob_out_pre.tdata [4]);
tran (kme_cddip0_ob_out_pre[3], \kme_cddip0_ob_out_pre.tdata [3]);
tran (kme_cddip0_ob_out_pre[2], \kme_cddip0_ob_out_pre.tdata [2]);
tran (kme_cddip0_ob_out_pre[1], \kme_cddip0_ob_out_pre.tdata [1]);
tran (kme_cddip0_ob_out_pre[0], \kme_cddip0_ob_out_pre.tdata [0]);
tran (kme_cddip1_ob_out_pre[82], \kme_cddip1_ob_out_pre.tvalid );
tran (kme_cddip1_ob_out_pre[81], \kme_cddip1_ob_out_pre.tlast );
tran (kme_cddip1_ob_out_pre[80], \kme_cddip1_ob_out_pre.tid [0]);
tran (kme_cddip1_ob_out_pre[79], \kme_cddip1_ob_out_pre.tstrb [7]);
tran (kme_cddip1_ob_out_pre[78], \kme_cddip1_ob_out_pre.tstrb [6]);
tran (kme_cddip1_ob_out_pre[77], \kme_cddip1_ob_out_pre.tstrb [5]);
tran (kme_cddip1_ob_out_pre[76], \kme_cddip1_ob_out_pre.tstrb [4]);
tran (kme_cddip1_ob_out_pre[75], \kme_cddip1_ob_out_pre.tstrb [3]);
tran (kme_cddip1_ob_out_pre[74], \kme_cddip1_ob_out_pre.tstrb [2]);
tran (kme_cddip1_ob_out_pre[73], \kme_cddip1_ob_out_pre.tstrb [1]);
tran (kme_cddip1_ob_out_pre[72], \kme_cddip1_ob_out_pre.tstrb [0]);
tran (kme_cddip1_ob_out_pre[71], \kme_cddip1_ob_out_pre.tuser [7]);
tran (kme_cddip1_ob_out_pre[70], \kme_cddip1_ob_out_pre.tuser [6]);
tran (kme_cddip1_ob_out_pre[69], \kme_cddip1_ob_out_pre.tuser [5]);
tran (kme_cddip1_ob_out_pre[68], \kme_cddip1_ob_out_pre.tuser [4]);
tran (kme_cddip1_ob_out_pre[67], \kme_cddip1_ob_out_pre.tuser [3]);
tran (kme_cddip1_ob_out_pre[66], \kme_cddip1_ob_out_pre.tuser [2]);
tran (kme_cddip1_ob_out_pre[65], \kme_cddip1_ob_out_pre.tuser [1]);
tran (kme_cddip1_ob_out_pre[64], \kme_cddip1_ob_out_pre.tuser [0]);
tran (kme_cddip1_ob_out_pre[63], \kme_cddip1_ob_out_pre.tdata [63]);
tran (kme_cddip1_ob_out_pre[62], \kme_cddip1_ob_out_pre.tdata [62]);
tran (kme_cddip1_ob_out_pre[61], \kme_cddip1_ob_out_pre.tdata [61]);
tran (kme_cddip1_ob_out_pre[60], \kme_cddip1_ob_out_pre.tdata [60]);
tran (kme_cddip1_ob_out_pre[59], \kme_cddip1_ob_out_pre.tdata [59]);
tran (kme_cddip1_ob_out_pre[58], \kme_cddip1_ob_out_pre.tdata [58]);
tran (kme_cddip1_ob_out_pre[57], \kme_cddip1_ob_out_pre.tdata [57]);
tran (kme_cddip1_ob_out_pre[56], \kme_cddip1_ob_out_pre.tdata [56]);
tran (kme_cddip1_ob_out_pre[55], \kme_cddip1_ob_out_pre.tdata [55]);
tran (kme_cddip1_ob_out_pre[54], \kme_cddip1_ob_out_pre.tdata [54]);
tran (kme_cddip1_ob_out_pre[53], \kme_cddip1_ob_out_pre.tdata [53]);
tran (kme_cddip1_ob_out_pre[52], \kme_cddip1_ob_out_pre.tdata [52]);
tran (kme_cddip1_ob_out_pre[51], \kme_cddip1_ob_out_pre.tdata [51]);
tran (kme_cddip1_ob_out_pre[50], \kme_cddip1_ob_out_pre.tdata [50]);
tran (kme_cddip1_ob_out_pre[49], \kme_cddip1_ob_out_pre.tdata [49]);
tran (kme_cddip1_ob_out_pre[48], \kme_cddip1_ob_out_pre.tdata [48]);
tran (kme_cddip1_ob_out_pre[47], \kme_cddip1_ob_out_pre.tdata [47]);
tran (kme_cddip1_ob_out_pre[46], \kme_cddip1_ob_out_pre.tdata [46]);
tran (kme_cddip1_ob_out_pre[45], \kme_cddip1_ob_out_pre.tdata [45]);
tran (kme_cddip1_ob_out_pre[44], \kme_cddip1_ob_out_pre.tdata [44]);
tran (kme_cddip1_ob_out_pre[43], \kme_cddip1_ob_out_pre.tdata [43]);
tran (kme_cddip1_ob_out_pre[42], \kme_cddip1_ob_out_pre.tdata [42]);
tran (kme_cddip1_ob_out_pre[41], \kme_cddip1_ob_out_pre.tdata [41]);
tran (kme_cddip1_ob_out_pre[40], \kme_cddip1_ob_out_pre.tdata [40]);
tran (kme_cddip1_ob_out_pre[39], \kme_cddip1_ob_out_pre.tdata [39]);
tran (kme_cddip1_ob_out_pre[38], \kme_cddip1_ob_out_pre.tdata [38]);
tran (kme_cddip1_ob_out_pre[37], \kme_cddip1_ob_out_pre.tdata [37]);
tran (kme_cddip1_ob_out_pre[36], \kme_cddip1_ob_out_pre.tdata [36]);
tran (kme_cddip1_ob_out_pre[35], \kme_cddip1_ob_out_pre.tdata [35]);
tran (kme_cddip1_ob_out_pre[34], \kme_cddip1_ob_out_pre.tdata [34]);
tran (kme_cddip1_ob_out_pre[33], \kme_cddip1_ob_out_pre.tdata [33]);
tran (kme_cddip1_ob_out_pre[32], \kme_cddip1_ob_out_pre.tdata [32]);
tran (kme_cddip1_ob_out_pre[31], \kme_cddip1_ob_out_pre.tdata [31]);
tran (kme_cddip1_ob_out_pre[30], \kme_cddip1_ob_out_pre.tdata [30]);
tran (kme_cddip1_ob_out_pre[29], \kme_cddip1_ob_out_pre.tdata [29]);
tran (kme_cddip1_ob_out_pre[28], \kme_cddip1_ob_out_pre.tdata [28]);
tran (kme_cddip1_ob_out_pre[27], \kme_cddip1_ob_out_pre.tdata [27]);
tran (kme_cddip1_ob_out_pre[26], \kme_cddip1_ob_out_pre.tdata [26]);
tran (kme_cddip1_ob_out_pre[25], \kme_cddip1_ob_out_pre.tdata [25]);
tran (kme_cddip1_ob_out_pre[24], \kme_cddip1_ob_out_pre.tdata [24]);
tran (kme_cddip1_ob_out_pre[23], \kme_cddip1_ob_out_pre.tdata [23]);
tran (kme_cddip1_ob_out_pre[22], \kme_cddip1_ob_out_pre.tdata [22]);
tran (kme_cddip1_ob_out_pre[21], \kme_cddip1_ob_out_pre.tdata [21]);
tran (kme_cddip1_ob_out_pre[20], \kme_cddip1_ob_out_pre.tdata [20]);
tran (kme_cddip1_ob_out_pre[19], \kme_cddip1_ob_out_pre.tdata [19]);
tran (kme_cddip1_ob_out_pre[18], \kme_cddip1_ob_out_pre.tdata [18]);
tran (kme_cddip1_ob_out_pre[17], \kme_cddip1_ob_out_pre.tdata [17]);
tran (kme_cddip1_ob_out_pre[16], \kme_cddip1_ob_out_pre.tdata [16]);
tran (kme_cddip1_ob_out_pre[15], \kme_cddip1_ob_out_pre.tdata [15]);
tran (kme_cddip1_ob_out_pre[14], \kme_cddip1_ob_out_pre.tdata [14]);
tran (kme_cddip1_ob_out_pre[13], \kme_cddip1_ob_out_pre.tdata [13]);
tran (kme_cddip1_ob_out_pre[12], \kme_cddip1_ob_out_pre.tdata [12]);
tran (kme_cddip1_ob_out_pre[11], \kme_cddip1_ob_out_pre.tdata [11]);
tran (kme_cddip1_ob_out_pre[10], \kme_cddip1_ob_out_pre.tdata [10]);
tran (kme_cddip1_ob_out_pre[9], \kme_cddip1_ob_out_pre.tdata [9]);
tran (kme_cddip1_ob_out_pre[8], \kme_cddip1_ob_out_pre.tdata [8]);
tran (kme_cddip1_ob_out_pre[7], \kme_cddip1_ob_out_pre.tdata [7]);
tran (kme_cddip1_ob_out_pre[6], \kme_cddip1_ob_out_pre.tdata [6]);
tran (kme_cddip1_ob_out_pre[5], \kme_cddip1_ob_out_pre.tdata [5]);
tran (kme_cddip1_ob_out_pre[4], \kme_cddip1_ob_out_pre.tdata [4]);
tran (kme_cddip1_ob_out_pre[3], \kme_cddip1_ob_out_pre.tdata [3]);
tran (kme_cddip1_ob_out_pre[2], \kme_cddip1_ob_out_pre.tdata [2]);
tran (kme_cddip1_ob_out_pre[1], \kme_cddip1_ob_out_pre.tdata [1]);
tran (kme_cddip1_ob_out_pre[0], \kme_cddip1_ob_out_pre.tdata [0]);
tran (kme_cddip2_ob_out_pre[82], \kme_cddip2_ob_out_pre.tvalid );
tran (kme_cddip2_ob_out_pre[81], \kme_cddip2_ob_out_pre.tlast );
tran (kme_cddip2_ob_out_pre[80], \kme_cddip2_ob_out_pre.tid [0]);
tran (kme_cddip2_ob_out_pre[79], \kme_cddip2_ob_out_pre.tstrb [7]);
tran (kme_cddip2_ob_out_pre[78], \kme_cddip2_ob_out_pre.tstrb [6]);
tran (kme_cddip2_ob_out_pre[77], \kme_cddip2_ob_out_pre.tstrb [5]);
tran (kme_cddip2_ob_out_pre[76], \kme_cddip2_ob_out_pre.tstrb [4]);
tran (kme_cddip2_ob_out_pre[75], \kme_cddip2_ob_out_pre.tstrb [3]);
tran (kme_cddip2_ob_out_pre[74], \kme_cddip2_ob_out_pre.tstrb [2]);
tran (kme_cddip2_ob_out_pre[73], \kme_cddip2_ob_out_pre.tstrb [1]);
tran (kme_cddip2_ob_out_pre[72], \kme_cddip2_ob_out_pre.tstrb [0]);
tran (kme_cddip2_ob_out_pre[71], \kme_cddip2_ob_out_pre.tuser [7]);
tran (kme_cddip2_ob_out_pre[70], \kme_cddip2_ob_out_pre.tuser [6]);
tran (kme_cddip2_ob_out_pre[69], \kme_cddip2_ob_out_pre.tuser [5]);
tran (kme_cddip2_ob_out_pre[68], \kme_cddip2_ob_out_pre.tuser [4]);
tran (kme_cddip2_ob_out_pre[67], \kme_cddip2_ob_out_pre.tuser [3]);
tran (kme_cddip2_ob_out_pre[66], \kme_cddip2_ob_out_pre.tuser [2]);
tran (kme_cddip2_ob_out_pre[65], \kme_cddip2_ob_out_pre.tuser [1]);
tran (kme_cddip2_ob_out_pre[64], \kme_cddip2_ob_out_pre.tuser [0]);
tran (kme_cddip2_ob_out_pre[63], \kme_cddip2_ob_out_pre.tdata [63]);
tran (kme_cddip2_ob_out_pre[62], \kme_cddip2_ob_out_pre.tdata [62]);
tran (kme_cddip2_ob_out_pre[61], \kme_cddip2_ob_out_pre.tdata [61]);
tran (kme_cddip2_ob_out_pre[60], \kme_cddip2_ob_out_pre.tdata [60]);
tran (kme_cddip2_ob_out_pre[59], \kme_cddip2_ob_out_pre.tdata [59]);
tran (kme_cddip2_ob_out_pre[58], \kme_cddip2_ob_out_pre.tdata [58]);
tran (kme_cddip2_ob_out_pre[57], \kme_cddip2_ob_out_pre.tdata [57]);
tran (kme_cddip2_ob_out_pre[56], \kme_cddip2_ob_out_pre.tdata [56]);
tran (kme_cddip2_ob_out_pre[55], \kme_cddip2_ob_out_pre.tdata [55]);
tran (kme_cddip2_ob_out_pre[54], \kme_cddip2_ob_out_pre.tdata [54]);
tran (kme_cddip2_ob_out_pre[53], \kme_cddip2_ob_out_pre.tdata [53]);
tran (kme_cddip2_ob_out_pre[52], \kme_cddip2_ob_out_pre.tdata [52]);
tran (kme_cddip2_ob_out_pre[51], \kme_cddip2_ob_out_pre.tdata [51]);
tran (kme_cddip2_ob_out_pre[50], \kme_cddip2_ob_out_pre.tdata [50]);
tran (kme_cddip2_ob_out_pre[49], \kme_cddip2_ob_out_pre.tdata [49]);
tran (kme_cddip2_ob_out_pre[48], \kme_cddip2_ob_out_pre.tdata [48]);
tran (kme_cddip2_ob_out_pre[47], \kme_cddip2_ob_out_pre.tdata [47]);
tran (kme_cddip2_ob_out_pre[46], \kme_cddip2_ob_out_pre.tdata [46]);
tran (kme_cddip2_ob_out_pre[45], \kme_cddip2_ob_out_pre.tdata [45]);
tran (kme_cddip2_ob_out_pre[44], \kme_cddip2_ob_out_pre.tdata [44]);
tran (kme_cddip2_ob_out_pre[43], \kme_cddip2_ob_out_pre.tdata [43]);
tran (kme_cddip2_ob_out_pre[42], \kme_cddip2_ob_out_pre.tdata [42]);
tran (kme_cddip2_ob_out_pre[41], \kme_cddip2_ob_out_pre.tdata [41]);
tran (kme_cddip2_ob_out_pre[40], \kme_cddip2_ob_out_pre.tdata [40]);
tran (kme_cddip2_ob_out_pre[39], \kme_cddip2_ob_out_pre.tdata [39]);
tran (kme_cddip2_ob_out_pre[38], \kme_cddip2_ob_out_pre.tdata [38]);
tran (kme_cddip2_ob_out_pre[37], \kme_cddip2_ob_out_pre.tdata [37]);
tran (kme_cddip2_ob_out_pre[36], \kme_cddip2_ob_out_pre.tdata [36]);
tran (kme_cddip2_ob_out_pre[35], \kme_cddip2_ob_out_pre.tdata [35]);
tran (kme_cddip2_ob_out_pre[34], \kme_cddip2_ob_out_pre.tdata [34]);
tran (kme_cddip2_ob_out_pre[33], \kme_cddip2_ob_out_pre.tdata [33]);
tran (kme_cddip2_ob_out_pre[32], \kme_cddip2_ob_out_pre.tdata [32]);
tran (kme_cddip2_ob_out_pre[31], \kme_cddip2_ob_out_pre.tdata [31]);
tran (kme_cddip2_ob_out_pre[30], \kme_cddip2_ob_out_pre.tdata [30]);
tran (kme_cddip2_ob_out_pre[29], \kme_cddip2_ob_out_pre.tdata [29]);
tran (kme_cddip2_ob_out_pre[28], \kme_cddip2_ob_out_pre.tdata [28]);
tran (kme_cddip2_ob_out_pre[27], \kme_cddip2_ob_out_pre.tdata [27]);
tran (kme_cddip2_ob_out_pre[26], \kme_cddip2_ob_out_pre.tdata [26]);
tran (kme_cddip2_ob_out_pre[25], \kme_cddip2_ob_out_pre.tdata [25]);
tran (kme_cddip2_ob_out_pre[24], \kme_cddip2_ob_out_pre.tdata [24]);
tran (kme_cddip2_ob_out_pre[23], \kme_cddip2_ob_out_pre.tdata [23]);
tran (kme_cddip2_ob_out_pre[22], \kme_cddip2_ob_out_pre.tdata [22]);
tran (kme_cddip2_ob_out_pre[21], \kme_cddip2_ob_out_pre.tdata [21]);
tran (kme_cddip2_ob_out_pre[20], \kme_cddip2_ob_out_pre.tdata [20]);
tran (kme_cddip2_ob_out_pre[19], \kme_cddip2_ob_out_pre.tdata [19]);
tran (kme_cddip2_ob_out_pre[18], \kme_cddip2_ob_out_pre.tdata [18]);
tran (kme_cddip2_ob_out_pre[17], \kme_cddip2_ob_out_pre.tdata [17]);
tran (kme_cddip2_ob_out_pre[16], \kme_cddip2_ob_out_pre.tdata [16]);
tran (kme_cddip2_ob_out_pre[15], \kme_cddip2_ob_out_pre.tdata [15]);
tran (kme_cddip2_ob_out_pre[14], \kme_cddip2_ob_out_pre.tdata [14]);
tran (kme_cddip2_ob_out_pre[13], \kme_cddip2_ob_out_pre.tdata [13]);
tran (kme_cddip2_ob_out_pre[12], \kme_cddip2_ob_out_pre.tdata [12]);
tran (kme_cddip2_ob_out_pre[11], \kme_cddip2_ob_out_pre.tdata [11]);
tran (kme_cddip2_ob_out_pre[10], \kme_cddip2_ob_out_pre.tdata [10]);
tran (kme_cddip2_ob_out_pre[9], \kme_cddip2_ob_out_pre.tdata [9]);
tran (kme_cddip2_ob_out_pre[8], \kme_cddip2_ob_out_pre.tdata [8]);
tran (kme_cddip2_ob_out_pre[7], \kme_cddip2_ob_out_pre.tdata [7]);
tran (kme_cddip2_ob_out_pre[6], \kme_cddip2_ob_out_pre.tdata [6]);
tran (kme_cddip2_ob_out_pre[5], \kme_cddip2_ob_out_pre.tdata [5]);
tran (kme_cddip2_ob_out_pre[4], \kme_cddip2_ob_out_pre.tdata [4]);
tran (kme_cddip2_ob_out_pre[3], \kme_cddip2_ob_out_pre.tdata [3]);
tran (kme_cddip2_ob_out_pre[2], \kme_cddip2_ob_out_pre.tdata [2]);
tran (kme_cddip2_ob_out_pre[1], \kme_cddip2_ob_out_pre.tdata [1]);
tran (kme_cddip2_ob_out_pre[0], \kme_cddip2_ob_out_pre.tdata [0]);
tran (kme_cddip3_ob_out_pre[82], \kme_cddip3_ob_out_pre.tvalid );
tran (kme_cddip3_ob_out_pre[81], \kme_cddip3_ob_out_pre.tlast );
tran (kme_cddip3_ob_out_pre[80], \kme_cddip3_ob_out_pre.tid [0]);
tran (kme_cddip3_ob_out_pre[79], \kme_cddip3_ob_out_pre.tstrb [7]);
tran (kme_cddip3_ob_out_pre[78], \kme_cddip3_ob_out_pre.tstrb [6]);
tran (kme_cddip3_ob_out_pre[77], \kme_cddip3_ob_out_pre.tstrb [5]);
tran (kme_cddip3_ob_out_pre[76], \kme_cddip3_ob_out_pre.tstrb [4]);
tran (kme_cddip3_ob_out_pre[75], \kme_cddip3_ob_out_pre.tstrb [3]);
tran (kme_cddip3_ob_out_pre[74], \kme_cddip3_ob_out_pre.tstrb [2]);
tran (kme_cddip3_ob_out_pre[73], \kme_cddip3_ob_out_pre.tstrb [1]);
tran (kme_cddip3_ob_out_pre[72], \kme_cddip3_ob_out_pre.tstrb [0]);
tran (kme_cddip3_ob_out_pre[71], \kme_cddip3_ob_out_pre.tuser [7]);
tran (kme_cddip3_ob_out_pre[70], \kme_cddip3_ob_out_pre.tuser [6]);
tran (kme_cddip3_ob_out_pre[69], \kme_cddip3_ob_out_pre.tuser [5]);
tran (kme_cddip3_ob_out_pre[68], \kme_cddip3_ob_out_pre.tuser [4]);
tran (kme_cddip3_ob_out_pre[67], \kme_cddip3_ob_out_pre.tuser [3]);
tran (kme_cddip3_ob_out_pre[66], \kme_cddip3_ob_out_pre.tuser [2]);
tran (kme_cddip3_ob_out_pre[65], \kme_cddip3_ob_out_pre.tuser [1]);
tran (kme_cddip3_ob_out_pre[64], \kme_cddip3_ob_out_pre.tuser [0]);
tran (kme_cddip3_ob_out_pre[63], \kme_cddip3_ob_out_pre.tdata [63]);
tran (kme_cddip3_ob_out_pre[62], \kme_cddip3_ob_out_pre.tdata [62]);
tran (kme_cddip3_ob_out_pre[61], \kme_cddip3_ob_out_pre.tdata [61]);
tran (kme_cddip3_ob_out_pre[60], \kme_cddip3_ob_out_pre.tdata [60]);
tran (kme_cddip3_ob_out_pre[59], \kme_cddip3_ob_out_pre.tdata [59]);
tran (kme_cddip3_ob_out_pre[58], \kme_cddip3_ob_out_pre.tdata [58]);
tran (kme_cddip3_ob_out_pre[57], \kme_cddip3_ob_out_pre.tdata [57]);
tran (kme_cddip3_ob_out_pre[56], \kme_cddip3_ob_out_pre.tdata [56]);
tran (kme_cddip3_ob_out_pre[55], \kme_cddip3_ob_out_pre.tdata [55]);
tran (kme_cddip3_ob_out_pre[54], \kme_cddip3_ob_out_pre.tdata [54]);
tran (kme_cddip3_ob_out_pre[53], \kme_cddip3_ob_out_pre.tdata [53]);
tran (kme_cddip3_ob_out_pre[52], \kme_cddip3_ob_out_pre.tdata [52]);
tran (kme_cddip3_ob_out_pre[51], \kme_cddip3_ob_out_pre.tdata [51]);
tran (kme_cddip3_ob_out_pre[50], \kme_cddip3_ob_out_pre.tdata [50]);
tran (kme_cddip3_ob_out_pre[49], \kme_cddip3_ob_out_pre.tdata [49]);
tran (kme_cddip3_ob_out_pre[48], \kme_cddip3_ob_out_pre.tdata [48]);
tran (kme_cddip3_ob_out_pre[47], \kme_cddip3_ob_out_pre.tdata [47]);
tran (kme_cddip3_ob_out_pre[46], \kme_cddip3_ob_out_pre.tdata [46]);
tran (kme_cddip3_ob_out_pre[45], \kme_cddip3_ob_out_pre.tdata [45]);
tran (kme_cddip3_ob_out_pre[44], \kme_cddip3_ob_out_pre.tdata [44]);
tran (kme_cddip3_ob_out_pre[43], \kme_cddip3_ob_out_pre.tdata [43]);
tran (kme_cddip3_ob_out_pre[42], \kme_cddip3_ob_out_pre.tdata [42]);
tran (kme_cddip3_ob_out_pre[41], \kme_cddip3_ob_out_pre.tdata [41]);
tran (kme_cddip3_ob_out_pre[40], \kme_cddip3_ob_out_pre.tdata [40]);
tran (kme_cddip3_ob_out_pre[39], \kme_cddip3_ob_out_pre.tdata [39]);
tran (kme_cddip3_ob_out_pre[38], \kme_cddip3_ob_out_pre.tdata [38]);
tran (kme_cddip3_ob_out_pre[37], \kme_cddip3_ob_out_pre.tdata [37]);
tran (kme_cddip3_ob_out_pre[36], \kme_cddip3_ob_out_pre.tdata [36]);
tran (kme_cddip3_ob_out_pre[35], \kme_cddip3_ob_out_pre.tdata [35]);
tran (kme_cddip3_ob_out_pre[34], \kme_cddip3_ob_out_pre.tdata [34]);
tran (kme_cddip3_ob_out_pre[33], \kme_cddip3_ob_out_pre.tdata [33]);
tran (kme_cddip3_ob_out_pre[32], \kme_cddip3_ob_out_pre.tdata [32]);
tran (kme_cddip3_ob_out_pre[31], \kme_cddip3_ob_out_pre.tdata [31]);
tran (kme_cddip3_ob_out_pre[30], \kme_cddip3_ob_out_pre.tdata [30]);
tran (kme_cddip3_ob_out_pre[29], \kme_cddip3_ob_out_pre.tdata [29]);
tran (kme_cddip3_ob_out_pre[28], \kme_cddip3_ob_out_pre.tdata [28]);
tran (kme_cddip3_ob_out_pre[27], \kme_cddip3_ob_out_pre.tdata [27]);
tran (kme_cddip3_ob_out_pre[26], \kme_cddip3_ob_out_pre.tdata [26]);
tran (kme_cddip3_ob_out_pre[25], \kme_cddip3_ob_out_pre.tdata [25]);
tran (kme_cddip3_ob_out_pre[24], \kme_cddip3_ob_out_pre.tdata [24]);
tran (kme_cddip3_ob_out_pre[23], \kme_cddip3_ob_out_pre.tdata [23]);
tran (kme_cddip3_ob_out_pre[22], \kme_cddip3_ob_out_pre.tdata [22]);
tran (kme_cddip3_ob_out_pre[21], \kme_cddip3_ob_out_pre.tdata [21]);
tran (kme_cddip3_ob_out_pre[20], \kme_cddip3_ob_out_pre.tdata [20]);
tran (kme_cddip3_ob_out_pre[19], \kme_cddip3_ob_out_pre.tdata [19]);
tran (kme_cddip3_ob_out_pre[18], \kme_cddip3_ob_out_pre.tdata [18]);
tran (kme_cddip3_ob_out_pre[17], \kme_cddip3_ob_out_pre.tdata [17]);
tran (kme_cddip3_ob_out_pre[16], \kme_cddip3_ob_out_pre.tdata [16]);
tran (kme_cddip3_ob_out_pre[15], \kme_cddip3_ob_out_pre.tdata [15]);
tran (kme_cddip3_ob_out_pre[14], \kme_cddip3_ob_out_pre.tdata [14]);
tran (kme_cddip3_ob_out_pre[13], \kme_cddip3_ob_out_pre.tdata [13]);
tran (kme_cddip3_ob_out_pre[12], \kme_cddip3_ob_out_pre.tdata [12]);
tran (kme_cddip3_ob_out_pre[11], \kme_cddip3_ob_out_pre.tdata [11]);
tran (kme_cddip3_ob_out_pre[10], \kme_cddip3_ob_out_pre.tdata [10]);
tran (kme_cddip3_ob_out_pre[9], \kme_cddip3_ob_out_pre.tdata [9]);
tran (kme_cddip3_ob_out_pre[8], \kme_cddip3_ob_out_pre.tdata [8]);
tran (kme_cddip3_ob_out_pre[7], \kme_cddip3_ob_out_pre.tdata [7]);
tran (kme_cddip3_ob_out_pre[6], \kme_cddip3_ob_out_pre.tdata [6]);
tran (kme_cddip3_ob_out_pre[5], \kme_cddip3_ob_out_pre.tdata [5]);
tran (kme_cddip3_ob_out_pre[4], \kme_cddip3_ob_out_pre.tdata [4]);
tran (kme_cddip3_ob_out_pre[3], \kme_cddip3_ob_out_pre.tdata [3]);
tran (kme_cddip3_ob_out_pre[2], \kme_cddip3_ob_out_pre.tdata [2]);
tran (kme_cddip3_ob_out_pre[1], \kme_cddip3_ob_out_pre.tdata [1]);
tran (kme_cddip3_ob_out_pre[0], \kme_cddip3_ob_out_pre.tdata [0]);
tran (idle_components[31], \idle_components.r.part0 [31]);
tran (idle_components[31], \idle_components.f.num_key_tlvs_in_flight [19]);
tran (idle_components[30], \idle_components.r.part0 [30]);
tran (idle_components[30], \idle_components.f.num_key_tlvs_in_flight [18]);
tran (idle_components[29], \idle_components.r.part0 [29]);
tran (idle_components[29], \idle_components.f.num_key_tlvs_in_flight [17]);
tran (idle_components[28], \idle_components.r.part0 [28]);
tran (idle_components[28], \idle_components.f.num_key_tlvs_in_flight [16]);
tran (idle_components[27], \idle_components.r.part0 [27]);
tran (idle_components[27], \idle_components.f.num_key_tlvs_in_flight [15]);
tran (idle_components[26], \idle_components.r.part0 [26]);
tran (idle_components[26], \idle_components.f.num_key_tlvs_in_flight [14]);
tran (idle_components[25], \idle_components.r.part0 [25]);
tran (idle_components[25], \idle_components.f.num_key_tlvs_in_flight [13]);
tran (idle_components[24], \idle_components.r.part0 [24]);
tran (idle_components[24], \idle_components.f.num_key_tlvs_in_flight [12]);
tran (idle_components[23], \idle_components.r.part0 [23]);
tran (idle_components[23], \idle_components.f.num_key_tlvs_in_flight [11]);
tran (idle_components[22], \idle_components.r.part0 [22]);
tran (idle_components[22], \idle_components.f.num_key_tlvs_in_flight [10]);
tran (idle_components[21], \idle_components.r.part0 [21]);
tran (idle_components[21], \idle_components.f.num_key_tlvs_in_flight [9]);
tran (idle_components[20], \idle_components.r.part0 [20]);
tran (idle_components[20], \idle_components.f.num_key_tlvs_in_flight [8]);
tran (idle_components[19], \idle_components.r.part0 [19]);
tran (idle_components[19], \idle_components.f.num_key_tlvs_in_flight [7]);
tran (idle_components[18], \idle_components.r.part0 [18]);
tran (idle_components[18], \idle_components.f.num_key_tlvs_in_flight [6]);
tran (idle_components[17], \idle_components.r.part0 [17]);
tran (idle_components[17], \idle_components.f.num_key_tlvs_in_flight [5]);
tran (idle_components[16], \idle_components.r.part0 [16]);
tran (idle_components[16], \idle_components.f.num_key_tlvs_in_flight [4]);
tran (idle_components[15], \idle_components.r.part0 [15]);
tran (idle_components[15], \idle_components.f.num_key_tlvs_in_flight [3]);
tran (idle_components[14], \idle_components.r.part0 [14]);
tran (idle_components[14], \idle_components.f.num_key_tlvs_in_flight [2]);
tran (idle_components[13], \idle_components.r.part0 [13]);
tran (idle_components[13], \idle_components.f.num_key_tlvs_in_flight [1]);
tran (idle_components[12], \idle_components.r.part0 [12]);
tran (idle_components[12], \idle_components.f.num_key_tlvs_in_flight [0]);
tran (idle_components[11], \idle_components.r.part0 [11]);
tran (idle_components[11], \idle_components.f.cddip0_key_tlv_rsm_idle );
tran (idle_components[10], \idle_components.r.part0 [10]);
tran (idle_components[10], \idle_components.f.cddip1_key_tlv_rsm_idle );
tran (idle_components[9], \idle_components.r.part0 [9]);
tran (idle_components[9], \idle_components.f.cddip2_key_tlv_rsm_idle );
tran (idle_components[8], \idle_components.r.part0 [8]);
tran (idle_components[8], \idle_components.f.cddip3_key_tlv_rsm_idle );
tran (idle_components[7], \idle_components.r.part0 [7]);
tran (idle_components[7], \idle_components.f.cceip0_key_tlv_rsm_idle );
tran (idle_components[6], \idle_components.r.part0 [6]);
tran (idle_components[6], \idle_components.f.cceip1_key_tlv_rsm_idle );
tran (idle_components[5], \idle_components.r.part0 [5]);
tran (idle_components[5], \idle_components.f.cceip2_key_tlv_rsm_idle );
tran (idle_components[4], \idle_components.r.part0 [4]);
tran (idle_components[4], \idle_components.f.cceip3_key_tlv_rsm_idle );
tran (idle_components[3], \idle_components.r.part0 [3]);
tran (idle_components[3], \idle_components.f.no_key_tlv_in_flight );
tran (idle_components[2], \idle_components.r.part0 [2]);
tran (idle_components[2], \idle_components.f.tlv_parser_idle );
tran (idle_components[1], \idle_components.r.part0 [1]);
tran (idle_components[1], \idle_components.f.drng_idle );
tran (idle_components[0], \idle_components.r.part0 [0]);
tran (idle_components[0], \idle_components.f.kme_slv_empty );
tran (\_zy_simnet_tvar_20[7][271] , \_zy_simnet_tvar_20[7].guid_size[0] );
tran (\_zy_simnet_tvar_20[7][270] , \_zy_simnet_tvar_20[7].label_size[5] );
tran (\_zy_simnet_tvar_20[7][269] , \_zy_simnet_tvar_20[7].label_size[4] );
tran (\_zy_simnet_tvar_20[7][268] , \_zy_simnet_tvar_20[7].label_size[3] );
tran (\_zy_simnet_tvar_20[7][267] , \_zy_simnet_tvar_20[7].label_size[2] );
tran (\_zy_simnet_tvar_20[7][266] , \_zy_simnet_tvar_20[7].label_size[1] );
tran (\_zy_simnet_tvar_20[7][265] , \_zy_simnet_tvar_20[7].label_size[0] );
tran (\_zy_simnet_tvar_20[7][264] , \_zy_simnet_tvar_20[7].label[255] );
tran (\_zy_simnet_tvar_20[7][263] , \_zy_simnet_tvar_20[7].label[254] );
tran (\_zy_simnet_tvar_20[7][262] , \_zy_simnet_tvar_20[7].label[253] );
tran (\_zy_simnet_tvar_20[7][261] , \_zy_simnet_tvar_20[7].label[252] );
tran (\_zy_simnet_tvar_20[7][260] , \_zy_simnet_tvar_20[7].label[251] );
tran (\_zy_simnet_tvar_20[7][259] , \_zy_simnet_tvar_20[7].label[250] );
tran (\_zy_simnet_tvar_20[7][258] , \_zy_simnet_tvar_20[7].label[249] );
tran (\_zy_simnet_tvar_20[7][257] , \_zy_simnet_tvar_20[7].label[248] );
tran (\_zy_simnet_tvar_20[7][256] , \_zy_simnet_tvar_20[7].label[247] );
tran (\_zy_simnet_tvar_20[7][255] , \_zy_simnet_tvar_20[7].label[246] );
tran (\_zy_simnet_tvar_20[7][254] , \_zy_simnet_tvar_20[7].label[245] );
tran (\_zy_simnet_tvar_20[7][253] , \_zy_simnet_tvar_20[7].label[244] );
tran (\_zy_simnet_tvar_20[7][252] , \_zy_simnet_tvar_20[7].label[243] );
tran (\_zy_simnet_tvar_20[7][251] , \_zy_simnet_tvar_20[7].label[242] );
tran (\_zy_simnet_tvar_20[7][250] , \_zy_simnet_tvar_20[7].label[241] );
tran (\_zy_simnet_tvar_20[7][249] , \_zy_simnet_tvar_20[7].label[240] );
tran (\_zy_simnet_tvar_20[7][248] , \_zy_simnet_tvar_20[7].label[239] );
tran (\_zy_simnet_tvar_20[7][247] , \_zy_simnet_tvar_20[7].label[238] );
tran (\_zy_simnet_tvar_20[7][246] , \_zy_simnet_tvar_20[7].label[237] );
tran (\_zy_simnet_tvar_20[7][245] , \_zy_simnet_tvar_20[7].label[236] );
tran (\_zy_simnet_tvar_20[7][244] , \_zy_simnet_tvar_20[7].label[235] );
tran (\_zy_simnet_tvar_20[7][243] , \_zy_simnet_tvar_20[7].label[234] );
tran (\_zy_simnet_tvar_20[7][242] , \_zy_simnet_tvar_20[7].label[233] );
tran (\_zy_simnet_tvar_20[7][241] , \_zy_simnet_tvar_20[7].label[232] );
tran (\_zy_simnet_tvar_20[7][240] , \_zy_simnet_tvar_20[7].label[231] );
tran (\_zy_simnet_tvar_20[7][239] , \_zy_simnet_tvar_20[7].label[230] );
tran (\_zy_simnet_tvar_20[7][238] , \_zy_simnet_tvar_20[7].label[229] );
tran (\_zy_simnet_tvar_20[7][237] , \_zy_simnet_tvar_20[7].label[228] );
tran (\_zy_simnet_tvar_20[7][236] , \_zy_simnet_tvar_20[7].label[227] );
tran (\_zy_simnet_tvar_20[7][235] , \_zy_simnet_tvar_20[7].label[226] );
tran (\_zy_simnet_tvar_20[7][234] , \_zy_simnet_tvar_20[7].label[225] );
tran (\_zy_simnet_tvar_20[7][233] , \_zy_simnet_tvar_20[7].label[224] );
tran (\_zy_simnet_tvar_20[7][232] , \_zy_simnet_tvar_20[7].label[223] );
tran (\_zy_simnet_tvar_20[7][231] , \_zy_simnet_tvar_20[7].label[222] );
tran (\_zy_simnet_tvar_20[7][230] , \_zy_simnet_tvar_20[7].label[221] );
tran (\_zy_simnet_tvar_20[7][229] , \_zy_simnet_tvar_20[7].label[220] );
tran (\_zy_simnet_tvar_20[7][228] , \_zy_simnet_tvar_20[7].label[219] );
tran (\_zy_simnet_tvar_20[7][227] , \_zy_simnet_tvar_20[7].label[218] );
tran (\_zy_simnet_tvar_20[7][226] , \_zy_simnet_tvar_20[7].label[217] );
tran (\_zy_simnet_tvar_20[7][225] , \_zy_simnet_tvar_20[7].label[216] );
tran (\_zy_simnet_tvar_20[7][224] , \_zy_simnet_tvar_20[7].label[215] );
tran (\_zy_simnet_tvar_20[7][223] , \_zy_simnet_tvar_20[7].label[214] );
tran (\_zy_simnet_tvar_20[7][222] , \_zy_simnet_tvar_20[7].label[213] );
tran (\_zy_simnet_tvar_20[7][221] , \_zy_simnet_tvar_20[7].label[212] );
tran (\_zy_simnet_tvar_20[7][220] , \_zy_simnet_tvar_20[7].label[211] );
tran (\_zy_simnet_tvar_20[7][219] , \_zy_simnet_tvar_20[7].label[210] );
tran (\_zy_simnet_tvar_20[7][218] , \_zy_simnet_tvar_20[7].label[209] );
tran (\_zy_simnet_tvar_20[7][217] , \_zy_simnet_tvar_20[7].label[208] );
tran (\_zy_simnet_tvar_20[7][216] , \_zy_simnet_tvar_20[7].label[207] );
tran (\_zy_simnet_tvar_20[7][215] , \_zy_simnet_tvar_20[7].label[206] );
tran (\_zy_simnet_tvar_20[7][214] , \_zy_simnet_tvar_20[7].label[205] );
tran (\_zy_simnet_tvar_20[7][213] , \_zy_simnet_tvar_20[7].label[204] );
tran (\_zy_simnet_tvar_20[7][212] , \_zy_simnet_tvar_20[7].label[203] );
tran (\_zy_simnet_tvar_20[7][211] , \_zy_simnet_tvar_20[7].label[202] );
tran (\_zy_simnet_tvar_20[7][210] , \_zy_simnet_tvar_20[7].label[201] );
tran (\_zy_simnet_tvar_20[7][209] , \_zy_simnet_tvar_20[7].label[200] );
tran (\_zy_simnet_tvar_20[7][208] , \_zy_simnet_tvar_20[7].label[199] );
tran (\_zy_simnet_tvar_20[7][207] , \_zy_simnet_tvar_20[7].label[198] );
tran (\_zy_simnet_tvar_20[7][206] , \_zy_simnet_tvar_20[7].label[197] );
tran (\_zy_simnet_tvar_20[7][205] , \_zy_simnet_tvar_20[7].label[196] );
tran (\_zy_simnet_tvar_20[7][204] , \_zy_simnet_tvar_20[7].label[195] );
tran (\_zy_simnet_tvar_20[7][203] , \_zy_simnet_tvar_20[7].label[194] );
tran (\_zy_simnet_tvar_20[7][202] , \_zy_simnet_tvar_20[7].label[193] );
tran (\_zy_simnet_tvar_20[7][201] , \_zy_simnet_tvar_20[7].label[192] );
tran (\_zy_simnet_tvar_20[7][200] , \_zy_simnet_tvar_20[7].label[191] );
tran (\_zy_simnet_tvar_20[7][199] , \_zy_simnet_tvar_20[7].label[190] );
tran (\_zy_simnet_tvar_20[7][198] , \_zy_simnet_tvar_20[7].label[189] );
tran (\_zy_simnet_tvar_20[7][197] , \_zy_simnet_tvar_20[7].label[188] );
tran (\_zy_simnet_tvar_20[7][196] , \_zy_simnet_tvar_20[7].label[187] );
tran (\_zy_simnet_tvar_20[7][195] , \_zy_simnet_tvar_20[7].label[186] );
tran (\_zy_simnet_tvar_20[7][194] , \_zy_simnet_tvar_20[7].label[185] );
tran (\_zy_simnet_tvar_20[7][193] , \_zy_simnet_tvar_20[7].label[184] );
tran (\_zy_simnet_tvar_20[7][192] , \_zy_simnet_tvar_20[7].label[183] );
tran (\_zy_simnet_tvar_20[7][191] , \_zy_simnet_tvar_20[7].label[182] );
tran (\_zy_simnet_tvar_20[7][190] , \_zy_simnet_tvar_20[7].label[181] );
tran (\_zy_simnet_tvar_20[7][189] , \_zy_simnet_tvar_20[7].label[180] );
tran (\_zy_simnet_tvar_20[7][188] , \_zy_simnet_tvar_20[7].label[179] );
tran (\_zy_simnet_tvar_20[7][187] , \_zy_simnet_tvar_20[7].label[178] );
tran (\_zy_simnet_tvar_20[7][186] , \_zy_simnet_tvar_20[7].label[177] );
tran (\_zy_simnet_tvar_20[7][185] , \_zy_simnet_tvar_20[7].label[176] );
tran (\_zy_simnet_tvar_20[7][184] , \_zy_simnet_tvar_20[7].label[175] );
tran (\_zy_simnet_tvar_20[7][183] , \_zy_simnet_tvar_20[7].label[174] );
tran (\_zy_simnet_tvar_20[7][182] , \_zy_simnet_tvar_20[7].label[173] );
tran (\_zy_simnet_tvar_20[7][181] , \_zy_simnet_tvar_20[7].label[172] );
tran (\_zy_simnet_tvar_20[7][180] , \_zy_simnet_tvar_20[7].label[171] );
tran (\_zy_simnet_tvar_20[7][179] , \_zy_simnet_tvar_20[7].label[170] );
tran (\_zy_simnet_tvar_20[7][178] , \_zy_simnet_tvar_20[7].label[169] );
tran (\_zy_simnet_tvar_20[7][177] , \_zy_simnet_tvar_20[7].label[168] );
tran (\_zy_simnet_tvar_20[7][176] , \_zy_simnet_tvar_20[7].label[167] );
tran (\_zy_simnet_tvar_20[7][175] , \_zy_simnet_tvar_20[7].label[166] );
tran (\_zy_simnet_tvar_20[7][174] , \_zy_simnet_tvar_20[7].label[165] );
tran (\_zy_simnet_tvar_20[7][173] , \_zy_simnet_tvar_20[7].label[164] );
tran (\_zy_simnet_tvar_20[7][172] , \_zy_simnet_tvar_20[7].label[163] );
tran (\_zy_simnet_tvar_20[7][171] , \_zy_simnet_tvar_20[7].label[162] );
tran (\_zy_simnet_tvar_20[7][170] , \_zy_simnet_tvar_20[7].label[161] );
tran (\_zy_simnet_tvar_20[7][169] , \_zy_simnet_tvar_20[7].label[160] );
tran (\_zy_simnet_tvar_20[7][168] , \_zy_simnet_tvar_20[7].label[159] );
tran (\_zy_simnet_tvar_20[7][167] , \_zy_simnet_tvar_20[7].label[158] );
tran (\_zy_simnet_tvar_20[7][166] , \_zy_simnet_tvar_20[7].label[157] );
tran (\_zy_simnet_tvar_20[7][165] , \_zy_simnet_tvar_20[7].label[156] );
tran (\_zy_simnet_tvar_20[7][164] , \_zy_simnet_tvar_20[7].label[155] );
tran (\_zy_simnet_tvar_20[7][163] , \_zy_simnet_tvar_20[7].label[154] );
tran (\_zy_simnet_tvar_20[7][162] , \_zy_simnet_tvar_20[7].label[153] );
tran (\_zy_simnet_tvar_20[7][161] , \_zy_simnet_tvar_20[7].label[152] );
tran (\_zy_simnet_tvar_20[7][160] , \_zy_simnet_tvar_20[7].label[151] );
tran (\_zy_simnet_tvar_20[7][159] , \_zy_simnet_tvar_20[7].label[150] );
tran (\_zy_simnet_tvar_20[7][158] , \_zy_simnet_tvar_20[7].label[149] );
tran (\_zy_simnet_tvar_20[7][157] , \_zy_simnet_tvar_20[7].label[148] );
tran (\_zy_simnet_tvar_20[7][156] , \_zy_simnet_tvar_20[7].label[147] );
tran (\_zy_simnet_tvar_20[7][155] , \_zy_simnet_tvar_20[7].label[146] );
tran (\_zy_simnet_tvar_20[7][154] , \_zy_simnet_tvar_20[7].label[145] );
tran (\_zy_simnet_tvar_20[7][153] , \_zy_simnet_tvar_20[7].label[144] );
tran (\_zy_simnet_tvar_20[7][152] , \_zy_simnet_tvar_20[7].label[143] );
tran (\_zy_simnet_tvar_20[7][151] , \_zy_simnet_tvar_20[7].label[142] );
tran (\_zy_simnet_tvar_20[7][150] , \_zy_simnet_tvar_20[7].label[141] );
tran (\_zy_simnet_tvar_20[7][149] , \_zy_simnet_tvar_20[7].label[140] );
tran (\_zy_simnet_tvar_20[7][148] , \_zy_simnet_tvar_20[7].label[139] );
tran (\_zy_simnet_tvar_20[7][147] , \_zy_simnet_tvar_20[7].label[138] );
tran (\_zy_simnet_tvar_20[7][146] , \_zy_simnet_tvar_20[7].label[137] );
tran (\_zy_simnet_tvar_20[7][145] , \_zy_simnet_tvar_20[7].label[136] );
tran (\_zy_simnet_tvar_20[7][144] , \_zy_simnet_tvar_20[7].label[135] );
tran (\_zy_simnet_tvar_20[7][143] , \_zy_simnet_tvar_20[7].label[134] );
tran (\_zy_simnet_tvar_20[7][142] , \_zy_simnet_tvar_20[7].label[133] );
tran (\_zy_simnet_tvar_20[7][141] , \_zy_simnet_tvar_20[7].label[132] );
tran (\_zy_simnet_tvar_20[7][140] , \_zy_simnet_tvar_20[7].label[131] );
tran (\_zy_simnet_tvar_20[7][139] , \_zy_simnet_tvar_20[7].label[130] );
tran (\_zy_simnet_tvar_20[7][138] , \_zy_simnet_tvar_20[7].label[129] );
tran (\_zy_simnet_tvar_20[7][137] , \_zy_simnet_tvar_20[7].label[128] );
tran (\_zy_simnet_tvar_20[7][136] , \_zy_simnet_tvar_20[7].label[127] );
tran (\_zy_simnet_tvar_20[7][135] , \_zy_simnet_tvar_20[7].label[126] );
tran (\_zy_simnet_tvar_20[7][134] , \_zy_simnet_tvar_20[7].label[125] );
tran (\_zy_simnet_tvar_20[7][133] , \_zy_simnet_tvar_20[7].label[124] );
tran (\_zy_simnet_tvar_20[7][132] , \_zy_simnet_tvar_20[7].label[123] );
tran (\_zy_simnet_tvar_20[7][131] , \_zy_simnet_tvar_20[7].label[122] );
tran (\_zy_simnet_tvar_20[7][130] , \_zy_simnet_tvar_20[7].label[121] );
tran (\_zy_simnet_tvar_20[7][129] , \_zy_simnet_tvar_20[7].label[120] );
tran (\_zy_simnet_tvar_20[7][128] , \_zy_simnet_tvar_20[7].label[119] );
tran (\_zy_simnet_tvar_20[7][127] , \_zy_simnet_tvar_20[7].label[118] );
tran (\_zy_simnet_tvar_20[7][126] , \_zy_simnet_tvar_20[7].label[117] );
tran (\_zy_simnet_tvar_20[7][125] , \_zy_simnet_tvar_20[7].label[116] );
tran (\_zy_simnet_tvar_20[7][124] , \_zy_simnet_tvar_20[7].label[115] );
tran (\_zy_simnet_tvar_20[7][123] , \_zy_simnet_tvar_20[7].label[114] );
tran (\_zy_simnet_tvar_20[7][122] , \_zy_simnet_tvar_20[7].label[113] );
tran (\_zy_simnet_tvar_20[7][121] , \_zy_simnet_tvar_20[7].label[112] );
tran (\_zy_simnet_tvar_20[7][120] , \_zy_simnet_tvar_20[7].label[111] );
tran (\_zy_simnet_tvar_20[7][119] , \_zy_simnet_tvar_20[7].label[110] );
tran (\_zy_simnet_tvar_20[7][118] , \_zy_simnet_tvar_20[7].label[109] );
tran (\_zy_simnet_tvar_20[7][117] , \_zy_simnet_tvar_20[7].label[108] );
tran (\_zy_simnet_tvar_20[7][116] , \_zy_simnet_tvar_20[7].label[107] );
tran (\_zy_simnet_tvar_20[7][115] , \_zy_simnet_tvar_20[7].label[106] );
tran (\_zy_simnet_tvar_20[7][114] , \_zy_simnet_tvar_20[7].label[105] );
tran (\_zy_simnet_tvar_20[7][113] , \_zy_simnet_tvar_20[7].label[104] );
tran (\_zy_simnet_tvar_20[7][112] , \_zy_simnet_tvar_20[7].label[103] );
tran (\_zy_simnet_tvar_20[7][111] , \_zy_simnet_tvar_20[7].label[102] );
tran (\_zy_simnet_tvar_20[7][110] , \_zy_simnet_tvar_20[7].label[101] );
tran (\_zy_simnet_tvar_20[7][109] , \_zy_simnet_tvar_20[7].label[100] );
tran (\_zy_simnet_tvar_20[7][108] , \_zy_simnet_tvar_20[7].label[99] );
tran (\_zy_simnet_tvar_20[7][107] , \_zy_simnet_tvar_20[7].label[98] );
tran (\_zy_simnet_tvar_20[7][106] , \_zy_simnet_tvar_20[7].label[97] );
tran (\_zy_simnet_tvar_20[7][105] , \_zy_simnet_tvar_20[7].label[96] );
tran (\_zy_simnet_tvar_20[7][104] , \_zy_simnet_tvar_20[7].label[95] );
tran (\_zy_simnet_tvar_20[7][103] , \_zy_simnet_tvar_20[7].label[94] );
tran (\_zy_simnet_tvar_20[7][102] , \_zy_simnet_tvar_20[7].label[93] );
tran (\_zy_simnet_tvar_20[7][101] , \_zy_simnet_tvar_20[7].label[92] );
tran (\_zy_simnet_tvar_20[7][100] , \_zy_simnet_tvar_20[7].label[91] );
tran (\_zy_simnet_tvar_20[7][99] , \_zy_simnet_tvar_20[7].label[90] );
tran (\_zy_simnet_tvar_20[7][98] , \_zy_simnet_tvar_20[7].label[89] );
tran (\_zy_simnet_tvar_20[7][97] , \_zy_simnet_tvar_20[7].label[88] );
tran (\_zy_simnet_tvar_20[7][96] , \_zy_simnet_tvar_20[7].label[87] );
tran (\_zy_simnet_tvar_20[7][95] , \_zy_simnet_tvar_20[7].label[86] );
tran (\_zy_simnet_tvar_20[7][94] , \_zy_simnet_tvar_20[7].label[85] );
tran (\_zy_simnet_tvar_20[7][93] , \_zy_simnet_tvar_20[7].label[84] );
tran (\_zy_simnet_tvar_20[7][92] , \_zy_simnet_tvar_20[7].label[83] );
tran (\_zy_simnet_tvar_20[7][91] , \_zy_simnet_tvar_20[7].label[82] );
tran (\_zy_simnet_tvar_20[7][90] , \_zy_simnet_tvar_20[7].label[81] );
tran (\_zy_simnet_tvar_20[7][89] , \_zy_simnet_tvar_20[7].label[80] );
tran (\_zy_simnet_tvar_20[7][88] , \_zy_simnet_tvar_20[7].label[79] );
tran (\_zy_simnet_tvar_20[7][87] , \_zy_simnet_tvar_20[7].label[78] );
tran (\_zy_simnet_tvar_20[7][86] , \_zy_simnet_tvar_20[7].label[77] );
tran (\_zy_simnet_tvar_20[7][85] , \_zy_simnet_tvar_20[7].label[76] );
tran (\_zy_simnet_tvar_20[7][84] , \_zy_simnet_tvar_20[7].label[75] );
tran (\_zy_simnet_tvar_20[7][83] , \_zy_simnet_tvar_20[7].label[74] );
tran (\_zy_simnet_tvar_20[7][82] , \_zy_simnet_tvar_20[7].label[73] );
tran (\_zy_simnet_tvar_20[7][81] , \_zy_simnet_tvar_20[7].label[72] );
tran (\_zy_simnet_tvar_20[7][80] , \_zy_simnet_tvar_20[7].label[71] );
tran (\_zy_simnet_tvar_20[7][79] , \_zy_simnet_tvar_20[7].label[70] );
tran (\_zy_simnet_tvar_20[7][78] , \_zy_simnet_tvar_20[7].label[69] );
tran (\_zy_simnet_tvar_20[7][77] , \_zy_simnet_tvar_20[7].label[68] );
tran (\_zy_simnet_tvar_20[7][76] , \_zy_simnet_tvar_20[7].label[67] );
tran (\_zy_simnet_tvar_20[7][75] , \_zy_simnet_tvar_20[7].label[66] );
tran (\_zy_simnet_tvar_20[7][74] , \_zy_simnet_tvar_20[7].label[65] );
tran (\_zy_simnet_tvar_20[7][73] , \_zy_simnet_tvar_20[7].label[64] );
tran (\_zy_simnet_tvar_20[7][72] , \_zy_simnet_tvar_20[7].label[63] );
tran (\_zy_simnet_tvar_20[7][71] , \_zy_simnet_tvar_20[7].label[62] );
tran (\_zy_simnet_tvar_20[7][70] , \_zy_simnet_tvar_20[7].label[61] );
tran (\_zy_simnet_tvar_20[7][69] , \_zy_simnet_tvar_20[7].label[60] );
tran (\_zy_simnet_tvar_20[7][68] , \_zy_simnet_tvar_20[7].label[59] );
tran (\_zy_simnet_tvar_20[7][67] , \_zy_simnet_tvar_20[7].label[58] );
tran (\_zy_simnet_tvar_20[7][66] , \_zy_simnet_tvar_20[7].label[57] );
tran (\_zy_simnet_tvar_20[7][65] , \_zy_simnet_tvar_20[7].label[56] );
tran (\_zy_simnet_tvar_20[7][64] , \_zy_simnet_tvar_20[7].label[55] );
tran (\_zy_simnet_tvar_20[7][63] , \_zy_simnet_tvar_20[7].label[54] );
tran (\_zy_simnet_tvar_20[7][62] , \_zy_simnet_tvar_20[7].label[53] );
tran (\_zy_simnet_tvar_20[7][61] , \_zy_simnet_tvar_20[7].label[52] );
tran (\_zy_simnet_tvar_20[7][60] , \_zy_simnet_tvar_20[7].label[51] );
tran (\_zy_simnet_tvar_20[7][59] , \_zy_simnet_tvar_20[7].label[50] );
tran (\_zy_simnet_tvar_20[7][58] , \_zy_simnet_tvar_20[7].label[49] );
tran (\_zy_simnet_tvar_20[7][57] , \_zy_simnet_tvar_20[7].label[48] );
tran (\_zy_simnet_tvar_20[7][56] , \_zy_simnet_tvar_20[7].label[47] );
tran (\_zy_simnet_tvar_20[7][55] , \_zy_simnet_tvar_20[7].label[46] );
tran (\_zy_simnet_tvar_20[7][54] , \_zy_simnet_tvar_20[7].label[45] );
tran (\_zy_simnet_tvar_20[7][53] , \_zy_simnet_tvar_20[7].label[44] );
tran (\_zy_simnet_tvar_20[7][52] , \_zy_simnet_tvar_20[7].label[43] );
tran (\_zy_simnet_tvar_20[7][51] , \_zy_simnet_tvar_20[7].label[42] );
tran (\_zy_simnet_tvar_20[7][50] , \_zy_simnet_tvar_20[7].label[41] );
tran (\_zy_simnet_tvar_20[7][49] , \_zy_simnet_tvar_20[7].label[40] );
tran (\_zy_simnet_tvar_20[7][48] , \_zy_simnet_tvar_20[7].label[39] );
tran (\_zy_simnet_tvar_20[7][47] , \_zy_simnet_tvar_20[7].label[38] );
tran (\_zy_simnet_tvar_20[7][46] , \_zy_simnet_tvar_20[7].label[37] );
tran (\_zy_simnet_tvar_20[7][45] , \_zy_simnet_tvar_20[7].label[36] );
tran (\_zy_simnet_tvar_20[7][44] , \_zy_simnet_tvar_20[7].label[35] );
tran (\_zy_simnet_tvar_20[7][43] , \_zy_simnet_tvar_20[7].label[34] );
tran (\_zy_simnet_tvar_20[7][42] , \_zy_simnet_tvar_20[7].label[33] );
tran (\_zy_simnet_tvar_20[7][41] , \_zy_simnet_tvar_20[7].label[32] );
tran (\_zy_simnet_tvar_20[7][40] , \_zy_simnet_tvar_20[7].label[31] );
tran (\_zy_simnet_tvar_20[7][39] , \_zy_simnet_tvar_20[7].label[30] );
tran (\_zy_simnet_tvar_20[7][38] , \_zy_simnet_tvar_20[7].label[29] );
tran (\_zy_simnet_tvar_20[7][37] , \_zy_simnet_tvar_20[7].label[28] );
tran (\_zy_simnet_tvar_20[7][36] , \_zy_simnet_tvar_20[7].label[27] );
tran (\_zy_simnet_tvar_20[7][35] , \_zy_simnet_tvar_20[7].label[26] );
tran (\_zy_simnet_tvar_20[7][34] , \_zy_simnet_tvar_20[7].label[25] );
tran (\_zy_simnet_tvar_20[7][33] , \_zy_simnet_tvar_20[7].label[24] );
tran (\_zy_simnet_tvar_20[7][32] , \_zy_simnet_tvar_20[7].label[23] );
tran (\_zy_simnet_tvar_20[7][31] , \_zy_simnet_tvar_20[7].label[22] );
tran (\_zy_simnet_tvar_20[7][30] , \_zy_simnet_tvar_20[7].label[21] );
tran (\_zy_simnet_tvar_20[7][29] , \_zy_simnet_tvar_20[7].label[20] );
tran (\_zy_simnet_tvar_20[7][28] , \_zy_simnet_tvar_20[7].label[19] );
tran (\_zy_simnet_tvar_20[7][27] , \_zy_simnet_tvar_20[7].label[18] );
tran (\_zy_simnet_tvar_20[7][26] , \_zy_simnet_tvar_20[7].label[17] );
tran (\_zy_simnet_tvar_20[7][25] , \_zy_simnet_tvar_20[7].label[16] );
tran (\_zy_simnet_tvar_20[7][24] , \_zy_simnet_tvar_20[7].label[15] );
tran (\_zy_simnet_tvar_20[7][23] , \_zy_simnet_tvar_20[7].label[14] );
tran (\_zy_simnet_tvar_20[7][22] , \_zy_simnet_tvar_20[7].label[13] );
tran (\_zy_simnet_tvar_20[7][21] , \_zy_simnet_tvar_20[7].label[12] );
tran (\_zy_simnet_tvar_20[7][20] , \_zy_simnet_tvar_20[7].label[11] );
tran (\_zy_simnet_tvar_20[7][19] , \_zy_simnet_tvar_20[7].label[10] );
tran (\_zy_simnet_tvar_20[7][18] , \_zy_simnet_tvar_20[7].label[9] );
tran (\_zy_simnet_tvar_20[7][17] , \_zy_simnet_tvar_20[7].label[8] );
tran (\_zy_simnet_tvar_20[7][16] , \_zy_simnet_tvar_20[7].label[7] );
tran (\_zy_simnet_tvar_20[7][15] , \_zy_simnet_tvar_20[7].label[6] );
tran (\_zy_simnet_tvar_20[7][14] , \_zy_simnet_tvar_20[7].label[5] );
tran (\_zy_simnet_tvar_20[7][13] , \_zy_simnet_tvar_20[7].label[4] );
tran (\_zy_simnet_tvar_20[7][12] , \_zy_simnet_tvar_20[7].label[3] );
tran (\_zy_simnet_tvar_20[7][11] , \_zy_simnet_tvar_20[7].label[2] );
tran (\_zy_simnet_tvar_20[7][10] , \_zy_simnet_tvar_20[7].label[1] );
tran (\_zy_simnet_tvar_20[7][9] , \_zy_simnet_tvar_20[7].label[0] );
tran (\_zy_simnet_tvar_20[7][8] , \_zy_simnet_tvar_20[7].delimiter_valid[0] );
tran (\_zy_simnet_tvar_20[7][7] , \_zy_simnet_tvar_20[7].delimiter[7] );
tran (\_zy_simnet_tvar_20[7][6] , \_zy_simnet_tvar_20[7].delimiter[6] );
tran (\_zy_simnet_tvar_20[7][5] , \_zy_simnet_tvar_20[7].delimiter[5] );
tran (\_zy_simnet_tvar_20[7][4] , \_zy_simnet_tvar_20[7].delimiter[4] );
tran (\_zy_simnet_tvar_20[7][3] , \_zy_simnet_tvar_20[7].delimiter[3] );
tran (\_zy_simnet_tvar_20[7][2] , \_zy_simnet_tvar_20[7].delimiter[2] );
tran (\_zy_simnet_tvar_20[7][1] , \_zy_simnet_tvar_20[7].delimiter[1] );
tran (\_zy_simnet_tvar_20[7][0] , \_zy_simnet_tvar_20[7].delimiter[0] );
tran (\_zy_simnet_tvar_20[6][271] , \_zy_simnet_tvar_20[6].guid_size[0] );
tran (\_zy_simnet_tvar_20[6][270] , \_zy_simnet_tvar_20[6].label_size[5] );
tran (\_zy_simnet_tvar_20[6][269] , \_zy_simnet_tvar_20[6].label_size[4] );
tran (\_zy_simnet_tvar_20[6][268] , \_zy_simnet_tvar_20[6].label_size[3] );
tran (\_zy_simnet_tvar_20[6][267] , \_zy_simnet_tvar_20[6].label_size[2] );
tran (\_zy_simnet_tvar_20[6][266] , \_zy_simnet_tvar_20[6].label_size[1] );
tran (\_zy_simnet_tvar_20[6][265] , \_zy_simnet_tvar_20[6].label_size[0] );
tran (\_zy_simnet_tvar_20[6][264] , \_zy_simnet_tvar_20[6].label[255] );
tran (\_zy_simnet_tvar_20[6][263] , \_zy_simnet_tvar_20[6].label[254] );
tran (\_zy_simnet_tvar_20[6][262] , \_zy_simnet_tvar_20[6].label[253] );
tran (\_zy_simnet_tvar_20[6][261] , \_zy_simnet_tvar_20[6].label[252] );
tran (\_zy_simnet_tvar_20[6][260] , \_zy_simnet_tvar_20[6].label[251] );
tran (\_zy_simnet_tvar_20[6][259] , \_zy_simnet_tvar_20[6].label[250] );
tran (\_zy_simnet_tvar_20[6][258] , \_zy_simnet_tvar_20[6].label[249] );
tran (\_zy_simnet_tvar_20[6][257] , \_zy_simnet_tvar_20[6].label[248] );
tran (\_zy_simnet_tvar_20[6][256] , \_zy_simnet_tvar_20[6].label[247] );
tran (\_zy_simnet_tvar_20[6][255] , \_zy_simnet_tvar_20[6].label[246] );
tran (\_zy_simnet_tvar_20[6][254] , \_zy_simnet_tvar_20[6].label[245] );
tran (\_zy_simnet_tvar_20[6][253] , \_zy_simnet_tvar_20[6].label[244] );
tran (\_zy_simnet_tvar_20[6][252] , \_zy_simnet_tvar_20[6].label[243] );
tran (\_zy_simnet_tvar_20[6][251] , \_zy_simnet_tvar_20[6].label[242] );
tran (\_zy_simnet_tvar_20[6][250] , \_zy_simnet_tvar_20[6].label[241] );
tran (\_zy_simnet_tvar_20[6][249] , \_zy_simnet_tvar_20[6].label[240] );
tran (\_zy_simnet_tvar_20[6][248] , \_zy_simnet_tvar_20[6].label[239] );
tran (\_zy_simnet_tvar_20[6][247] , \_zy_simnet_tvar_20[6].label[238] );
tran (\_zy_simnet_tvar_20[6][246] , \_zy_simnet_tvar_20[6].label[237] );
tran (\_zy_simnet_tvar_20[6][245] , \_zy_simnet_tvar_20[6].label[236] );
tran (\_zy_simnet_tvar_20[6][244] , \_zy_simnet_tvar_20[6].label[235] );
tran (\_zy_simnet_tvar_20[6][243] , \_zy_simnet_tvar_20[6].label[234] );
tran (\_zy_simnet_tvar_20[6][242] , \_zy_simnet_tvar_20[6].label[233] );
tran (\_zy_simnet_tvar_20[6][241] , \_zy_simnet_tvar_20[6].label[232] );
tran (\_zy_simnet_tvar_20[6][240] , \_zy_simnet_tvar_20[6].label[231] );
tran (\_zy_simnet_tvar_20[6][239] , \_zy_simnet_tvar_20[6].label[230] );
tran (\_zy_simnet_tvar_20[6][238] , \_zy_simnet_tvar_20[6].label[229] );
tran (\_zy_simnet_tvar_20[6][237] , \_zy_simnet_tvar_20[6].label[228] );
tran (\_zy_simnet_tvar_20[6][236] , \_zy_simnet_tvar_20[6].label[227] );
tran (\_zy_simnet_tvar_20[6][235] , \_zy_simnet_tvar_20[6].label[226] );
tran (\_zy_simnet_tvar_20[6][234] , \_zy_simnet_tvar_20[6].label[225] );
tran (\_zy_simnet_tvar_20[6][233] , \_zy_simnet_tvar_20[6].label[224] );
tran (\_zy_simnet_tvar_20[6][232] , \_zy_simnet_tvar_20[6].label[223] );
tran (\_zy_simnet_tvar_20[6][231] , \_zy_simnet_tvar_20[6].label[222] );
tran (\_zy_simnet_tvar_20[6][230] , \_zy_simnet_tvar_20[6].label[221] );
tran (\_zy_simnet_tvar_20[6][229] , \_zy_simnet_tvar_20[6].label[220] );
tran (\_zy_simnet_tvar_20[6][228] , \_zy_simnet_tvar_20[6].label[219] );
tran (\_zy_simnet_tvar_20[6][227] , \_zy_simnet_tvar_20[6].label[218] );
tran (\_zy_simnet_tvar_20[6][226] , \_zy_simnet_tvar_20[6].label[217] );
tran (\_zy_simnet_tvar_20[6][225] , \_zy_simnet_tvar_20[6].label[216] );
tran (\_zy_simnet_tvar_20[6][224] , \_zy_simnet_tvar_20[6].label[215] );
tran (\_zy_simnet_tvar_20[6][223] , \_zy_simnet_tvar_20[6].label[214] );
tran (\_zy_simnet_tvar_20[6][222] , \_zy_simnet_tvar_20[6].label[213] );
tran (\_zy_simnet_tvar_20[6][221] , \_zy_simnet_tvar_20[6].label[212] );
tran (\_zy_simnet_tvar_20[6][220] , \_zy_simnet_tvar_20[6].label[211] );
tran (\_zy_simnet_tvar_20[6][219] , \_zy_simnet_tvar_20[6].label[210] );
tran (\_zy_simnet_tvar_20[6][218] , \_zy_simnet_tvar_20[6].label[209] );
tran (\_zy_simnet_tvar_20[6][217] , \_zy_simnet_tvar_20[6].label[208] );
tran (\_zy_simnet_tvar_20[6][216] , \_zy_simnet_tvar_20[6].label[207] );
tran (\_zy_simnet_tvar_20[6][215] , \_zy_simnet_tvar_20[6].label[206] );
tran (\_zy_simnet_tvar_20[6][214] , \_zy_simnet_tvar_20[6].label[205] );
tran (\_zy_simnet_tvar_20[6][213] , \_zy_simnet_tvar_20[6].label[204] );
tran (\_zy_simnet_tvar_20[6][212] , \_zy_simnet_tvar_20[6].label[203] );
tran (\_zy_simnet_tvar_20[6][211] , \_zy_simnet_tvar_20[6].label[202] );
tran (\_zy_simnet_tvar_20[6][210] , \_zy_simnet_tvar_20[6].label[201] );
tran (\_zy_simnet_tvar_20[6][209] , \_zy_simnet_tvar_20[6].label[200] );
tran (\_zy_simnet_tvar_20[6][208] , \_zy_simnet_tvar_20[6].label[199] );
tran (\_zy_simnet_tvar_20[6][207] , \_zy_simnet_tvar_20[6].label[198] );
tran (\_zy_simnet_tvar_20[6][206] , \_zy_simnet_tvar_20[6].label[197] );
tran (\_zy_simnet_tvar_20[6][205] , \_zy_simnet_tvar_20[6].label[196] );
tran (\_zy_simnet_tvar_20[6][204] , \_zy_simnet_tvar_20[6].label[195] );
tran (\_zy_simnet_tvar_20[6][203] , \_zy_simnet_tvar_20[6].label[194] );
tran (\_zy_simnet_tvar_20[6][202] , \_zy_simnet_tvar_20[6].label[193] );
tran (\_zy_simnet_tvar_20[6][201] , \_zy_simnet_tvar_20[6].label[192] );
tran (\_zy_simnet_tvar_20[6][200] , \_zy_simnet_tvar_20[6].label[191] );
tran (\_zy_simnet_tvar_20[6][199] , \_zy_simnet_tvar_20[6].label[190] );
tran (\_zy_simnet_tvar_20[6][198] , \_zy_simnet_tvar_20[6].label[189] );
tran (\_zy_simnet_tvar_20[6][197] , \_zy_simnet_tvar_20[6].label[188] );
tran (\_zy_simnet_tvar_20[6][196] , \_zy_simnet_tvar_20[6].label[187] );
tran (\_zy_simnet_tvar_20[6][195] , \_zy_simnet_tvar_20[6].label[186] );
tran (\_zy_simnet_tvar_20[6][194] , \_zy_simnet_tvar_20[6].label[185] );
tran (\_zy_simnet_tvar_20[6][193] , \_zy_simnet_tvar_20[6].label[184] );
tran (\_zy_simnet_tvar_20[6][192] , \_zy_simnet_tvar_20[6].label[183] );
tran (\_zy_simnet_tvar_20[6][191] , \_zy_simnet_tvar_20[6].label[182] );
tran (\_zy_simnet_tvar_20[6][190] , \_zy_simnet_tvar_20[6].label[181] );
tran (\_zy_simnet_tvar_20[6][189] , \_zy_simnet_tvar_20[6].label[180] );
tran (\_zy_simnet_tvar_20[6][188] , \_zy_simnet_tvar_20[6].label[179] );
tran (\_zy_simnet_tvar_20[6][187] , \_zy_simnet_tvar_20[6].label[178] );
tran (\_zy_simnet_tvar_20[6][186] , \_zy_simnet_tvar_20[6].label[177] );
tran (\_zy_simnet_tvar_20[6][185] , \_zy_simnet_tvar_20[6].label[176] );
tran (\_zy_simnet_tvar_20[6][184] , \_zy_simnet_tvar_20[6].label[175] );
tran (\_zy_simnet_tvar_20[6][183] , \_zy_simnet_tvar_20[6].label[174] );
tran (\_zy_simnet_tvar_20[6][182] , \_zy_simnet_tvar_20[6].label[173] );
tran (\_zy_simnet_tvar_20[6][181] , \_zy_simnet_tvar_20[6].label[172] );
tran (\_zy_simnet_tvar_20[6][180] , \_zy_simnet_tvar_20[6].label[171] );
tran (\_zy_simnet_tvar_20[6][179] , \_zy_simnet_tvar_20[6].label[170] );
tran (\_zy_simnet_tvar_20[6][178] , \_zy_simnet_tvar_20[6].label[169] );
tran (\_zy_simnet_tvar_20[6][177] , \_zy_simnet_tvar_20[6].label[168] );
tran (\_zy_simnet_tvar_20[6][176] , \_zy_simnet_tvar_20[6].label[167] );
tran (\_zy_simnet_tvar_20[6][175] , \_zy_simnet_tvar_20[6].label[166] );
tran (\_zy_simnet_tvar_20[6][174] , \_zy_simnet_tvar_20[6].label[165] );
tran (\_zy_simnet_tvar_20[6][173] , \_zy_simnet_tvar_20[6].label[164] );
tran (\_zy_simnet_tvar_20[6][172] , \_zy_simnet_tvar_20[6].label[163] );
tran (\_zy_simnet_tvar_20[6][171] , \_zy_simnet_tvar_20[6].label[162] );
tran (\_zy_simnet_tvar_20[6][170] , \_zy_simnet_tvar_20[6].label[161] );
tran (\_zy_simnet_tvar_20[6][169] , \_zy_simnet_tvar_20[6].label[160] );
tran (\_zy_simnet_tvar_20[6][168] , \_zy_simnet_tvar_20[6].label[159] );
tran (\_zy_simnet_tvar_20[6][167] , \_zy_simnet_tvar_20[6].label[158] );
tran (\_zy_simnet_tvar_20[6][166] , \_zy_simnet_tvar_20[6].label[157] );
tran (\_zy_simnet_tvar_20[6][165] , \_zy_simnet_tvar_20[6].label[156] );
tran (\_zy_simnet_tvar_20[6][164] , \_zy_simnet_tvar_20[6].label[155] );
tran (\_zy_simnet_tvar_20[6][163] , \_zy_simnet_tvar_20[6].label[154] );
tran (\_zy_simnet_tvar_20[6][162] , \_zy_simnet_tvar_20[6].label[153] );
tran (\_zy_simnet_tvar_20[6][161] , \_zy_simnet_tvar_20[6].label[152] );
tran (\_zy_simnet_tvar_20[6][160] , \_zy_simnet_tvar_20[6].label[151] );
tran (\_zy_simnet_tvar_20[6][159] , \_zy_simnet_tvar_20[6].label[150] );
tran (\_zy_simnet_tvar_20[6][158] , \_zy_simnet_tvar_20[6].label[149] );
tran (\_zy_simnet_tvar_20[6][157] , \_zy_simnet_tvar_20[6].label[148] );
tran (\_zy_simnet_tvar_20[6][156] , \_zy_simnet_tvar_20[6].label[147] );
tran (\_zy_simnet_tvar_20[6][155] , \_zy_simnet_tvar_20[6].label[146] );
tran (\_zy_simnet_tvar_20[6][154] , \_zy_simnet_tvar_20[6].label[145] );
tran (\_zy_simnet_tvar_20[6][153] , \_zy_simnet_tvar_20[6].label[144] );
tran (\_zy_simnet_tvar_20[6][152] , \_zy_simnet_tvar_20[6].label[143] );
tran (\_zy_simnet_tvar_20[6][151] , \_zy_simnet_tvar_20[6].label[142] );
tran (\_zy_simnet_tvar_20[6][150] , \_zy_simnet_tvar_20[6].label[141] );
tran (\_zy_simnet_tvar_20[6][149] , \_zy_simnet_tvar_20[6].label[140] );
tran (\_zy_simnet_tvar_20[6][148] , \_zy_simnet_tvar_20[6].label[139] );
tran (\_zy_simnet_tvar_20[6][147] , \_zy_simnet_tvar_20[6].label[138] );
tran (\_zy_simnet_tvar_20[6][146] , \_zy_simnet_tvar_20[6].label[137] );
tran (\_zy_simnet_tvar_20[6][145] , \_zy_simnet_tvar_20[6].label[136] );
tran (\_zy_simnet_tvar_20[6][144] , \_zy_simnet_tvar_20[6].label[135] );
tran (\_zy_simnet_tvar_20[6][143] , \_zy_simnet_tvar_20[6].label[134] );
tran (\_zy_simnet_tvar_20[6][142] , \_zy_simnet_tvar_20[6].label[133] );
tran (\_zy_simnet_tvar_20[6][141] , \_zy_simnet_tvar_20[6].label[132] );
tran (\_zy_simnet_tvar_20[6][140] , \_zy_simnet_tvar_20[6].label[131] );
tran (\_zy_simnet_tvar_20[6][139] , \_zy_simnet_tvar_20[6].label[130] );
tran (\_zy_simnet_tvar_20[6][138] , \_zy_simnet_tvar_20[6].label[129] );
tran (\_zy_simnet_tvar_20[6][137] , \_zy_simnet_tvar_20[6].label[128] );
tran (\_zy_simnet_tvar_20[6][136] , \_zy_simnet_tvar_20[6].label[127] );
tran (\_zy_simnet_tvar_20[6][135] , \_zy_simnet_tvar_20[6].label[126] );
tran (\_zy_simnet_tvar_20[6][134] , \_zy_simnet_tvar_20[6].label[125] );
tran (\_zy_simnet_tvar_20[6][133] , \_zy_simnet_tvar_20[6].label[124] );
tran (\_zy_simnet_tvar_20[6][132] , \_zy_simnet_tvar_20[6].label[123] );
tran (\_zy_simnet_tvar_20[6][131] , \_zy_simnet_tvar_20[6].label[122] );
tran (\_zy_simnet_tvar_20[6][130] , \_zy_simnet_tvar_20[6].label[121] );
tran (\_zy_simnet_tvar_20[6][129] , \_zy_simnet_tvar_20[6].label[120] );
tran (\_zy_simnet_tvar_20[6][128] , \_zy_simnet_tvar_20[6].label[119] );
tran (\_zy_simnet_tvar_20[6][127] , \_zy_simnet_tvar_20[6].label[118] );
tran (\_zy_simnet_tvar_20[6][126] , \_zy_simnet_tvar_20[6].label[117] );
tran (\_zy_simnet_tvar_20[6][125] , \_zy_simnet_tvar_20[6].label[116] );
tran (\_zy_simnet_tvar_20[6][124] , \_zy_simnet_tvar_20[6].label[115] );
tran (\_zy_simnet_tvar_20[6][123] , \_zy_simnet_tvar_20[6].label[114] );
tran (\_zy_simnet_tvar_20[6][122] , \_zy_simnet_tvar_20[6].label[113] );
tran (\_zy_simnet_tvar_20[6][121] , \_zy_simnet_tvar_20[6].label[112] );
tran (\_zy_simnet_tvar_20[6][120] , \_zy_simnet_tvar_20[6].label[111] );
tran (\_zy_simnet_tvar_20[6][119] , \_zy_simnet_tvar_20[6].label[110] );
tran (\_zy_simnet_tvar_20[6][118] , \_zy_simnet_tvar_20[6].label[109] );
tran (\_zy_simnet_tvar_20[6][117] , \_zy_simnet_tvar_20[6].label[108] );
tran (\_zy_simnet_tvar_20[6][116] , \_zy_simnet_tvar_20[6].label[107] );
tran (\_zy_simnet_tvar_20[6][115] , \_zy_simnet_tvar_20[6].label[106] );
tran (\_zy_simnet_tvar_20[6][114] , \_zy_simnet_tvar_20[6].label[105] );
tran (\_zy_simnet_tvar_20[6][113] , \_zy_simnet_tvar_20[6].label[104] );
tran (\_zy_simnet_tvar_20[6][112] , \_zy_simnet_tvar_20[6].label[103] );
tran (\_zy_simnet_tvar_20[6][111] , \_zy_simnet_tvar_20[6].label[102] );
tran (\_zy_simnet_tvar_20[6][110] , \_zy_simnet_tvar_20[6].label[101] );
tran (\_zy_simnet_tvar_20[6][109] , \_zy_simnet_tvar_20[6].label[100] );
tran (\_zy_simnet_tvar_20[6][108] , \_zy_simnet_tvar_20[6].label[99] );
tran (\_zy_simnet_tvar_20[6][107] , \_zy_simnet_tvar_20[6].label[98] );
tran (\_zy_simnet_tvar_20[6][106] , \_zy_simnet_tvar_20[6].label[97] );
tran (\_zy_simnet_tvar_20[6][105] , \_zy_simnet_tvar_20[6].label[96] );
tran (\_zy_simnet_tvar_20[6][104] , \_zy_simnet_tvar_20[6].label[95] );
tran (\_zy_simnet_tvar_20[6][103] , \_zy_simnet_tvar_20[6].label[94] );
tran (\_zy_simnet_tvar_20[6][102] , \_zy_simnet_tvar_20[6].label[93] );
tran (\_zy_simnet_tvar_20[6][101] , \_zy_simnet_tvar_20[6].label[92] );
tran (\_zy_simnet_tvar_20[6][100] , \_zy_simnet_tvar_20[6].label[91] );
tran (\_zy_simnet_tvar_20[6][99] , \_zy_simnet_tvar_20[6].label[90] );
tran (\_zy_simnet_tvar_20[6][98] , \_zy_simnet_tvar_20[6].label[89] );
tran (\_zy_simnet_tvar_20[6][97] , \_zy_simnet_tvar_20[6].label[88] );
tran (\_zy_simnet_tvar_20[6][96] , \_zy_simnet_tvar_20[6].label[87] );
tran (\_zy_simnet_tvar_20[6][95] , \_zy_simnet_tvar_20[6].label[86] );
tran (\_zy_simnet_tvar_20[6][94] , \_zy_simnet_tvar_20[6].label[85] );
tran (\_zy_simnet_tvar_20[6][93] , \_zy_simnet_tvar_20[6].label[84] );
tran (\_zy_simnet_tvar_20[6][92] , \_zy_simnet_tvar_20[6].label[83] );
tran (\_zy_simnet_tvar_20[6][91] , \_zy_simnet_tvar_20[6].label[82] );
tran (\_zy_simnet_tvar_20[6][90] , \_zy_simnet_tvar_20[6].label[81] );
tran (\_zy_simnet_tvar_20[6][89] , \_zy_simnet_tvar_20[6].label[80] );
tran (\_zy_simnet_tvar_20[6][88] , \_zy_simnet_tvar_20[6].label[79] );
tran (\_zy_simnet_tvar_20[6][87] , \_zy_simnet_tvar_20[6].label[78] );
tran (\_zy_simnet_tvar_20[6][86] , \_zy_simnet_tvar_20[6].label[77] );
tran (\_zy_simnet_tvar_20[6][85] , \_zy_simnet_tvar_20[6].label[76] );
tran (\_zy_simnet_tvar_20[6][84] , \_zy_simnet_tvar_20[6].label[75] );
tran (\_zy_simnet_tvar_20[6][83] , \_zy_simnet_tvar_20[6].label[74] );
tran (\_zy_simnet_tvar_20[6][82] , \_zy_simnet_tvar_20[6].label[73] );
tran (\_zy_simnet_tvar_20[6][81] , \_zy_simnet_tvar_20[6].label[72] );
tran (\_zy_simnet_tvar_20[6][80] , \_zy_simnet_tvar_20[6].label[71] );
tran (\_zy_simnet_tvar_20[6][79] , \_zy_simnet_tvar_20[6].label[70] );
tran (\_zy_simnet_tvar_20[6][78] , \_zy_simnet_tvar_20[6].label[69] );
tran (\_zy_simnet_tvar_20[6][77] , \_zy_simnet_tvar_20[6].label[68] );
tran (\_zy_simnet_tvar_20[6][76] , \_zy_simnet_tvar_20[6].label[67] );
tran (\_zy_simnet_tvar_20[6][75] , \_zy_simnet_tvar_20[6].label[66] );
tran (\_zy_simnet_tvar_20[6][74] , \_zy_simnet_tvar_20[6].label[65] );
tran (\_zy_simnet_tvar_20[6][73] , \_zy_simnet_tvar_20[6].label[64] );
tran (\_zy_simnet_tvar_20[6][72] , \_zy_simnet_tvar_20[6].label[63] );
tran (\_zy_simnet_tvar_20[6][71] , \_zy_simnet_tvar_20[6].label[62] );
tran (\_zy_simnet_tvar_20[6][70] , \_zy_simnet_tvar_20[6].label[61] );
tran (\_zy_simnet_tvar_20[6][69] , \_zy_simnet_tvar_20[6].label[60] );
tran (\_zy_simnet_tvar_20[6][68] , \_zy_simnet_tvar_20[6].label[59] );
tran (\_zy_simnet_tvar_20[6][67] , \_zy_simnet_tvar_20[6].label[58] );
tran (\_zy_simnet_tvar_20[6][66] , \_zy_simnet_tvar_20[6].label[57] );
tran (\_zy_simnet_tvar_20[6][65] , \_zy_simnet_tvar_20[6].label[56] );
tran (\_zy_simnet_tvar_20[6][64] , \_zy_simnet_tvar_20[6].label[55] );
tran (\_zy_simnet_tvar_20[6][63] , \_zy_simnet_tvar_20[6].label[54] );
tran (\_zy_simnet_tvar_20[6][62] , \_zy_simnet_tvar_20[6].label[53] );
tran (\_zy_simnet_tvar_20[6][61] , \_zy_simnet_tvar_20[6].label[52] );
tran (\_zy_simnet_tvar_20[6][60] , \_zy_simnet_tvar_20[6].label[51] );
tran (\_zy_simnet_tvar_20[6][59] , \_zy_simnet_tvar_20[6].label[50] );
tran (\_zy_simnet_tvar_20[6][58] , \_zy_simnet_tvar_20[6].label[49] );
tran (\_zy_simnet_tvar_20[6][57] , \_zy_simnet_tvar_20[6].label[48] );
tran (\_zy_simnet_tvar_20[6][56] , \_zy_simnet_tvar_20[6].label[47] );
tran (\_zy_simnet_tvar_20[6][55] , \_zy_simnet_tvar_20[6].label[46] );
tran (\_zy_simnet_tvar_20[6][54] , \_zy_simnet_tvar_20[6].label[45] );
tran (\_zy_simnet_tvar_20[6][53] , \_zy_simnet_tvar_20[6].label[44] );
tran (\_zy_simnet_tvar_20[6][52] , \_zy_simnet_tvar_20[6].label[43] );
tran (\_zy_simnet_tvar_20[6][51] , \_zy_simnet_tvar_20[6].label[42] );
tran (\_zy_simnet_tvar_20[6][50] , \_zy_simnet_tvar_20[6].label[41] );
tran (\_zy_simnet_tvar_20[6][49] , \_zy_simnet_tvar_20[6].label[40] );
tran (\_zy_simnet_tvar_20[6][48] , \_zy_simnet_tvar_20[6].label[39] );
tran (\_zy_simnet_tvar_20[6][47] , \_zy_simnet_tvar_20[6].label[38] );
tran (\_zy_simnet_tvar_20[6][46] , \_zy_simnet_tvar_20[6].label[37] );
tran (\_zy_simnet_tvar_20[6][45] , \_zy_simnet_tvar_20[6].label[36] );
tran (\_zy_simnet_tvar_20[6][44] , \_zy_simnet_tvar_20[6].label[35] );
tran (\_zy_simnet_tvar_20[6][43] , \_zy_simnet_tvar_20[6].label[34] );
tran (\_zy_simnet_tvar_20[6][42] , \_zy_simnet_tvar_20[6].label[33] );
tran (\_zy_simnet_tvar_20[6][41] , \_zy_simnet_tvar_20[6].label[32] );
tran (\_zy_simnet_tvar_20[6][40] , \_zy_simnet_tvar_20[6].label[31] );
tran (\_zy_simnet_tvar_20[6][39] , \_zy_simnet_tvar_20[6].label[30] );
tran (\_zy_simnet_tvar_20[6][38] , \_zy_simnet_tvar_20[6].label[29] );
tran (\_zy_simnet_tvar_20[6][37] , \_zy_simnet_tvar_20[6].label[28] );
tran (\_zy_simnet_tvar_20[6][36] , \_zy_simnet_tvar_20[6].label[27] );
tran (\_zy_simnet_tvar_20[6][35] , \_zy_simnet_tvar_20[6].label[26] );
tran (\_zy_simnet_tvar_20[6][34] , \_zy_simnet_tvar_20[6].label[25] );
tran (\_zy_simnet_tvar_20[6][33] , \_zy_simnet_tvar_20[6].label[24] );
tran (\_zy_simnet_tvar_20[6][32] , \_zy_simnet_tvar_20[6].label[23] );
tran (\_zy_simnet_tvar_20[6][31] , \_zy_simnet_tvar_20[6].label[22] );
tran (\_zy_simnet_tvar_20[6][30] , \_zy_simnet_tvar_20[6].label[21] );
tran (\_zy_simnet_tvar_20[6][29] , \_zy_simnet_tvar_20[6].label[20] );
tran (\_zy_simnet_tvar_20[6][28] , \_zy_simnet_tvar_20[6].label[19] );
tran (\_zy_simnet_tvar_20[6][27] , \_zy_simnet_tvar_20[6].label[18] );
tran (\_zy_simnet_tvar_20[6][26] , \_zy_simnet_tvar_20[6].label[17] );
tran (\_zy_simnet_tvar_20[6][25] , \_zy_simnet_tvar_20[6].label[16] );
tran (\_zy_simnet_tvar_20[6][24] , \_zy_simnet_tvar_20[6].label[15] );
tran (\_zy_simnet_tvar_20[6][23] , \_zy_simnet_tvar_20[6].label[14] );
tran (\_zy_simnet_tvar_20[6][22] , \_zy_simnet_tvar_20[6].label[13] );
tran (\_zy_simnet_tvar_20[6][21] , \_zy_simnet_tvar_20[6].label[12] );
tran (\_zy_simnet_tvar_20[6][20] , \_zy_simnet_tvar_20[6].label[11] );
tran (\_zy_simnet_tvar_20[6][19] , \_zy_simnet_tvar_20[6].label[10] );
tran (\_zy_simnet_tvar_20[6][18] , \_zy_simnet_tvar_20[6].label[9] );
tran (\_zy_simnet_tvar_20[6][17] , \_zy_simnet_tvar_20[6].label[8] );
tran (\_zy_simnet_tvar_20[6][16] , \_zy_simnet_tvar_20[6].label[7] );
tran (\_zy_simnet_tvar_20[6][15] , \_zy_simnet_tvar_20[6].label[6] );
tran (\_zy_simnet_tvar_20[6][14] , \_zy_simnet_tvar_20[6].label[5] );
tran (\_zy_simnet_tvar_20[6][13] , \_zy_simnet_tvar_20[6].label[4] );
tran (\_zy_simnet_tvar_20[6][12] , \_zy_simnet_tvar_20[6].label[3] );
tran (\_zy_simnet_tvar_20[6][11] , \_zy_simnet_tvar_20[6].label[2] );
tran (\_zy_simnet_tvar_20[6][10] , \_zy_simnet_tvar_20[6].label[1] );
tran (\_zy_simnet_tvar_20[6][9] , \_zy_simnet_tvar_20[6].label[0] );
tran (\_zy_simnet_tvar_20[6][8] , \_zy_simnet_tvar_20[6].delimiter_valid[0] );
tran (\_zy_simnet_tvar_20[6][7] , \_zy_simnet_tvar_20[6].delimiter[7] );
tran (\_zy_simnet_tvar_20[6][6] , \_zy_simnet_tvar_20[6].delimiter[6] );
tran (\_zy_simnet_tvar_20[6][5] , \_zy_simnet_tvar_20[6].delimiter[5] );
tran (\_zy_simnet_tvar_20[6][4] , \_zy_simnet_tvar_20[6].delimiter[4] );
tran (\_zy_simnet_tvar_20[6][3] , \_zy_simnet_tvar_20[6].delimiter[3] );
tran (\_zy_simnet_tvar_20[6][2] , \_zy_simnet_tvar_20[6].delimiter[2] );
tran (\_zy_simnet_tvar_20[6][1] , \_zy_simnet_tvar_20[6].delimiter[1] );
tran (\_zy_simnet_tvar_20[6][0] , \_zy_simnet_tvar_20[6].delimiter[0] );
tran (\_zy_simnet_tvar_20[5][271] , \_zy_simnet_tvar_20[5].guid_size[0] );
tran (\_zy_simnet_tvar_20[5][270] , \_zy_simnet_tvar_20[5].label_size[5] );
tran (\_zy_simnet_tvar_20[5][269] , \_zy_simnet_tvar_20[5].label_size[4] );
tran (\_zy_simnet_tvar_20[5][268] , \_zy_simnet_tvar_20[5].label_size[3] );
tran (\_zy_simnet_tvar_20[5][267] , \_zy_simnet_tvar_20[5].label_size[2] );
tran (\_zy_simnet_tvar_20[5][266] , \_zy_simnet_tvar_20[5].label_size[1] );
tran (\_zy_simnet_tvar_20[5][265] , \_zy_simnet_tvar_20[5].label_size[0] );
tran (\_zy_simnet_tvar_20[5][264] , \_zy_simnet_tvar_20[5].label[255] );
tran (\_zy_simnet_tvar_20[5][263] , \_zy_simnet_tvar_20[5].label[254] );
tran (\_zy_simnet_tvar_20[5][262] , \_zy_simnet_tvar_20[5].label[253] );
tran (\_zy_simnet_tvar_20[5][261] , \_zy_simnet_tvar_20[5].label[252] );
tran (\_zy_simnet_tvar_20[5][260] , \_zy_simnet_tvar_20[5].label[251] );
tran (\_zy_simnet_tvar_20[5][259] , \_zy_simnet_tvar_20[5].label[250] );
tran (\_zy_simnet_tvar_20[5][258] , \_zy_simnet_tvar_20[5].label[249] );
tran (\_zy_simnet_tvar_20[5][257] , \_zy_simnet_tvar_20[5].label[248] );
tran (\_zy_simnet_tvar_20[5][256] , \_zy_simnet_tvar_20[5].label[247] );
tran (\_zy_simnet_tvar_20[5][255] , \_zy_simnet_tvar_20[5].label[246] );
tran (\_zy_simnet_tvar_20[5][254] , \_zy_simnet_tvar_20[5].label[245] );
tran (\_zy_simnet_tvar_20[5][253] , \_zy_simnet_tvar_20[5].label[244] );
tran (\_zy_simnet_tvar_20[5][252] , \_zy_simnet_tvar_20[5].label[243] );
tran (\_zy_simnet_tvar_20[5][251] , \_zy_simnet_tvar_20[5].label[242] );
tran (\_zy_simnet_tvar_20[5][250] , \_zy_simnet_tvar_20[5].label[241] );
tran (\_zy_simnet_tvar_20[5][249] , \_zy_simnet_tvar_20[5].label[240] );
tran (\_zy_simnet_tvar_20[5][248] , \_zy_simnet_tvar_20[5].label[239] );
tran (\_zy_simnet_tvar_20[5][247] , \_zy_simnet_tvar_20[5].label[238] );
tran (\_zy_simnet_tvar_20[5][246] , \_zy_simnet_tvar_20[5].label[237] );
tran (\_zy_simnet_tvar_20[5][245] , \_zy_simnet_tvar_20[5].label[236] );
tran (\_zy_simnet_tvar_20[5][244] , \_zy_simnet_tvar_20[5].label[235] );
tran (\_zy_simnet_tvar_20[5][243] , \_zy_simnet_tvar_20[5].label[234] );
tran (\_zy_simnet_tvar_20[5][242] , \_zy_simnet_tvar_20[5].label[233] );
tran (\_zy_simnet_tvar_20[5][241] , \_zy_simnet_tvar_20[5].label[232] );
tran (\_zy_simnet_tvar_20[5][240] , \_zy_simnet_tvar_20[5].label[231] );
tran (\_zy_simnet_tvar_20[5][239] , \_zy_simnet_tvar_20[5].label[230] );
tran (\_zy_simnet_tvar_20[5][238] , \_zy_simnet_tvar_20[5].label[229] );
tran (\_zy_simnet_tvar_20[5][237] , \_zy_simnet_tvar_20[5].label[228] );
tran (\_zy_simnet_tvar_20[5][236] , \_zy_simnet_tvar_20[5].label[227] );
tran (\_zy_simnet_tvar_20[5][235] , \_zy_simnet_tvar_20[5].label[226] );
tran (\_zy_simnet_tvar_20[5][234] , \_zy_simnet_tvar_20[5].label[225] );
tran (\_zy_simnet_tvar_20[5][233] , \_zy_simnet_tvar_20[5].label[224] );
tran (\_zy_simnet_tvar_20[5][232] , \_zy_simnet_tvar_20[5].label[223] );
tran (\_zy_simnet_tvar_20[5][231] , \_zy_simnet_tvar_20[5].label[222] );
tran (\_zy_simnet_tvar_20[5][230] , \_zy_simnet_tvar_20[5].label[221] );
tran (\_zy_simnet_tvar_20[5][229] , \_zy_simnet_tvar_20[5].label[220] );
tran (\_zy_simnet_tvar_20[5][228] , \_zy_simnet_tvar_20[5].label[219] );
tran (\_zy_simnet_tvar_20[5][227] , \_zy_simnet_tvar_20[5].label[218] );
tran (\_zy_simnet_tvar_20[5][226] , \_zy_simnet_tvar_20[5].label[217] );
tran (\_zy_simnet_tvar_20[5][225] , \_zy_simnet_tvar_20[5].label[216] );
tran (\_zy_simnet_tvar_20[5][224] , \_zy_simnet_tvar_20[5].label[215] );
tran (\_zy_simnet_tvar_20[5][223] , \_zy_simnet_tvar_20[5].label[214] );
tran (\_zy_simnet_tvar_20[5][222] , \_zy_simnet_tvar_20[5].label[213] );
tran (\_zy_simnet_tvar_20[5][221] , \_zy_simnet_tvar_20[5].label[212] );
tran (\_zy_simnet_tvar_20[5][220] , \_zy_simnet_tvar_20[5].label[211] );
tran (\_zy_simnet_tvar_20[5][219] , \_zy_simnet_tvar_20[5].label[210] );
tran (\_zy_simnet_tvar_20[5][218] , \_zy_simnet_tvar_20[5].label[209] );
tran (\_zy_simnet_tvar_20[5][217] , \_zy_simnet_tvar_20[5].label[208] );
tran (\_zy_simnet_tvar_20[5][216] , \_zy_simnet_tvar_20[5].label[207] );
tran (\_zy_simnet_tvar_20[5][215] , \_zy_simnet_tvar_20[5].label[206] );
tran (\_zy_simnet_tvar_20[5][214] , \_zy_simnet_tvar_20[5].label[205] );
tran (\_zy_simnet_tvar_20[5][213] , \_zy_simnet_tvar_20[5].label[204] );
tran (\_zy_simnet_tvar_20[5][212] , \_zy_simnet_tvar_20[5].label[203] );
tran (\_zy_simnet_tvar_20[5][211] , \_zy_simnet_tvar_20[5].label[202] );
tran (\_zy_simnet_tvar_20[5][210] , \_zy_simnet_tvar_20[5].label[201] );
tran (\_zy_simnet_tvar_20[5][209] , \_zy_simnet_tvar_20[5].label[200] );
tran (\_zy_simnet_tvar_20[5][208] , \_zy_simnet_tvar_20[5].label[199] );
tran (\_zy_simnet_tvar_20[5][207] , \_zy_simnet_tvar_20[5].label[198] );
tran (\_zy_simnet_tvar_20[5][206] , \_zy_simnet_tvar_20[5].label[197] );
tran (\_zy_simnet_tvar_20[5][205] , \_zy_simnet_tvar_20[5].label[196] );
tran (\_zy_simnet_tvar_20[5][204] , \_zy_simnet_tvar_20[5].label[195] );
tran (\_zy_simnet_tvar_20[5][203] , \_zy_simnet_tvar_20[5].label[194] );
tran (\_zy_simnet_tvar_20[5][202] , \_zy_simnet_tvar_20[5].label[193] );
tran (\_zy_simnet_tvar_20[5][201] , \_zy_simnet_tvar_20[5].label[192] );
tran (\_zy_simnet_tvar_20[5][200] , \_zy_simnet_tvar_20[5].label[191] );
tran (\_zy_simnet_tvar_20[5][199] , \_zy_simnet_tvar_20[5].label[190] );
tran (\_zy_simnet_tvar_20[5][198] , \_zy_simnet_tvar_20[5].label[189] );
tran (\_zy_simnet_tvar_20[5][197] , \_zy_simnet_tvar_20[5].label[188] );
tran (\_zy_simnet_tvar_20[5][196] , \_zy_simnet_tvar_20[5].label[187] );
tran (\_zy_simnet_tvar_20[5][195] , \_zy_simnet_tvar_20[5].label[186] );
tran (\_zy_simnet_tvar_20[5][194] , \_zy_simnet_tvar_20[5].label[185] );
tran (\_zy_simnet_tvar_20[5][193] , \_zy_simnet_tvar_20[5].label[184] );
tran (\_zy_simnet_tvar_20[5][192] , \_zy_simnet_tvar_20[5].label[183] );
tran (\_zy_simnet_tvar_20[5][191] , \_zy_simnet_tvar_20[5].label[182] );
tran (\_zy_simnet_tvar_20[5][190] , \_zy_simnet_tvar_20[5].label[181] );
tran (\_zy_simnet_tvar_20[5][189] , \_zy_simnet_tvar_20[5].label[180] );
tran (\_zy_simnet_tvar_20[5][188] , \_zy_simnet_tvar_20[5].label[179] );
tran (\_zy_simnet_tvar_20[5][187] , \_zy_simnet_tvar_20[5].label[178] );
tran (\_zy_simnet_tvar_20[5][186] , \_zy_simnet_tvar_20[5].label[177] );
tran (\_zy_simnet_tvar_20[5][185] , \_zy_simnet_tvar_20[5].label[176] );
tran (\_zy_simnet_tvar_20[5][184] , \_zy_simnet_tvar_20[5].label[175] );
tran (\_zy_simnet_tvar_20[5][183] , \_zy_simnet_tvar_20[5].label[174] );
tran (\_zy_simnet_tvar_20[5][182] , \_zy_simnet_tvar_20[5].label[173] );
tran (\_zy_simnet_tvar_20[5][181] , \_zy_simnet_tvar_20[5].label[172] );
tran (\_zy_simnet_tvar_20[5][180] , \_zy_simnet_tvar_20[5].label[171] );
tran (\_zy_simnet_tvar_20[5][179] , \_zy_simnet_tvar_20[5].label[170] );
tran (\_zy_simnet_tvar_20[5][178] , \_zy_simnet_tvar_20[5].label[169] );
tran (\_zy_simnet_tvar_20[5][177] , \_zy_simnet_tvar_20[5].label[168] );
tran (\_zy_simnet_tvar_20[5][176] , \_zy_simnet_tvar_20[5].label[167] );
tran (\_zy_simnet_tvar_20[5][175] , \_zy_simnet_tvar_20[5].label[166] );
tran (\_zy_simnet_tvar_20[5][174] , \_zy_simnet_tvar_20[5].label[165] );
tran (\_zy_simnet_tvar_20[5][173] , \_zy_simnet_tvar_20[5].label[164] );
tran (\_zy_simnet_tvar_20[5][172] , \_zy_simnet_tvar_20[5].label[163] );
tran (\_zy_simnet_tvar_20[5][171] , \_zy_simnet_tvar_20[5].label[162] );
tran (\_zy_simnet_tvar_20[5][170] , \_zy_simnet_tvar_20[5].label[161] );
tran (\_zy_simnet_tvar_20[5][169] , \_zy_simnet_tvar_20[5].label[160] );
tran (\_zy_simnet_tvar_20[5][168] , \_zy_simnet_tvar_20[5].label[159] );
tran (\_zy_simnet_tvar_20[5][167] , \_zy_simnet_tvar_20[5].label[158] );
tran (\_zy_simnet_tvar_20[5][166] , \_zy_simnet_tvar_20[5].label[157] );
tran (\_zy_simnet_tvar_20[5][165] , \_zy_simnet_tvar_20[5].label[156] );
tran (\_zy_simnet_tvar_20[5][164] , \_zy_simnet_tvar_20[5].label[155] );
tran (\_zy_simnet_tvar_20[5][163] , \_zy_simnet_tvar_20[5].label[154] );
tran (\_zy_simnet_tvar_20[5][162] , \_zy_simnet_tvar_20[5].label[153] );
tran (\_zy_simnet_tvar_20[5][161] , \_zy_simnet_tvar_20[5].label[152] );
tran (\_zy_simnet_tvar_20[5][160] , \_zy_simnet_tvar_20[5].label[151] );
tran (\_zy_simnet_tvar_20[5][159] , \_zy_simnet_tvar_20[5].label[150] );
tran (\_zy_simnet_tvar_20[5][158] , \_zy_simnet_tvar_20[5].label[149] );
tran (\_zy_simnet_tvar_20[5][157] , \_zy_simnet_tvar_20[5].label[148] );
tran (\_zy_simnet_tvar_20[5][156] , \_zy_simnet_tvar_20[5].label[147] );
tran (\_zy_simnet_tvar_20[5][155] , \_zy_simnet_tvar_20[5].label[146] );
tran (\_zy_simnet_tvar_20[5][154] , \_zy_simnet_tvar_20[5].label[145] );
tran (\_zy_simnet_tvar_20[5][153] , \_zy_simnet_tvar_20[5].label[144] );
tran (\_zy_simnet_tvar_20[5][152] , \_zy_simnet_tvar_20[5].label[143] );
tran (\_zy_simnet_tvar_20[5][151] , \_zy_simnet_tvar_20[5].label[142] );
tran (\_zy_simnet_tvar_20[5][150] , \_zy_simnet_tvar_20[5].label[141] );
tran (\_zy_simnet_tvar_20[5][149] , \_zy_simnet_tvar_20[5].label[140] );
tran (\_zy_simnet_tvar_20[5][148] , \_zy_simnet_tvar_20[5].label[139] );
tran (\_zy_simnet_tvar_20[5][147] , \_zy_simnet_tvar_20[5].label[138] );
tran (\_zy_simnet_tvar_20[5][146] , \_zy_simnet_tvar_20[5].label[137] );
tran (\_zy_simnet_tvar_20[5][145] , \_zy_simnet_tvar_20[5].label[136] );
tran (\_zy_simnet_tvar_20[5][144] , \_zy_simnet_tvar_20[5].label[135] );
tran (\_zy_simnet_tvar_20[5][143] , \_zy_simnet_tvar_20[5].label[134] );
tran (\_zy_simnet_tvar_20[5][142] , \_zy_simnet_tvar_20[5].label[133] );
tran (\_zy_simnet_tvar_20[5][141] , \_zy_simnet_tvar_20[5].label[132] );
tran (\_zy_simnet_tvar_20[5][140] , \_zy_simnet_tvar_20[5].label[131] );
tran (\_zy_simnet_tvar_20[5][139] , \_zy_simnet_tvar_20[5].label[130] );
tran (\_zy_simnet_tvar_20[5][138] , \_zy_simnet_tvar_20[5].label[129] );
tran (\_zy_simnet_tvar_20[5][137] , \_zy_simnet_tvar_20[5].label[128] );
tran (\_zy_simnet_tvar_20[5][136] , \_zy_simnet_tvar_20[5].label[127] );
tran (\_zy_simnet_tvar_20[5][135] , \_zy_simnet_tvar_20[5].label[126] );
tran (\_zy_simnet_tvar_20[5][134] , \_zy_simnet_tvar_20[5].label[125] );
tran (\_zy_simnet_tvar_20[5][133] , \_zy_simnet_tvar_20[5].label[124] );
tran (\_zy_simnet_tvar_20[5][132] , \_zy_simnet_tvar_20[5].label[123] );
tran (\_zy_simnet_tvar_20[5][131] , \_zy_simnet_tvar_20[5].label[122] );
tran (\_zy_simnet_tvar_20[5][130] , \_zy_simnet_tvar_20[5].label[121] );
tran (\_zy_simnet_tvar_20[5][129] , \_zy_simnet_tvar_20[5].label[120] );
tran (\_zy_simnet_tvar_20[5][128] , \_zy_simnet_tvar_20[5].label[119] );
tran (\_zy_simnet_tvar_20[5][127] , \_zy_simnet_tvar_20[5].label[118] );
tran (\_zy_simnet_tvar_20[5][126] , \_zy_simnet_tvar_20[5].label[117] );
tran (\_zy_simnet_tvar_20[5][125] , \_zy_simnet_tvar_20[5].label[116] );
tran (\_zy_simnet_tvar_20[5][124] , \_zy_simnet_tvar_20[5].label[115] );
tran (\_zy_simnet_tvar_20[5][123] , \_zy_simnet_tvar_20[5].label[114] );
tran (\_zy_simnet_tvar_20[5][122] , \_zy_simnet_tvar_20[5].label[113] );
tran (\_zy_simnet_tvar_20[5][121] , \_zy_simnet_tvar_20[5].label[112] );
tran (\_zy_simnet_tvar_20[5][120] , \_zy_simnet_tvar_20[5].label[111] );
tran (\_zy_simnet_tvar_20[5][119] , \_zy_simnet_tvar_20[5].label[110] );
tran (\_zy_simnet_tvar_20[5][118] , \_zy_simnet_tvar_20[5].label[109] );
tran (\_zy_simnet_tvar_20[5][117] , \_zy_simnet_tvar_20[5].label[108] );
tran (\_zy_simnet_tvar_20[5][116] , \_zy_simnet_tvar_20[5].label[107] );
tran (\_zy_simnet_tvar_20[5][115] , \_zy_simnet_tvar_20[5].label[106] );
tran (\_zy_simnet_tvar_20[5][114] , \_zy_simnet_tvar_20[5].label[105] );
tran (\_zy_simnet_tvar_20[5][113] , \_zy_simnet_tvar_20[5].label[104] );
tran (\_zy_simnet_tvar_20[5][112] , \_zy_simnet_tvar_20[5].label[103] );
tran (\_zy_simnet_tvar_20[5][111] , \_zy_simnet_tvar_20[5].label[102] );
tran (\_zy_simnet_tvar_20[5][110] , \_zy_simnet_tvar_20[5].label[101] );
tran (\_zy_simnet_tvar_20[5][109] , \_zy_simnet_tvar_20[5].label[100] );
tran (\_zy_simnet_tvar_20[5][108] , \_zy_simnet_tvar_20[5].label[99] );
tran (\_zy_simnet_tvar_20[5][107] , \_zy_simnet_tvar_20[5].label[98] );
tran (\_zy_simnet_tvar_20[5][106] , \_zy_simnet_tvar_20[5].label[97] );
tran (\_zy_simnet_tvar_20[5][105] , \_zy_simnet_tvar_20[5].label[96] );
tran (\_zy_simnet_tvar_20[5][104] , \_zy_simnet_tvar_20[5].label[95] );
tran (\_zy_simnet_tvar_20[5][103] , \_zy_simnet_tvar_20[5].label[94] );
tran (\_zy_simnet_tvar_20[5][102] , \_zy_simnet_tvar_20[5].label[93] );
tran (\_zy_simnet_tvar_20[5][101] , \_zy_simnet_tvar_20[5].label[92] );
tran (\_zy_simnet_tvar_20[5][100] , \_zy_simnet_tvar_20[5].label[91] );
tran (\_zy_simnet_tvar_20[5][99] , \_zy_simnet_tvar_20[5].label[90] );
tran (\_zy_simnet_tvar_20[5][98] , \_zy_simnet_tvar_20[5].label[89] );
tran (\_zy_simnet_tvar_20[5][97] , \_zy_simnet_tvar_20[5].label[88] );
tran (\_zy_simnet_tvar_20[5][96] , \_zy_simnet_tvar_20[5].label[87] );
tran (\_zy_simnet_tvar_20[5][95] , \_zy_simnet_tvar_20[5].label[86] );
tran (\_zy_simnet_tvar_20[5][94] , \_zy_simnet_tvar_20[5].label[85] );
tran (\_zy_simnet_tvar_20[5][93] , \_zy_simnet_tvar_20[5].label[84] );
tran (\_zy_simnet_tvar_20[5][92] , \_zy_simnet_tvar_20[5].label[83] );
tran (\_zy_simnet_tvar_20[5][91] , \_zy_simnet_tvar_20[5].label[82] );
tran (\_zy_simnet_tvar_20[5][90] , \_zy_simnet_tvar_20[5].label[81] );
tran (\_zy_simnet_tvar_20[5][89] , \_zy_simnet_tvar_20[5].label[80] );
tran (\_zy_simnet_tvar_20[5][88] , \_zy_simnet_tvar_20[5].label[79] );
tran (\_zy_simnet_tvar_20[5][87] , \_zy_simnet_tvar_20[5].label[78] );
tran (\_zy_simnet_tvar_20[5][86] , \_zy_simnet_tvar_20[5].label[77] );
tran (\_zy_simnet_tvar_20[5][85] , \_zy_simnet_tvar_20[5].label[76] );
tran (\_zy_simnet_tvar_20[5][84] , \_zy_simnet_tvar_20[5].label[75] );
tran (\_zy_simnet_tvar_20[5][83] , \_zy_simnet_tvar_20[5].label[74] );
tran (\_zy_simnet_tvar_20[5][82] , \_zy_simnet_tvar_20[5].label[73] );
tran (\_zy_simnet_tvar_20[5][81] , \_zy_simnet_tvar_20[5].label[72] );
tran (\_zy_simnet_tvar_20[5][80] , \_zy_simnet_tvar_20[5].label[71] );
tran (\_zy_simnet_tvar_20[5][79] , \_zy_simnet_tvar_20[5].label[70] );
tran (\_zy_simnet_tvar_20[5][78] , \_zy_simnet_tvar_20[5].label[69] );
tran (\_zy_simnet_tvar_20[5][77] , \_zy_simnet_tvar_20[5].label[68] );
tran (\_zy_simnet_tvar_20[5][76] , \_zy_simnet_tvar_20[5].label[67] );
tran (\_zy_simnet_tvar_20[5][75] , \_zy_simnet_tvar_20[5].label[66] );
tran (\_zy_simnet_tvar_20[5][74] , \_zy_simnet_tvar_20[5].label[65] );
tran (\_zy_simnet_tvar_20[5][73] , \_zy_simnet_tvar_20[5].label[64] );
tran (\_zy_simnet_tvar_20[5][72] , \_zy_simnet_tvar_20[5].label[63] );
tran (\_zy_simnet_tvar_20[5][71] , \_zy_simnet_tvar_20[5].label[62] );
tran (\_zy_simnet_tvar_20[5][70] , \_zy_simnet_tvar_20[5].label[61] );
tran (\_zy_simnet_tvar_20[5][69] , \_zy_simnet_tvar_20[5].label[60] );
tran (\_zy_simnet_tvar_20[5][68] , \_zy_simnet_tvar_20[5].label[59] );
tran (\_zy_simnet_tvar_20[5][67] , \_zy_simnet_tvar_20[5].label[58] );
tran (\_zy_simnet_tvar_20[5][66] , \_zy_simnet_tvar_20[5].label[57] );
tran (\_zy_simnet_tvar_20[5][65] , \_zy_simnet_tvar_20[5].label[56] );
tran (\_zy_simnet_tvar_20[5][64] , \_zy_simnet_tvar_20[5].label[55] );
tran (\_zy_simnet_tvar_20[5][63] , \_zy_simnet_tvar_20[5].label[54] );
tran (\_zy_simnet_tvar_20[5][62] , \_zy_simnet_tvar_20[5].label[53] );
tran (\_zy_simnet_tvar_20[5][61] , \_zy_simnet_tvar_20[5].label[52] );
tran (\_zy_simnet_tvar_20[5][60] , \_zy_simnet_tvar_20[5].label[51] );
tran (\_zy_simnet_tvar_20[5][59] , \_zy_simnet_tvar_20[5].label[50] );
tran (\_zy_simnet_tvar_20[5][58] , \_zy_simnet_tvar_20[5].label[49] );
tran (\_zy_simnet_tvar_20[5][57] , \_zy_simnet_tvar_20[5].label[48] );
tran (\_zy_simnet_tvar_20[5][56] , \_zy_simnet_tvar_20[5].label[47] );
tran (\_zy_simnet_tvar_20[5][55] , \_zy_simnet_tvar_20[5].label[46] );
tran (\_zy_simnet_tvar_20[5][54] , \_zy_simnet_tvar_20[5].label[45] );
tran (\_zy_simnet_tvar_20[5][53] , \_zy_simnet_tvar_20[5].label[44] );
tran (\_zy_simnet_tvar_20[5][52] , \_zy_simnet_tvar_20[5].label[43] );
tran (\_zy_simnet_tvar_20[5][51] , \_zy_simnet_tvar_20[5].label[42] );
tran (\_zy_simnet_tvar_20[5][50] , \_zy_simnet_tvar_20[5].label[41] );
tran (\_zy_simnet_tvar_20[5][49] , \_zy_simnet_tvar_20[5].label[40] );
tran (\_zy_simnet_tvar_20[5][48] , \_zy_simnet_tvar_20[5].label[39] );
tran (\_zy_simnet_tvar_20[5][47] , \_zy_simnet_tvar_20[5].label[38] );
tran (\_zy_simnet_tvar_20[5][46] , \_zy_simnet_tvar_20[5].label[37] );
tran (\_zy_simnet_tvar_20[5][45] , \_zy_simnet_tvar_20[5].label[36] );
tran (\_zy_simnet_tvar_20[5][44] , \_zy_simnet_tvar_20[5].label[35] );
tran (\_zy_simnet_tvar_20[5][43] , \_zy_simnet_tvar_20[5].label[34] );
tran (\_zy_simnet_tvar_20[5][42] , \_zy_simnet_tvar_20[5].label[33] );
tran (\_zy_simnet_tvar_20[5][41] , \_zy_simnet_tvar_20[5].label[32] );
tran (\_zy_simnet_tvar_20[5][40] , \_zy_simnet_tvar_20[5].label[31] );
tran (\_zy_simnet_tvar_20[5][39] , \_zy_simnet_tvar_20[5].label[30] );
tran (\_zy_simnet_tvar_20[5][38] , \_zy_simnet_tvar_20[5].label[29] );
tran (\_zy_simnet_tvar_20[5][37] , \_zy_simnet_tvar_20[5].label[28] );
tran (\_zy_simnet_tvar_20[5][36] , \_zy_simnet_tvar_20[5].label[27] );
tran (\_zy_simnet_tvar_20[5][35] , \_zy_simnet_tvar_20[5].label[26] );
tran (\_zy_simnet_tvar_20[5][34] , \_zy_simnet_tvar_20[5].label[25] );
tran (\_zy_simnet_tvar_20[5][33] , \_zy_simnet_tvar_20[5].label[24] );
tran (\_zy_simnet_tvar_20[5][32] , \_zy_simnet_tvar_20[5].label[23] );
tran (\_zy_simnet_tvar_20[5][31] , \_zy_simnet_tvar_20[5].label[22] );
tran (\_zy_simnet_tvar_20[5][30] , \_zy_simnet_tvar_20[5].label[21] );
tran (\_zy_simnet_tvar_20[5][29] , \_zy_simnet_tvar_20[5].label[20] );
tran (\_zy_simnet_tvar_20[5][28] , \_zy_simnet_tvar_20[5].label[19] );
tran (\_zy_simnet_tvar_20[5][27] , \_zy_simnet_tvar_20[5].label[18] );
tran (\_zy_simnet_tvar_20[5][26] , \_zy_simnet_tvar_20[5].label[17] );
tran (\_zy_simnet_tvar_20[5][25] , \_zy_simnet_tvar_20[5].label[16] );
tran (\_zy_simnet_tvar_20[5][24] , \_zy_simnet_tvar_20[5].label[15] );
tran (\_zy_simnet_tvar_20[5][23] , \_zy_simnet_tvar_20[5].label[14] );
tran (\_zy_simnet_tvar_20[5][22] , \_zy_simnet_tvar_20[5].label[13] );
tran (\_zy_simnet_tvar_20[5][21] , \_zy_simnet_tvar_20[5].label[12] );
tran (\_zy_simnet_tvar_20[5][20] , \_zy_simnet_tvar_20[5].label[11] );
tran (\_zy_simnet_tvar_20[5][19] , \_zy_simnet_tvar_20[5].label[10] );
tran (\_zy_simnet_tvar_20[5][18] , \_zy_simnet_tvar_20[5].label[9] );
tran (\_zy_simnet_tvar_20[5][17] , \_zy_simnet_tvar_20[5].label[8] );
tran (\_zy_simnet_tvar_20[5][16] , \_zy_simnet_tvar_20[5].label[7] );
tran (\_zy_simnet_tvar_20[5][15] , \_zy_simnet_tvar_20[5].label[6] );
tran (\_zy_simnet_tvar_20[5][14] , \_zy_simnet_tvar_20[5].label[5] );
tran (\_zy_simnet_tvar_20[5][13] , \_zy_simnet_tvar_20[5].label[4] );
tran (\_zy_simnet_tvar_20[5][12] , \_zy_simnet_tvar_20[5].label[3] );
tran (\_zy_simnet_tvar_20[5][11] , \_zy_simnet_tvar_20[5].label[2] );
tran (\_zy_simnet_tvar_20[5][10] , \_zy_simnet_tvar_20[5].label[1] );
tran (\_zy_simnet_tvar_20[5][9] , \_zy_simnet_tvar_20[5].label[0] );
tran (\_zy_simnet_tvar_20[5][8] , \_zy_simnet_tvar_20[5].delimiter_valid[0] );
tran (\_zy_simnet_tvar_20[5][7] , \_zy_simnet_tvar_20[5].delimiter[7] );
tran (\_zy_simnet_tvar_20[5][6] , \_zy_simnet_tvar_20[5].delimiter[6] );
tran (\_zy_simnet_tvar_20[5][5] , \_zy_simnet_tvar_20[5].delimiter[5] );
tran (\_zy_simnet_tvar_20[5][4] , \_zy_simnet_tvar_20[5].delimiter[4] );
tran (\_zy_simnet_tvar_20[5][3] , \_zy_simnet_tvar_20[5].delimiter[3] );
tran (\_zy_simnet_tvar_20[5][2] , \_zy_simnet_tvar_20[5].delimiter[2] );
tran (\_zy_simnet_tvar_20[5][1] , \_zy_simnet_tvar_20[5].delimiter[1] );
tran (\_zy_simnet_tvar_20[5][0] , \_zy_simnet_tvar_20[5].delimiter[0] );
tran (\_zy_simnet_tvar_20[4][271] , \_zy_simnet_tvar_20[4].guid_size[0] );
tran (\_zy_simnet_tvar_20[4][270] , \_zy_simnet_tvar_20[4].label_size[5] );
tran (\_zy_simnet_tvar_20[4][269] , \_zy_simnet_tvar_20[4].label_size[4] );
tran (\_zy_simnet_tvar_20[4][268] , \_zy_simnet_tvar_20[4].label_size[3] );
tran (\_zy_simnet_tvar_20[4][267] , \_zy_simnet_tvar_20[4].label_size[2] );
tran (\_zy_simnet_tvar_20[4][266] , \_zy_simnet_tvar_20[4].label_size[1] );
tran (\_zy_simnet_tvar_20[4][265] , \_zy_simnet_tvar_20[4].label_size[0] );
tran (\_zy_simnet_tvar_20[4][264] , \_zy_simnet_tvar_20[4].label[255] );
tran (\_zy_simnet_tvar_20[4][263] , \_zy_simnet_tvar_20[4].label[254] );
tran (\_zy_simnet_tvar_20[4][262] , \_zy_simnet_tvar_20[4].label[253] );
tran (\_zy_simnet_tvar_20[4][261] , \_zy_simnet_tvar_20[4].label[252] );
tran (\_zy_simnet_tvar_20[4][260] , \_zy_simnet_tvar_20[4].label[251] );
tran (\_zy_simnet_tvar_20[4][259] , \_zy_simnet_tvar_20[4].label[250] );
tran (\_zy_simnet_tvar_20[4][258] , \_zy_simnet_tvar_20[4].label[249] );
tran (\_zy_simnet_tvar_20[4][257] , \_zy_simnet_tvar_20[4].label[248] );
tran (\_zy_simnet_tvar_20[4][256] , \_zy_simnet_tvar_20[4].label[247] );
tran (\_zy_simnet_tvar_20[4][255] , \_zy_simnet_tvar_20[4].label[246] );
tran (\_zy_simnet_tvar_20[4][254] , \_zy_simnet_tvar_20[4].label[245] );
tran (\_zy_simnet_tvar_20[4][253] , \_zy_simnet_tvar_20[4].label[244] );
tran (\_zy_simnet_tvar_20[4][252] , \_zy_simnet_tvar_20[4].label[243] );
tran (\_zy_simnet_tvar_20[4][251] , \_zy_simnet_tvar_20[4].label[242] );
tran (\_zy_simnet_tvar_20[4][250] , \_zy_simnet_tvar_20[4].label[241] );
tran (\_zy_simnet_tvar_20[4][249] , \_zy_simnet_tvar_20[4].label[240] );
tran (\_zy_simnet_tvar_20[4][248] , \_zy_simnet_tvar_20[4].label[239] );
tran (\_zy_simnet_tvar_20[4][247] , \_zy_simnet_tvar_20[4].label[238] );
tran (\_zy_simnet_tvar_20[4][246] , \_zy_simnet_tvar_20[4].label[237] );
tran (\_zy_simnet_tvar_20[4][245] , \_zy_simnet_tvar_20[4].label[236] );
tran (\_zy_simnet_tvar_20[4][244] , \_zy_simnet_tvar_20[4].label[235] );
tran (\_zy_simnet_tvar_20[4][243] , \_zy_simnet_tvar_20[4].label[234] );
tran (\_zy_simnet_tvar_20[4][242] , \_zy_simnet_tvar_20[4].label[233] );
tran (\_zy_simnet_tvar_20[4][241] , \_zy_simnet_tvar_20[4].label[232] );
tran (\_zy_simnet_tvar_20[4][240] , \_zy_simnet_tvar_20[4].label[231] );
tran (\_zy_simnet_tvar_20[4][239] , \_zy_simnet_tvar_20[4].label[230] );
tran (\_zy_simnet_tvar_20[4][238] , \_zy_simnet_tvar_20[4].label[229] );
tran (\_zy_simnet_tvar_20[4][237] , \_zy_simnet_tvar_20[4].label[228] );
tran (\_zy_simnet_tvar_20[4][236] , \_zy_simnet_tvar_20[4].label[227] );
tran (\_zy_simnet_tvar_20[4][235] , \_zy_simnet_tvar_20[4].label[226] );
tran (\_zy_simnet_tvar_20[4][234] , \_zy_simnet_tvar_20[4].label[225] );
tran (\_zy_simnet_tvar_20[4][233] , \_zy_simnet_tvar_20[4].label[224] );
tran (\_zy_simnet_tvar_20[4][232] , \_zy_simnet_tvar_20[4].label[223] );
tran (\_zy_simnet_tvar_20[4][231] , \_zy_simnet_tvar_20[4].label[222] );
tran (\_zy_simnet_tvar_20[4][230] , \_zy_simnet_tvar_20[4].label[221] );
tran (\_zy_simnet_tvar_20[4][229] , \_zy_simnet_tvar_20[4].label[220] );
tran (\_zy_simnet_tvar_20[4][228] , \_zy_simnet_tvar_20[4].label[219] );
tran (\_zy_simnet_tvar_20[4][227] , \_zy_simnet_tvar_20[4].label[218] );
tran (\_zy_simnet_tvar_20[4][226] , \_zy_simnet_tvar_20[4].label[217] );
tran (\_zy_simnet_tvar_20[4][225] , \_zy_simnet_tvar_20[4].label[216] );
tran (\_zy_simnet_tvar_20[4][224] , \_zy_simnet_tvar_20[4].label[215] );
tran (\_zy_simnet_tvar_20[4][223] , \_zy_simnet_tvar_20[4].label[214] );
tran (\_zy_simnet_tvar_20[4][222] , \_zy_simnet_tvar_20[4].label[213] );
tran (\_zy_simnet_tvar_20[4][221] , \_zy_simnet_tvar_20[4].label[212] );
tran (\_zy_simnet_tvar_20[4][220] , \_zy_simnet_tvar_20[4].label[211] );
tran (\_zy_simnet_tvar_20[4][219] , \_zy_simnet_tvar_20[4].label[210] );
tran (\_zy_simnet_tvar_20[4][218] , \_zy_simnet_tvar_20[4].label[209] );
tran (\_zy_simnet_tvar_20[4][217] , \_zy_simnet_tvar_20[4].label[208] );
tran (\_zy_simnet_tvar_20[4][216] , \_zy_simnet_tvar_20[4].label[207] );
tran (\_zy_simnet_tvar_20[4][215] , \_zy_simnet_tvar_20[4].label[206] );
tran (\_zy_simnet_tvar_20[4][214] , \_zy_simnet_tvar_20[4].label[205] );
tran (\_zy_simnet_tvar_20[4][213] , \_zy_simnet_tvar_20[4].label[204] );
tran (\_zy_simnet_tvar_20[4][212] , \_zy_simnet_tvar_20[4].label[203] );
tran (\_zy_simnet_tvar_20[4][211] , \_zy_simnet_tvar_20[4].label[202] );
tran (\_zy_simnet_tvar_20[4][210] , \_zy_simnet_tvar_20[4].label[201] );
tran (\_zy_simnet_tvar_20[4][209] , \_zy_simnet_tvar_20[4].label[200] );
tran (\_zy_simnet_tvar_20[4][208] , \_zy_simnet_tvar_20[4].label[199] );
tran (\_zy_simnet_tvar_20[4][207] , \_zy_simnet_tvar_20[4].label[198] );
tran (\_zy_simnet_tvar_20[4][206] , \_zy_simnet_tvar_20[4].label[197] );
tran (\_zy_simnet_tvar_20[4][205] , \_zy_simnet_tvar_20[4].label[196] );
tran (\_zy_simnet_tvar_20[4][204] , \_zy_simnet_tvar_20[4].label[195] );
tran (\_zy_simnet_tvar_20[4][203] , \_zy_simnet_tvar_20[4].label[194] );
tran (\_zy_simnet_tvar_20[4][202] , \_zy_simnet_tvar_20[4].label[193] );
tran (\_zy_simnet_tvar_20[4][201] , \_zy_simnet_tvar_20[4].label[192] );
tran (\_zy_simnet_tvar_20[4][200] , \_zy_simnet_tvar_20[4].label[191] );
tran (\_zy_simnet_tvar_20[4][199] , \_zy_simnet_tvar_20[4].label[190] );
tran (\_zy_simnet_tvar_20[4][198] , \_zy_simnet_tvar_20[4].label[189] );
tran (\_zy_simnet_tvar_20[4][197] , \_zy_simnet_tvar_20[4].label[188] );
tran (\_zy_simnet_tvar_20[4][196] , \_zy_simnet_tvar_20[4].label[187] );
tran (\_zy_simnet_tvar_20[4][195] , \_zy_simnet_tvar_20[4].label[186] );
tran (\_zy_simnet_tvar_20[4][194] , \_zy_simnet_tvar_20[4].label[185] );
tran (\_zy_simnet_tvar_20[4][193] , \_zy_simnet_tvar_20[4].label[184] );
tran (\_zy_simnet_tvar_20[4][192] , \_zy_simnet_tvar_20[4].label[183] );
tran (\_zy_simnet_tvar_20[4][191] , \_zy_simnet_tvar_20[4].label[182] );
tran (\_zy_simnet_tvar_20[4][190] , \_zy_simnet_tvar_20[4].label[181] );
tran (\_zy_simnet_tvar_20[4][189] , \_zy_simnet_tvar_20[4].label[180] );
tran (\_zy_simnet_tvar_20[4][188] , \_zy_simnet_tvar_20[4].label[179] );
tran (\_zy_simnet_tvar_20[4][187] , \_zy_simnet_tvar_20[4].label[178] );
tran (\_zy_simnet_tvar_20[4][186] , \_zy_simnet_tvar_20[4].label[177] );
tran (\_zy_simnet_tvar_20[4][185] , \_zy_simnet_tvar_20[4].label[176] );
tran (\_zy_simnet_tvar_20[4][184] , \_zy_simnet_tvar_20[4].label[175] );
tran (\_zy_simnet_tvar_20[4][183] , \_zy_simnet_tvar_20[4].label[174] );
tran (\_zy_simnet_tvar_20[4][182] , \_zy_simnet_tvar_20[4].label[173] );
tran (\_zy_simnet_tvar_20[4][181] , \_zy_simnet_tvar_20[4].label[172] );
tran (\_zy_simnet_tvar_20[4][180] , \_zy_simnet_tvar_20[4].label[171] );
tran (\_zy_simnet_tvar_20[4][179] , \_zy_simnet_tvar_20[4].label[170] );
tran (\_zy_simnet_tvar_20[4][178] , \_zy_simnet_tvar_20[4].label[169] );
tran (\_zy_simnet_tvar_20[4][177] , \_zy_simnet_tvar_20[4].label[168] );
tran (\_zy_simnet_tvar_20[4][176] , \_zy_simnet_tvar_20[4].label[167] );
tran (\_zy_simnet_tvar_20[4][175] , \_zy_simnet_tvar_20[4].label[166] );
tran (\_zy_simnet_tvar_20[4][174] , \_zy_simnet_tvar_20[4].label[165] );
tran (\_zy_simnet_tvar_20[4][173] , \_zy_simnet_tvar_20[4].label[164] );
tran (\_zy_simnet_tvar_20[4][172] , \_zy_simnet_tvar_20[4].label[163] );
tran (\_zy_simnet_tvar_20[4][171] , \_zy_simnet_tvar_20[4].label[162] );
tran (\_zy_simnet_tvar_20[4][170] , \_zy_simnet_tvar_20[4].label[161] );
tran (\_zy_simnet_tvar_20[4][169] , \_zy_simnet_tvar_20[4].label[160] );
tran (\_zy_simnet_tvar_20[4][168] , \_zy_simnet_tvar_20[4].label[159] );
tran (\_zy_simnet_tvar_20[4][167] , \_zy_simnet_tvar_20[4].label[158] );
tran (\_zy_simnet_tvar_20[4][166] , \_zy_simnet_tvar_20[4].label[157] );
tran (\_zy_simnet_tvar_20[4][165] , \_zy_simnet_tvar_20[4].label[156] );
tran (\_zy_simnet_tvar_20[4][164] , \_zy_simnet_tvar_20[4].label[155] );
tran (\_zy_simnet_tvar_20[4][163] , \_zy_simnet_tvar_20[4].label[154] );
tran (\_zy_simnet_tvar_20[4][162] , \_zy_simnet_tvar_20[4].label[153] );
tran (\_zy_simnet_tvar_20[4][161] , \_zy_simnet_tvar_20[4].label[152] );
tran (\_zy_simnet_tvar_20[4][160] , \_zy_simnet_tvar_20[4].label[151] );
tran (\_zy_simnet_tvar_20[4][159] , \_zy_simnet_tvar_20[4].label[150] );
tran (\_zy_simnet_tvar_20[4][158] , \_zy_simnet_tvar_20[4].label[149] );
tran (\_zy_simnet_tvar_20[4][157] , \_zy_simnet_tvar_20[4].label[148] );
tran (\_zy_simnet_tvar_20[4][156] , \_zy_simnet_tvar_20[4].label[147] );
tran (\_zy_simnet_tvar_20[4][155] , \_zy_simnet_tvar_20[4].label[146] );
tran (\_zy_simnet_tvar_20[4][154] , \_zy_simnet_tvar_20[4].label[145] );
tran (\_zy_simnet_tvar_20[4][153] , \_zy_simnet_tvar_20[4].label[144] );
tran (\_zy_simnet_tvar_20[4][152] , \_zy_simnet_tvar_20[4].label[143] );
tran (\_zy_simnet_tvar_20[4][151] , \_zy_simnet_tvar_20[4].label[142] );
tran (\_zy_simnet_tvar_20[4][150] , \_zy_simnet_tvar_20[4].label[141] );
tran (\_zy_simnet_tvar_20[4][149] , \_zy_simnet_tvar_20[4].label[140] );
tran (\_zy_simnet_tvar_20[4][148] , \_zy_simnet_tvar_20[4].label[139] );
tran (\_zy_simnet_tvar_20[4][147] , \_zy_simnet_tvar_20[4].label[138] );
tran (\_zy_simnet_tvar_20[4][146] , \_zy_simnet_tvar_20[4].label[137] );
tran (\_zy_simnet_tvar_20[4][145] , \_zy_simnet_tvar_20[4].label[136] );
tran (\_zy_simnet_tvar_20[4][144] , \_zy_simnet_tvar_20[4].label[135] );
tran (\_zy_simnet_tvar_20[4][143] , \_zy_simnet_tvar_20[4].label[134] );
tran (\_zy_simnet_tvar_20[4][142] , \_zy_simnet_tvar_20[4].label[133] );
tran (\_zy_simnet_tvar_20[4][141] , \_zy_simnet_tvar_20[4].label[132] );
tran (\_zy_simnet_tvar_20[4][140] , \_zy_simnet_tvar_20[4].label[131] );
tran (\_zy_simnet_tvar_20[4][139] , \_zy_simnet_tvar_20[4].label[130] );
tran (\_zy_simnet_tvar_20[4][138] , \_zy_simnet_tvar_20[4].label[129] );
tran (\_zy_simnet_tvar_20[4][137] , \_zy_simnet_tvar_20[4].label[128] );
tran (\_zy_simnet_tvar_20[4][136] , \_zy_simnet_tvar_20[4].label[127] );
tran (\_zy_simnet_tvar_20[4][135] , \_zy_simnet_tvar_20[4].label[126] );
tran (\_zy_simnet_tvar_20[4][134] , \_zy_simnet_tvar_20[4].label[125] );
tran (\_zy_simnet_tvar_20[4][133] , \_zy_simnet_tvar_20[4].label[124] );
tran (\_zy_simnet_tvar_20[4][132] , \_zy_simnet_tvar_20[4].label[123] );
tran (\_zy_simnet_tvar_20[4][131] , \_zy_simnet_tvar_20[4].label[122] );
tran (\_zy_simnet_tvar_20[4][130] , \_zy_simnet_tvar_20[4].label[121] );
tran (\_zy_simnet_tvar_20[4][129] , \_zy_simnet_tvar_20[4].label[120] );
tran (\_zy_simnet_tvar_20[4][128] , \_zy_simnet_tvar_20[4].label[119] );
tran (\_zy_simnet_tvar_20[4][127] , \_zy_simnet_tvar_20[4].label[118] );
tran (\_zy_simnet_tvar_20[4][126] , \_zy_simnet_tvar_20[4].label[117] );
tran (\_zy_simnet_tvar_20[4][125] , \_zy_simnet_tvar_20[4].label[116] );
tran (\_zy_simnet_tvar_20[4][124] , \_zy_simnet_tvar_20[4].label[115] );
tran (\_zy_simnet_tvar_20[4][123] , \_zy_simnet_tvar_20[4].label[114] );
tran (\_zy_simnet_tvar_20[4][122] , \_zy_simnet_tvar_20[4].label[113] );
tran (\_zy_simnet_tvar_20[4][121] , \_zy_simnet_tvar_20[4].label[112] );
tran (\_zy_simnet_tvar_20[4][120] , \_zy_simnet_tvar_20[4].label[111] );
tran (\_zy_simnet_tvar_20[4][119] , \_zy_simnet_tvar_20[4].label[110] );
tran (\_zy_simnet_tvar_20[4][118] , \_zy_simnet_tvar_20[4].label[109] );
tran (\_zy_simnet_tvar_20[4][117] , \_zy_simnet_tvar_20[4].label[108] );
tran (\_zy_simnet_tvar_20[4][116] , \_zy_simnet_tvar_20[4].label[107] );
tran (\_zy_simnet_tvar_20[4][115] , \_zy_simnet_tvar_20[4].label[106] );
tran (\_zy_simnet_tvar_20[4][114] , \_zy_simnet_tvar_20[4].label[105] );
tran (\_zy_simnet_tvar_20[4][113] , \_zy_simnet_tvar_20[4].label[104] );
tran (\_zy_simnet_tvar_20[4][112] , \_zy_simnet_tvar_20[4].label[103] );
tran (\_zy_simnet_tvar_20[4][111] , \_zy_simnet_tvar_20[4].label[102] );
tran (\_zy_simnet_tvar_20[4][110] , \_zy_simnet_tvar_20[4].label[101] );
tran (\_zy_simnet_tvar_20[4][109] , \_zy_simnet_tvar_20[4].label[100] );
tran (\_zy_simnet_tvar_20[4][108] , \_zy_simnet_tvar_20[4].label[99] );
tran (\_zy_simnet_tvar_20[4][107] , \_zy_simnet_tvar_20[4].label[98] );
tran (\_zy_simnet_tvar_20[4][106] , \_zy_simnet_tvar_20[4].label[97] );
tran (\_zy_simnet_tvar_20[4][105] , \_zy_simnet_tvar_20[4].label[96] );
tran (\_zy_simnet_tvar_20[4][104] , \_zy_simnet_tvar_20[4].label[95] );
tran (\_zy_simnet_tvar_20[4][103] , \_zy_simnet_tvar_20[4].label[94] );
tran (\_zy_simnet_tvar_20[4][102] , \_zy_simnet_tvar_20[4].label[93] );
tran (\_zy_simnet_tvar_20[4][101] , \_zy_simnet_tvar_20[4].label[92] );
tran (\_zy_simnet_tvar_20[4][100] , \_zy_simnet_tvar_20[4].label[91] );
tran (\_zy_simnet_tvar_20[4][99] , \_zy_simnet_tvar_20[4].label[90] );
tran (\_zy_simnet_tvar_20[4][98] , \_zy_simnet_tvar_20[4].label[89] );
tran (\_zy_simnet_tvar_20[4][97] , \_zy_simnet_tvar_20[4].label[88] );
tran (\_zy_simnet_tvar_20[4][96] , \_zy_simnet_tvar_20[4].label[87] );
tran (\_zy_simnet_tvar_20[4][95] , \_zy_simnet_tvar_20[4].label[86] );
tran (\_zy_simnet_tvar_20[4][94] , \_zy_simnet_tvar_20[4].label[85] );
tran (\_zy_simnet_tvar_20[4][93] , \_zy_simnet_tvar_20[4].label[84] );
tran (\_zy_simnet_tvar_20[4][92] , \_zy_simnet_tvar_20[4].label[83] );
tran (\_zy_simnet_tvar_20[4][91] , \_zy_simnet_tvar_20[4].label[82] );
tran (\_zy_simnet_tvar_20[4][90] , \_zy_simnet_tvar_20[4].label[81] );
tran (\_zy_simnet_tvar_20[4][89] , \_zy_simnet_tvar_20[4].label[80] );
tran (\_zy_simnet_tvar_20[4][88] , \_zy_simnet_tvar_20[4].label[79] );
tran (\_zy_simnet_tvar_20[4][87] , \_zy_simnet_tvar_20[4].label[78] );
tran (\_zy_simnet_tvar_20[4][86] , \_zy_simnet_tvar_20[4].label[77] );
tran (\_zy_simnet_tvar_20[4][85] , \_zy_simnet_tvar_20[4].label[76] );
tran (\_zy_simnet_tvar_20[4][84] , \_zy_simnet_tvar_20[4].label[75] );
tran (\_zy_simnet_tvar_20[4][83] , \_zy_simnet_tvar_20[4].label[74] );
tran (\_zy_simnet_tvar_20[4][82] , \_zy_simnet_tvar_20[4].label[73] );
tran (\_zy_simnet_tvar_20[4][81] , \_zy_simnet_tvar_20[4].label[72] );
tran (\_zy_simnet_tvar_20[4][80] , \_zy_simnet_tvar_20[4].label[71] );
tran (\_zy_simnet_tvar_20[4][79] , \_zy_simnet_tvar_20[4].label[70] );
tran (\_zy_simnet_tvar_20[4][78] , \_zy_simnet_tvar_20[4].label[69] );
tran (\_zy_simnet_tvar_20[4][77] , \_zy_simnet_tvar_20[4].label[68] );
tran (\_zy_simnet_tvar_20[4][76] , \_zy_simnet_tvar_20[4].label[67] );
tran (\_zy_simnet_tvar_20[4][75] , \_zy_simnet_tvar_20[4].label[66] );
tran (\_zy_simnet_tvar_20[4][74] , \_zy_simnet_tvar_20[4].label[65] );
tran (\_zy_simnet_tvar_20[4][73] , \_zy_simnet_tvar_20[4].label[64] );
tran (\_zy_simnet_tvar_20[4][72] , \_zy_simnet_tvar_20[4].label[63] );
tran (\_zy_simnet_tvar_20[4][71] , \_zy_simnet_tvar_20[4].label[62] );
tran (\_zy_simnet_tvar_20[4][70] , \_zy_simnet_tvar_20[4].label[61] );
tran (\_zy_simnet_tvar_20[4][69] , \_zy_simnet_tvar_20[4].label[60] );
tran (\_zy_simnet_tvar_20[4][68] , \_zy_simnet_tvar_20[4].label[59] );
tran (\_zy_simnet_tvar_20[4][67] , \_zy_simnet_tvar_20[4].label[58] );
tran (\_zy_simnet_tvar_20[4][66] , \_zy_simnet_tvar_20[4].label[57] );
tran (\_zy_simnet_tvar_20[4][65] , \_zy_simnet_tvar_20[4].label[56] );
tran (\_zy_simnet_tvar_20[4][64] , \_zy_simnet_tvar_20[4].label[55] );
tran (\_zy_simnet_tvar_20[4][63] , \_zy_simnet_tvar_20[4].label[54] );
tran (\_zy_simnet_tvar_20[4][62] , \_zy_simnet_tvar_20[4].label[53] );
tran (\_zy_simnet_tvar_20[4][61] , \_zy_simnet_tvar_20[4].label[52] );
tran (\_zy_simnet_tvar_20[4][60] , \_zy_simnet_tvar_20[4].label[51] );
tran (\_zy_simnet_tvar_20[4][59] , \_zy_simnet_tvar_20[4].label[50] );
tran (\_zy_simnet_tvar_20[4][58] , \_zy_simnet_tvar_20[4].label[49] );
tran (\_zy_simnet_tvar_20[4][57] , \_zy_simnet_tvar_20[4].label[48] );
tran (\_zy_simnet_tvar_20[4][56] , \_zy_simnet_tvar_20[4].label[47] );
tran (\_zy_simnet_tvar_20[4][55] , \_zy_simnet_tvar_20[4].label[46] );
tran (\_zy_simnet_tvar_20[4][54] , \_zy_simnet_tvar_20[4].label[45] );
tran (\_zy_simnet_tvar_20[4][53] , \_zy_simnet_tvar_20[4].label[44] );
tran (\_zy_simnet_tvar_20[4][52] , \_zy_simnet_tvar_20[4].label[43] );
tran (\_zy_simnet_tvar_20[4][51] , \_zy_simnet_tvar_20[4].label[42] );
tran (\_zy_simnet_tvar_20[4][50] , \_zy_simnet_tvar_20[4].label[41] );
tran (\_zy_simnet_tvar_20[4][49] , \_zy_simnet_tvar_20[4].label[40] );
tran (\_zy_simnet_tvar_20[4][48] , \_zy_simnet_tvar_20[4].label[39] );
tran (\_zy_simnet_tvar_20[4][47] , \_zy_simnet_tvar_20[4].label[38] );
tran (\_zy_simnet_tvar_20[4][46] , \_zy_simnet_tvar_20[4].label[37] );
tran (\_zy_simnet_tvar_20[4][45] , \_zy_simnet_tvar_20[4].label[36] );
tran (\_zy_simnet_tvar_20[4][44] , \_zy_simnet_tvar_20[4].label[35] );
tran (\_zy_simnet_tvar_20[4][43] , \_zy_simnet_tvar_20[4].label[34] );
tran (\_zy_simnet_tvar_20[4][42] , \_zy_simnet_tvar_20[4].label[33] );
tran (\_zy_simnet_tvar_20[4][41] , \_zy_simnet_tvar_20[4].label[32] );
tran (\_zy_simnet_tvar_20[4][40] , \_zy_simnet_tvar_20[4].label[31] );
tran (\_zy_simnet_tvar_20[4][39] , \_zy_simnet_tvar_20[4].label[30] );
tran (\_zy_simnet_tvar_20[4][38] , \_zy_simnet_tvar_20[4].label[29] );
tran (\_zy_simnet_tvar_20[4][37] , \_zy_simnet_tvar_20[4].label[28] );
tran (\_zy_simnet_tvar_20[4][36] , \_zy_simnet_tvar_20[4].label[27] );
tran (\_zy_simnet_tvar_20[4][35] , \_zy_simnet_tvar_20[4].label[26] );
tran (\_zy_simnet_tvar_20[4][34] , \_zy_simnet_tvar_20[4].label[25] );
tran (\_zy_simnet_tvar_20[4][33] , \_zy_simnet_tvar_20[4].label[24] );
tran (\_zy_simnet_tvar_20[4][32] , \_zy_simnet_tvar_20[4].label[23] );
tran (\_zy_simnet_tvar_20[4][31] , \_zy_simnet_tvar_20[4].label[22] );
tran (\_zy_simnet_tvar_20[4][30] , \_zy_simnet_tvar_20[4].label[21] );
tran (\_zy_simnet_tvar_20[4][29] , \_zy_simnet_tvar_20[4].label[20] );
tran (\_zy_simnet_tvar_20[4][28] , \_zy_simnet_tvar_20[4].label[19] );
tran (\_zy_simnet_tvar_20[4][27] , \_zy_simnet_tvar_20[4].label[18] );
tran (\_zy_simnet_tvar_20[4][26] , \_zy_simnet_tvar_20[4].label[17] );
tran (\_zy_simnet_tvar_20[4][25] , \_zy_simnet_tvar_20[4].label[16] );
tran (\_zy_simnet_tvar_20[4][24] , \_zy_simnet_tvar_20[4].label[15] );
tran (\_zy_simnet_tvar_20[4][23] , \_zy_simnet_tvar_20[4].label[14] );
tran (\_zy_simnet_tvar_20[4][22] , \_zy_simnet_tvar_20[4].label[13] );
tran (\_zy_simnet_tvar_20[4][21] , \_zy_simnet_tvar_20[4].label[12] );
tran (\_zy_simnet_tvar_20[4][20] , \_zy_simnet_tvar_20[4].label[11] );
tran (\_zy_simnet_tvar_20[4][19] , \_zy_simnet_tvar_20[4].label[10] );
tran (\_zy_simnet_tvar_20[4][18] , \_zy_simnet_tvar_20[4].label[9] );
tran (\_zy_simnet_tvar_20[4][17] , \_zy_simnet_tvar_20[4].label[8] );
tran (\_zy_simnet_tvar_20[4][16] , \_zy_simnet_tvar_20[4].label[7] );
tran (\_zy_simnet_tvar_20[4][15] , \_zy_simnet_tvar_20[4].label[6] );
tran (\_zy_simnet_tvar_20[4][14] , \_zy_simnet_tvar_20[4].label[5] );
tran (\_zy_simnet_tvar_20[4][13] , \_zy_simnet_tvar_20[4].label[4] );
tran (\_zy_simnet_tvar_20[4][12] , \_zy_simnet_tvar_20[4].label[3] );
tran (\_zy_simnet_tvar_20[4][11] , \_zy_simnet_tvar_20[4].label[2] );
tran (\_zy_simnet_tvar_20[4][10] , \_zy_simnet_tvar_20[4].label[1] );
tran (\_zy_simnet_tvar_20[4][9] , \_zy_simnet_tvar_20[4].label[0] );
tran (\_zy_simnet_tvar_20[4][8] , \_zy_simnet_tvar_20[4].delimiter_valid[0] );
tran (\_zy_simnet_tvar_20[4][7] , \_zy_simnet_tvar_20[4].delimiter[7] );
tran (\_zy_simnet_tvar_20[4][6] , \_zy_simnet_tvar_20[4].delimiter[6] );
tran (\_zy_simnet_tvar_20[4][5] , \_zy_simnet_tvar_20[4].delimiter[5] );
tran (\_zy_simnet_tvar_20[4][4] , \_zy_simnet_tvar_20[4].delimiter[4] );
tran (\_zy_simnet_tvar_20[4][3] , \_zy_simnet_tvar_20[4].delimiter[3] );
tran (\_zy_simnet_tvar_20[4][2] , \_zy_simnet_tvar_20[4].delimiter[2] );
tran (\_zy_simnet_tvar_20[4][1] , \_zy_simnet_tvar_20[4].delimiter[1] );
tran (\_zy_simnet_tvar_20[4][0] , \_zy_simnet_tvar_20[4].delimiter[0] );
tran (\_zy_simnet_tvar_20[3][271] , \_zy_simnet_tvar_20[3].guid_size[0] );
tran (\_zy_simnet_tvar_20[3][270] , \_zy_simnet_tvar_20[3].label_size[5] );
tran (\_zy_simnet_tvar_20[3][269] , \_zy_simnet_tvar_20[3].label_size[4] );
tran (\_zy_simnet_tvar_20[3][268] , \_zy_simnet_tvar_20[3].label_size[3] );
tran (\_zy_simnet_tvar_20[3][267] , \_zy_simnet_tvar_20[3].label_size[2] );
tran (\_zy_simnet_tvar_20[3][266] , \_zy_simnet_tvar_20[3].label_size[1] );
tran (\_zy_simnet_tvar_20[3][265] , \_zy_simnet_tvar_20[3].label_size[0] );
tran (\_zy_simnet_tvar_20[3][264] , \_zy_simnet_tvar_20[3].label[255] );
tran (\_zy_simnet_tvar_20[3][263] , \_zy_simnet_tvar_20[3].label[254] );
tran (\_zy_simnet_tvar_20[3][262] , \_zy_simnet_tvar_20[3].label[253] );
tran (\_zy_simnet_tvar_20[3][261] , \_zy_simnet_tvar_20[3].label[252] );
tran (\_zy_simnet_tvar_20[3][260] , \_zy_simnet_tvar_20[3].label[251] );
tran (\_zy_simnet_tvar_20[3][259] , \_zy_simnet_tvar_20[3].label[250] );
tran (\_zy_simnet_tvar_20[3][258] , \_zy_simnet_tvar_20[3].label[249] );
tran (\_zy_simnet_tvar_20[3][257] , \_zy_simnet_tvar_20[3].label[248] );
tran (\_zy_simnet_tvar_20[3][256] , \_zy_simnet_tvar_20[3].label[247] );
tran (\_zy_simnet_tvar_20[3][255] , \_zy_simnet_tvar_20[3].label[246] );
tran (\_zy_simnet_tvar_20[3][254] , \_zy_simnet_tvar_20[3].label[245] );
tran (\_zy_simnet_tvar_20[3][253] , \_zy_simnet_tvar_20[3].label[244] );
tran (\_zy_simnet_tvar_20[3][252] , \_zy_simnet_tvar_20[3].label[243] );
tran (\_zy_simnet_tvar_20[3][251] , \_zy_simnet_tvar_20[3].label[242] );
tran (\_zy_simnet_tvar_20[3][250] , \_zy_simnet_tvar_20[3].label[241] );
tran (\_zy_simnet_tvar_20[3][249] , \_zy_simnet_tvar_20[3].label[240] );
tran (\_zy_simnet_tvar_20[3][248] , \_zy_simnet_tvar_20[3].label[239] );
tran (\_zy_simnet_tvar_20[3][247] , \_zy_simnet_tvar_20[3].label[238] );
tran (\_zy_simnet_tvar_20[3][246] , \_zy_simnet_tvar_20[3].label[237] );
tran (\_zy_simnet_tvar_20[3][245] , \_zy_simnet_tvar_20[3].label[236] );
tran (\_zy_simnet_tvar_20[3][244] , \_zy_simnet_tvar_20[3].label[235] );
tran (\_zy_simnet_tvar_20[3][243] , \_zy_simnet_tvar_20[3].label[234] );
tran (\_zy_simnet_tvar_20[3][242] , \_zy_simnet_tvar_20[3].label[233] );
tran (\_zy_simnet_tvar_20[3][241] , \_zy_simnet_tvar_20[3].label[232] );
tran (\_zy_simnet_tvar_20[3][240] , \_zy_simnet_tvar_20[3].label[231] );
tran (\_zy_simnet_tvar_20[3][239] , \_zy_simnet_tvar_20[3].label[230] );
tran (\_zy_simnet_tvar_20[3][238] , \_zy_simnet_tvar_20[3].label[229] );
tran (\_zy_simnet_tvar_20[3][237] , \_zy_simnet_tvar_20[3].label[228] );
tran (\_zy_simnet_tvar_20[3][236] , \_zy_simnet_tvar_20[3].label[227] );
tran (\_zy_simnet_tvar_20[3][235] , \_zy_simnet_tvar_20[3].label[226] );
tran (\_zy_simnet_tvar_20[3][234] , \_zy_simnet_tvar_20[3].label[225] );
tran (\_zy_simnet_tvar_20[3][233] , \_zy_simnet_tvar_20[3].label[224] );
tran (\_zy_simnet_tvar_20[3][232] , \_zy_simnet_tvar_20[3].label[223] );
tran (\_zy_simnet_tvar_20[3][231] , \_zy_simnet_tvar_20[3].label[222] );
tran (\_zy_simnet_tvar_20[3][230] , \_zy_simnet_tvar_20[3].label[221] );
tran (\_zy_simnet_tvar_20[3][229] , \_zy_simnet_tvar_20[3].label[220] );
tran (\_zy_simnet_tvar_20[3][228] , \_zy_simnet_tvar_20[3].label[219] );
tran (\_zy_simnet_tvar_20[3][227] , \_zy_simnet_tvar_20[3].label[218] );
tran (\_zy_simnet_tvar_20[3][226] , \_zy_simnet_tvar_20[3].label[217] );
tran (\_zy_simnet_tvar_20[3][225] , \_zy_simnet_tvar_20[3].label[216] );
tran (\_zy_simnet_tvar_20[3][224] , \_zy_simnet_tvar_20[3].label[215] );
tran (\_zy_simnet_tvar_20[3][223] , \_zy_simnet_tvar_20[3].label[214] );
tran (\_zy_simnet_tvar_20[3][222] , \_zy_simnet_tvar_20[3].label[213] );
tran (\_zy_simnet_tvar_20[3][221] , \_zy_simnet_tvar_20[3].label[212] );
tran (\_zy_simnet_tvar_20[3][220] , \_zy_simnet_tvar_20[3].label[211] );
tran (\_zy_simnet_tvar_20[3][219] , \_zy_simnet_tvar_20[3].label[210] );
tran (\_zy_simnet_tvar_20[3][218] , \_zy_simnet_tvar_20[3].label[209] );
tran (\_zy_simnet_tvar_20[3][217] , \_zy_simnet_tvar_20[3].label[208] );
tran (\_zy_simnet_tvar_20[3][216] , \_zy_simnet_tvar_20[3].label[207] );
tran (\_zy_simnet_tvar_20[3][215] , \_zy_simnet_tvar_20[3].label[206] );
tran (\_zy_simnet_tvar_20[3][214] , \_zy_simnet_tvar_20[3].label[205] );
tran (\_zy_simnet_tvar_20[3][213] , \_zy_simnet_tvar_20[3].label[204] );
tran (\_zy_simnet_tvar_20[3][212] , \_zy_simnet_tvar_20[3].label[203] );
tran (\_zy_simnet_tvar_20[3][211] , \_zy_simnet_tvar_20[3].label[202] );
tran (\_zy_simnet_tvar_20[3][210] , \_zy_simnet_tvar_20[3].label[201] );
tran (\_zy_simnet_tvar_20[3][209] , \_zy_simnet_tvar_20[3].label[200] );
tran (\_zy_simnet_tvar_20[3][208] , \_zy_simnet_tvar_20[3].label[199] );
tran (\_zy_simnet_tvar_20[3][207] , \_zy_simnet_tvar_20[3].label[198] );
tran (\_zy_simnet_tvar_20[3][206] , \_zy_simnet_tvar_20[3].label[197] );
tran (\_zy_simnet_tvar_20[3][205] , \_zy_simnet_tvar_20[3].label[196] );
tran (\_zy_simnet_tvar_20[3][204] , \_zy_simnet_tvar_20[3].label[195] );
tran (\_zy_simnet_tvar_20[3][203] , \_zy_simnet_tvar_20[3].label[194] );
tran (\_zy_simnet_tvar_20[3][202] , \_zy_simnet_tvar_20[3].label[193] );
tran (\_zy_simnet_tvar_20[3][201] , \_zy_simnet_tvar_20[3].label[192] );
tran (\_zy_simnet_tvar_20[3][200] , \_zy_simnet_tvar_20[3].label[191] );
tran (\_zy_simnet_tvar_20[3][199] , \_zy_simnet_tvar_20[3].label[190] );
tran (\_zy_simnet_tvar_20[3][198] , \_zy_simnet_tvar_20[3].label[189] );
tran (\_zy_simnet_tvar_20[3][197] , \_zy_simnet_tvar_20[3].label[188] );
tran (\_zy_simnet_tvar_20[3][196] , \_zy_simnet_tvar_20[3].label[187] );
tran (\_zy_simnet_tvar_20[3][195] , \_zy_simnet_tvar_20[3].label[186] );
tran (\_zy_simnet_tvar_20[3][194] , \_zy_simnet_tvar_20[3].label[185] );
tran (\_zy_simnet_tvar_20[3][193] , \_zy_simnet_tvar_20[3].label[184] );
tran (\_zy_simnet_tvar_20[3][192] , \_zy_simnet_tvar_20[3].label[183] );
tran (\_zy_simnet_tvar_20[3][191] , \_zy_simnet_tvar_20[3].label[182] );
tran (\_zy_simnet_tvar_20[3][190] , \_zy_simnet_tvar_20[3].label[181] );
tran (\_zy_simnet_tvar_20[3][189] , \_zy_simnet_tvar_20[3].label[180] );
tran (\_zy_simnet_tvar_20[3][188] , \_zy_simnet_tvar_20[3].label[179] );
tran (\_zy_simnet_tvar_20[3][187] , \_zy_simnet_tvar_20[3].label[178] );
tran (\_zy_simnet_tvar_20[3][186] , \_zy_simnet_tvar_20[3].label[177] );
tran (\_zy_simnet_tvar_20[3][185] , \_zy_simnet_tvar_20[3].label[176] );
tran (\_zy_simnet_tvar_20[3][184] , \_zy_simnet_tvar_20[3].label[175] );
tran (\_zy_simnet_tvar_20[3][183] , \_zy_simnet_tvar_20[3].label[174] );
tran (\_zy_simnet_tvar_20[3][182] , \_zy_simnet_tvar_20[3].label[173] );
tran (\_zy_simnet_tvar_20[3][181] , \_zy_simnet_tvar_20[3].label[172] );
tran (\_zy_simnet_tvar_20[3][180] , \_zy_simnet_tvar_20[3].label[171] );
tran (\_zy_simnet_tvar_20[3][179] , \_zy_simnet_tvar_20[3].label[170] );
tran (\_zy_simnet_tvar_20[3][178] , \_zy_simnet_tvar_20[3].label[169] );
tran (\_zy_simnet_tvar_20[3][177] , \_zy_simnet_tvar_20[3].label[168] );
tran (\_zy_simnet_tvar_20[3][176] , \_zy_simnet_tvar_20[3].label[167] );
tran (\_zy_simnet_tvar_20[3][175] , \_zy_simnet_tvar_20[3].label[166] );
tran (\_zy_simnet_tvar_20[3][174] , \_zy_simnet_tvar_20[3].label[165] );
tran (\_zy_simnet_tvar_20[3][173] , \_zy_simnet_tvar_20[3].label[164] );
tran (\_zy_simnet_tvar_20[3][172] , \_zy_simnet_tvar_20[3].label[163] );
tran (\_zy_simnet_tvar_20[3][171] , \_zy_simnet_tvar_20[3].label[162] );
tran (\_zy_simnet_tvar_20[3][170] , \_zy_simnet_tvar_20[3].label[161] );
tran (\_zy_simnet_tvar_20[3][169] , \_zy_simnet_tvar_20[3].label[160] );
tran (\_zy_simnet_tvar_20[3][168] , \_zy_simnet_tvar_20[3].label[159] );
tran (\_zy_simnet_tvar_20[3][167] , \_zy_simnet_tvar_20[3].label[158] );
tran (\_zy_simnet_tvar_20[3][166] , \_zy_simnet_tvar_20[3].label[157] );
tran (\_zy_simnet_tvar_20[3][165] , \_zy_simnet_tvar_20[3].label[156] );
tran (\_zy_simnet_tvar_20[3][164] , \_zy_simnet_tvar_20[3].label[155] );
tran (\_zy_simnet_tvar_20[3][163] , \_zy_simnet_tvar_20[3].label[154] );
tran (\_zy_simnet_tvar_20[3][162] , \_zy_simnet_tvar_20[3].label[153] );
tran (\_zy_simnet_tvar_20[3][161] , \_zy_simnet_tvar_20[3].label[152] );
tran (\_zy_simnet_tvar_20[3][160] , \_zy_simnet_tvar_20[3].label[151] );
tran (\_zy_simnet_tvar_20[3][159] , \_zy_simnet_tvar_20[3].label[150] );
tran (\_zy_simnet_tvar_20[3][158] , \_zy_simnet_tvar_20[3].label[149] );
tran (\_zy_simnet_tvar_20[3][157] , \_zy_simnet_tvar_20[3].label[148] );
tran (\_zy_simnet_tvar_20[3][156] , \_zy_simnet_tvar_20[3].label[147] );
tran (\_zy_simnet_tvar_20[3][155] , \_zy_simnet_tvar_20[3].label[146] );
tran (\_zy_simnet_tvar_20[3][154] , \_zy_simnet_tvar_20[3].label[145] );
tran (\_zy_simnet_tvar_20[3][153] , \_zy_simnet_tvar_20[3].label[144] );
tran (\_zy_simnet_tvar_20[3][152] , \_zy_simnet_tvar_20[3].label[143] );
tran (\_zy_simnet_tvar_20[3][151] , \_zy_simnet_tvar_20[3].label[142] );
tran (\_zy_simnet_tvar_20[3][150] , \_zy_simnet_tvar_20[3].label[141] );
tran (\_zy_simnet_tvar_20[3][149] , \_zy_simnet_tvar_20[3].label[140] );
tran (\_zy_simnet_tvar_20[3][148] , \_zy_simnet_tvar_20[3].label[139] );
tran (\_zy_simnet_tvar_20[3][147] , \_zy_simnet_tvar_20[3].label[138] );
tran (\_zy_simnet_tvar_20[3][146] , \_zy_simnet_tvar_20[3].label[137] );
tran (\_zy_simnet_tvar_20[3][145] , \_zy_simnet_tvar_20[3].label[136] );
tran (\_zy_simnet_tvar_20[3][144] , \_zy_simnet_tvar_20[3].label[135] );
tran (\_zy_simnet_tvar_20[3][143] , \_zy_simnet_tvar_20[3].label[134] );
tran (\_zy_simnet_tvar_20[3][142] , \_zy_simnet_tvar_20[3].label[133] );
tran (\_zy_simnet_tvar_20[3][141] , \_zy_simnet_tvar_20[3].label[132] );
tran (\_zy_simnet_tvar_20[3][140] , \_zy_simnet_tvar_20[3].label[131] );
tran (\_zy_simnet_tvar_20[3][139] , \_zy_simnet_tvar_20[3].label[130] );
tran (\_zy_simnet_tvar_20[3][138] , \_zy_simnet_tvar_20[3].label[129] );
tran (\_zy_simnet_tvar_20[3][137] , \_zy_simnet_tvar_20[3].label[128] );
tran (\_zy_simnet_tvar_20[3][136] , \_zy_simnet_tvar_20[3].label[127] );
tran (\_zy_simnet_tvar_20[3][135] , \_zy_simnet_tvar_20[3].label[126] );
tran (\_zy_simnet_tvar_20[3][134] , \_zy_simnet_tvar_20[3].label[125] );
tran (\_zy_simnet_tvar_20[3][133] , \_zy_simnet_tvar_20[3].label[124] );
tran (\_zy_simnet_tvar_20[3][132] , \_zy_simnet_tvar_20[3].label[123] );
tran (\_zy_simnet_tvar_20[3][131] , \_zy_simnet_tvar_20[3].label[122] );
tran (\_zy_simnet_tvar_20[3][130] , \_zy_simnet_tvar_20[3].label[121] );
tran (\_zy_simnet_tvar_20[3][129] , \_zy_simnet_tvar_20[3].label[120] );
tran (\_zy_simnet_tvar_20[3][128] , \_zy_simnet_tvar_20[3].label[119] );
tran (\_zy_simnet_tvar_20[3][127] , \_zy_simnet_tvar_20[3].label[118] );
tran (\_zy_simnet_tvar_20[3][126] , \_zy_simnet_tvar_20[3].label[117] );
tran (\_zy_simnet_tvar_20[3][125] , \_zy_simnet_tvar_20[3].label[116] );
tran (\_zy_simnet_tvar_20[3][124] , \_zy_simnet_tvar_20[3].label[115] );
tran (\_zy_simnet_tvar_20[3][123] , \_zy_simnet_tvar_20[3].label[114] );
tran (\_zy_simnet_tvar_20[3][122] , \_zy_simnet_tvar_20[3].label[113] );
tran (\_zy_simnet_tvar_20[3][121] , \_zy_simnet_tvar_20[3].label[112] );
tran (\_zy_simnet_tvar_20[3][120] , \_zy_simnet_tvar_20[3].label[111] );
tran (\_zy_simnet_tvar_20[3][119] , \_zy_simnet_tvar_20[3].label[110] );
tran (\_zy_simnet_tvar_20[3][118] , \_zy_simnet_tvar_20[3].label[109] );
tran (\_zy_simnet_tvar_20[3][117] , \_zy_simnet_tvar_20[3].label[108] );
tran (\_zy_simnet_tvar_20[3][116] , \_zy_simnet_tvar_20[3].label[107] );
tran (\_zy_simnet_tvar_20[3][115] , \_zy_simnet_tvar_20[3].label[106] );
tran (\_zy_simnet_tvar_20[3][114] , \_zy_simnet_tvar_20[3].label[105] );
tran (\_zy_simnet_tvar_20[3][113] , \_zy_simnet_tvar_20[3].label[104] );
tran (\_zy_simnet_tvar_20[3][112] , \_zy_simnet_tvar_20[3].label[103] );
tran (\_zy_simnet_tvar_20[3][111] , \_zy_simnet_tvar_20[3].label[102] );
tran (\_zy_simnet_tvar_20[3][110] , \_zy_simnet_tvar_20[3].label[101] );
tran (\_zy_simnet_tvar_20[3][109] , \_zy_simnet_tvar_20[3].label[100] );
tran (\_zy_simnet_tvar_20[3][108] , \_zy_simnet_tvar_20[3].label[99] );
tran (\_zy_simnet_tvar_20[3][107] , \_zy_simnet_tvar_20[3].label[98] );
tran (\_zy_simnet_tvar_20[3][106] , \_zy_simnet_tvar_20[3].label[97] );
tran (\_zy_simnet_tvar_20[3][105] , \_zy_simnet_tvar_20[3].label[96] );
tran (\_zy_simnet_tvar_20[3][104] , \_zy_simnet_tvar_20[3].label[95] );
tran (\_zy_simnet_tvar_20[3][103] , \_zy_simnet_tvar_20[3].label[94] );
tran (\_zy_simnet_tvar_20[3][102] , \_zy_simnet_tvar_20[3].label[93] );
tran (\_zy_simnet_tvar_20[3][101] , \_zy_simnet_tvar_20[3].label[92] );
tran (\_zy_simnet_tvar_20[3][100] , \_zy_simnet_tvar_20[3].label[91] );
tran (\_zy_simnet_tvar_20[3][99] , \_zy_simnet_tvar_20[3].label[90] );
tran (\_zy_simnet_tvar_20[3][98] , \_zy_simnet_tvar_20[3].label[89] );
tran (\_zy_simnet_tvar_20[3][97] , \_zy_simnet_tvar_20[3].label[88] );
tran (\_zy_simnet_tvar_20[3][96] , \_zy_simnet_tvar_20[3].label[87] );
tran (\_zy_simnet_tvar_20[3][95] , \_zy_simnet_tvar_20[3].label[86] );
tran (\_zy_simnet_tvar_20[3][94] , \_zy_simnet_tvar_20[3].label[85] );
tran (\_zy_simnet_tvar_20[3][93] , \_zy_simnet_tvar_20[3].label[84] );
tran (\_zy_simnet_tvar_20[3][92] , \_zy_simnet_tvar_20[3].label[83] );
tran (\_zy_simnet_tvar_20[3][91] , \_zy_simnet_tvar_20[3].label[82] );
tran (\_zy_simnet_tvar_20[3][90] , \_zy_simnet_tvar_20[3].label[81] );
tran (\_zy_simnet_tvar_20[3][89] , \_zy_simnet_tvar_20[3].label[80] );
tran (\_zy_simnet_tvar_20[3][88] , \_zy_simnet_tvar_20[3].label[79] );
tran (\_zy_simnet_tvar_20[3][87] , \_zy_simnet_tvar_20[3].label[78] );
tran (\_zy_simnet_tvar_20[3][86] , \_zy_simnet_tvar_20[3].label[77] );
tran (\_zy_simnet_tvar_20[3][85] , \_zy_simnet_tvar_20[3].label[76] );
tran (\_zy_simnet_tvar_20[3][84] , \_zy_simnet_tvar_20[3].label[75] );
tran (\_zy_simnet_tvar_20[3][83] , \_zy_simnet_tvar_20[3].label[74] );
tran (\_zy_simnet_tvar_20[3][82] , \_zy_simnet_tvar_20[3].label[73] );
tran (\_zy_simnet_tvar_20[3][81] , \_zy_simnet_tvar_20[3].label[72] );
tran (\_zy_simnet_tvar_20[3][80] , \_zy_simnet_tvar_20[3].label[71] );
tran (\_zy_simnet_tvar_20[3][79] , \_zy_simnet_tvar_20[3].label[70] );
tran (\_zy_simnet_tvar_20[3][78] , \_zy_simnet_tvar_20[3].label[69] );
tran (\_zy_simnet_tvar_20[3][77] , \_zy_simnet_tvar_20[3].label[68] );
tran (\_zy_simnet_tvar_20[3][76] , \_zy_simnet_tvar_20[3].label[67] );
tran (\_zy_simnet_tvar_20[3][75] , \_zy_simnet_tvar_20[3].label[66] );
tran (\_zy_simnet_tvar_20[3][74] , \_zy_simnet_tvar_20[3].label[65] );
tran (\_zy_simnet_tvar_20[3][73] , \_zy_simnet_tvar_20[3].label[64] );
tran (\_zy_simnet_tvar_20[3][72] , \_zy_simnet_tvar_20[3].label[63] );
tran (\_zy_simnet_tvar_20[3][71] , \_zy_simnet_tvar_20[3].label[62] );
tran (\_zy_simnet_tvar_20[3][70] , \_zy_simnet_tvar_20[3].label[61] );
tran (\_zy_simnet_tvar_20[3][69] , \_zy_simnet_tvar_20[3].label[60] );
tran (\_zy_simnet_tvar_20[3][68] , \_zy_simnet_tvar_20[3].label[59] );
tran (\_zy_simnet_tvar_20[3][67] , \_zy_simnet_tvar_20[3].label[58] );
tran (\_zy_simnet_tvar_20[3][66] , \_zy_simnet_tvar_20[3].label[57] );
tran (\_zy_simnet_tvar_20[3][65] , \_zy_simnet_tvar_20[3].label[56] );
tran (\_zy_simnet_tvar_20[3][64] , \_zy_simnet_tvar_20[3].label[55] );
tran (\_zy_simnet_tvar_20[3][63] , \_zy_simnet_tvar_20[3].label[54] );
tran (\_zy_simnet_tvar_20[3][62] , \_zy_simnet_tvar_20[3].label[53] );
tran (\_zy_simnet_tvar_20[3][61] , \_zy_simnet_tvar_20[3].label[52] );
tran (\_zy_simnet_tvar_20[3][60] , \_zy_simnet_tvar_20[3].label[51] );
tran (\_zy_simnet_tvar_20[3][59] , \_zy_simnet_tvar_20[3].label[50] );
tran (\_zy_simnet_tvar_20[3][58] , \_zy_simnet_tvar_20[3].label[49] );
tran (\_zy_simnet_tvar_20[3][57] , \_zy_simnet_tvar_20[3].label[48] );
tran (\_zy_simnet_tvar_20[3][56] , \_zy_simnet_tvar_20[3].label[47] );
tran (\_zy_simnet_tvar_20[3][55] , \_zy_simnet_tvar_20[3].label[46] );
tran (\_zy_simnet_tvar_20[3][54] , \_zy_simnet_tvar_20[3].label[45] );
tran (\_zy_simnet_tvar_20[3][53] , \_zy_simnet_tvar_20[3].label[44] );
tran (\_zy_simnet_tvar_20[3][52] , \_zy_simnet_tvar_20[3].label[43] );
tran (\_zy_simnet_tvar_20[3][51] , \_zy_simnet_tvar_20[3].label[42] );
tran (\_zy_simnet_tvar_20[3][50] , \_zy_simnet_tvar_20[3].label[41] );
tran (\_zy_simnet_tvar_20[3][49] , \_zy_simnet_tvar_20[3].label[40] );
tran (\_zy_simnet_tvar_20[3][48] , \_zy_simnet_tvar_20[3].label[39] );
tran (\_zy_simnet_tvar_20[3][47] , \_zy_simnet_tvar_20[3].label[38] );
tran (\_zy_simnet_tvar_20[3][46] , \_zy_simnet_tvar_20[3].label[37] );
tran (\_zy_simnet_tvar_20[3][45] , \_zy_simnet_tvar_20[3].label[36] );
tran (\_zy_simnet_tvar_20[3][44] , \_zy_simnet_tvar_20[3].label[35] );
tran (\_zy_simnet_tvar_20[3][43] , \_zy_simnet_tvar_20[3].label[34] );
tran (\_zy_simnet_tvar_20[3][42] , \_zy_simnet_tvar_20[3].label[33] );
tran (\_zy_simnet_tvar_20[3][41] , \_zy_simnet_tvar_20[3].label[32] );
tran (\_zy_simnet_tvar_20[3][40] , \_zy_simnet_tvar_20[3].label[31] );
tran (\_zy_simnet_tvar_20[3][39] , \_zy_simnet_tvar_20[3].label[30] );
tran (\_zy_simnet_tvar_20[3][38] , \_zy_simnet_tvar_20[3].label[29] );
tran (\_zy_simnet_tvar_20[3][37] , \_zy_simnet_tvar_20[3].label[28] );
tran (\_zy_simnet_tvar_20[3][36] , \_zy_simnet_tvar_20[3].label[27] );
tran (\_zy_simnet_tvar_20[3][35] , \_zy_simnet_tvar_20[3].label[26] );
tran (\_zy_simnet_tvar_20[3][34] , \_zy_simnet_tvar_20[3].label[25] );
tran (\_zy_simnet_tvar_20[3][33] , \_zy_simnet_tvar_20[3].label[24] );
tran (\_zy_simnet_tvar_20[3][32] , \_zy_simnet_tvar_20[3].label[23] );
tran (\_zy_simnet_tvar_20[3][31] , \_zy_simnet_tvar_20[3].label[22] );
tran (\_zy_simnet_tvar_20[3][30] , \_zy_simnet_tvar_20[3].label[21] );
tran (\_zy_simnet_tvar_20[3][29] , \_zy_simnet_tvar_20[3].label[20] );
tran (\_zy_simnet_tvar_20[3][28] , \_zy_simnet_tvar_20[3].label[19] );
tran (\_zy_simnet_tvar_20[3][27] , \_zy_simnet_tvar_20[3].label[18] );
tran (\_zy_simnet_tvar_20[3][26] , \_zy_simnet_tvar_20[3].label[17] );
tran (\_zy_simnet_tvar_20[3][25] , \_zy_simnet_tvar_20[3].label[16] );
tran (\_zy_simnet_tvar_20[3][24] , \_zy_simnet_tvar_20[3].label[15] );
tran (\_zy_simnet_tvar_20[3][23] , \_zy_simnet_tvar_20[3].label[14] );
tran (\_zy_simnet_tvar_20[3][22] , \_zy_simnet_tvar_20[3].label[13] );
tran (\_zy_simnet_tvar_20[3][21] , \_zy_simnet_tvar_20[3].label[12] );
tran (\_zy_simnet_tvar_20[3][20] , \_zy_simnet_tvar_20[3].label[11] );
tran (\_zy_simnet_tvar_20[3][19] , \_zy_simnet_tvar_20[3].label[10] );
tran (\_zy_simnet_tvar_20[3][18] , \_zy_simnet_tvar_20[3].label[9] );
tran (\_zy_simnet_tvar_20[3][17] , \_zy_simnet_tvar_20[3].label[8] );
tran (\_zy_simnet_tvar_20[3][16] , \_zy_simnet_tvar_20[3].label[7] );
tran (\_zy_simnet_tvar_20[3][15] , \_zy_simnet_tvar_20[3].label[6] );
tran (\_zy_simnet_tvar_20[3][14] , \_zy_simnet_tvar_20[3].label[5] );
tran (\_zy_simnet_tvar_20[3][13] , \_zy_simnet_tvar_20[3].label[4] );
tran (\_zy_simnet_tvar_20[3][12] , \_zy_simnet_tvar_20[3].label[3] );
tran (\_zy_simnet_tvar_20[3][11] , \_zy_simnet_tvar_20[3].label[2] );
tran (\_zy_simnet_tvar_20[3][10] , \_zy_simnet_tvar_20[3].label[1] );
tran (\_zy_simnet_tvar_20[3][9] , \_zy_simnet_tvar_20[3].label[0] );
tran (\_zy_simnet_tvar_20[3][8] , \_zy_simnet_tvar_20[3].delimiter_valid[0] );
tran (\_zy_simnet_tvar_20[3][7] , \_zy_simnet_tvar_20[3].delimiter[7] );
tran (\_zy_simnet_tvar_20[3][6] , \_zy_simnet_tvar_20[3].delimiter[6] );
tran (\_zy_simnet_tvar_20[3][5] , \_zy_simnet_tvar_20[3].delimiter[5] );
tran (\_zy_simnet_tvar_20[3][4] , \_zy_simnet_tvar_20[3].delimiter[4] );
tran (\_zy_simnet_tvar_20[3][3] , \_zy_simnet_tvar_20[3].delimiter[3] );
tran (\_zy_simnet_tvar_20[3][2] , \_zy_simnet_tvar_20[3].delimiter[2] );
tran (\_zy_simnet_tvar_20[3][1] , \_zy_simnet_tvar_20[3].delimiter[1] );
tran (\_zy_simnet_tvar_20[3][0] , \_zy_simnet_tvar_20[3].delimiter[0] );
tran (\_zy_simnet_tvar_20[2][271] , \_zy_simnet_tvar_20[2].guid_size[0] );
tran (\_zy_simnet_tvar_20[2][270] , \_zy_simnet_tvar_20[2].label_size[5] );
tran (\_zy_simnet_tvar_20[2][269] , \_zy_simnet_tvar_20[2].label_size[4] );
tran (\_zy_simnet_tvar_20[2][268] , \_zy_simnet_tvar_20[2].label_size[3] );
tran (\_zy_simnet_tvar_20[2][267] , \_zy_simnet_tvar_20[2].label_size[2] );
tran (\_zy_simnet_tvar_20[2][266] , \_zy_simnet_tvar_20[2].label_size[1] );
tran (\_zy_simnet_tvar_20[2][265] , \_zy_simnet_tvar_20[2].label_size[0] );
tran (\_zy_simnet_tvar_20[2][264] , \_zy_simnet_tvar_20[2].label[255] );
tran (\_zy_simnet_tvar_20[2][263] , \_zy_simnet_tvar_20[2].label[254] );
tran (\_zy_simnet_tvar_20[2][262] , \_zy_simnet_tvar_20[2].label[253] );
tran (\_zy_simnet_tvar_20[2][261] , \_zy_simnet_tvar_20[2].label[252] );
tran (\_zy_simnet_tvar_20[2][260] , \_zy_simnet_tvar_20[2].label[251] );
tran (\_zy_simnet_tvar_20[2][259] , \_zy_simnet_tvar_20[2].label[250] );
tran (\_zy_simnet_tvar_20[2][258] , \_zy_simnet_tvar_20[2].label[249] );
tran (\_zy_simnet_tvar_20[2][257] , \_zy_simnet_tvar_20[2].label[248] );
tran (\_zy_simnet_tvar_20[2][256] , \_zy_simnet_tvar_20[2].label[247] );
tran (\_zy_simnet_tvar_20[2][255] , \_zy_simnet_tvar_20[2].label[246] );
tran (\_zy_simnet_tvar_20[2][254] , \_zy_simnet_tvar_20[2].label[245] );
tran (\_zy_simnet_tvar_20[2][253] , \_zy_simnet_tvar_20[2].label[244] );
tran (\_zy_simnet_tvar_20[2][252] , \_zy_simnet_tvar_20[2].label[243] );
tran (\_zy_simnet_tvar_20[2][251] , \_zy_simnet_tvar_20[2].label[242] );
tran (\_zy_simnet_tvar_20[2][250] , \_zy_simnet_tvar_20[2].label[241] );
tran (\_zy_simnet_tvar_20[2][249] , \_zy_simnet_tvar_20[2].label[240] );
tran (\_zy_simnet_tvar_20[2][248] , \_zy_simnet_tvar_20[2].label[239] );
tran (\_zy_simnet_tvar_20[2][247] , \_zy_simnet_tvar_20[2].label[238] );
tran (\_zy_simnet_tvar_20[2][246] , \_zy_simnet_tvar_20[2].label[237] );
tran (\_zy_simnet_tvar_20[2][245] , \_zy_simnet_tvar_20[2].label[236] );
tran (\_zy_simnet_tvar_20[2][244] , \_zy_simnet_tvar_20[2].label[235] );
tran (\_zy_simnet_tvar_20[2][243] , \_zy_simnet_tvar_20[2].label[234] );
tran (\_zy_simnet_tvar_20[2][242] , \_zy_simnet_tvar_20[2].label[233] );
tran (\_zy_simnet_tvar_20[2][241] , \_zy_simnet_tvar_20[2].label[232] );
tran (\_zy_simnet_tvar_20[2][240] , \_zy_simnet_tvar_20[2].label[231] );
tran (\_zy_simnet_tvar_20[2][239] , \_zy_simnet_tvar_20[2].label[230] );
tran (\_zy_simnet_tvar_20[2][238] , \_zy_simnet_tvar_20[2].label[229] );
tran (\_zy_simnet_tvar_20[2][237] , \_zy_simnet_tvar_20[2].label[228] );
tran (\_zy_simnet_tvar_20[2][236] , \_zy_simnet_tvar_20[2].label[227] );
tran (\_zy_simnet_tvar_20[2][235] , \_zy_simnet_tvar_20[2].label[226] );
tran (\_zy_simnet_tvar_20[2][234] , \_zy_simnet_tvar_20[2].label[225] );
tran (\_zy_simnet_tvar_20[2][233] , \_zy_simnet_tvar_20[2].label[224] );
tran (\_zy_simnet_tvar_20[2][232] , \_zy_simnet_tvar_20[2].label[223] );
tran (\_zy_simnet_tvar_20[2][231] , \_zy_simnet_tvar_20[2].label[222] );
tran (\_zy_simnet_tvar_20[2][230] , \_zy_simnet_tvar_20[2].label[221] );
tran (\_zy_simnet_tvar_20[2][229] , \_zy_simnet_tvar_20[2].label[220] );
tran (\_zy_simnet_tvar_20[2][228] , \_zy_simnet_tvar_20[2].label[219] );
tran (\_zy_simnet_tvar_20[2][227] , \_zy_simnet_tvar_20[2].label[218] );
tran (\_zy_simnet_tvar_20[2][226] , \_zy_simnet_tvar_20[2].label[217] );
tran (\_zy_simnet_tvar_20[2][225] , \_zy_simnet_tvar_20[2].label[216] );
tran (\_zy_simnet_tvar_20[2][224] , \_zy_simnet_tvar_20[2].label[215] );
tran (\_zy_simnet_tvar_20[2][223] , \_zy_simnet_tvar_20[2].label[214] );
tran (\_zy_simnet_tvar_20[2][222] , \_zy_simnet_tvar_20[2].label[213] );
tran (\_zy_simnet_tvar_20[2][221] , \_zy_simnet_tvar_20[2].label[212] );
tran (\_zy_simnet_tvar_20[2][220] , \_zy_simnet_tvar_20[2].label[211] );
tran (\_zy_simnet_tvar_20[2][219] , \_zy_simnet_tvar_20[2].label[210] );
tran (\_zy_simnet_tvar_20[2][218] , \_zy_simnet_tvar_20[2].label[209] );
tran (\_zy_simnet_tvar_20[2][217] , \_zy_simnet_tvar_20[2].label[208] );
tran (\_zy_simnet_tvar_20[2][216] , \_zy_simnet_tvar_20[2].label[207] );
tran (\_zy_simnet_tvar_20[2][215] , \_zy_simnet_tvar_20[2].label[206] );
tran (\_zy_simnet_tvar_20[2][214] , \_zy_simnet_tvar_20[2].label[205] );
tran (\_zy_simnet_tvar_20[2][213] , \_zy_simnet_tvar_20[2].label[204] );
tran (\_zy_simnet_tvar_20[2][212] , \_zy_simnet_tvar_20[2].label[203] );
tran (\_zy_simnet_tvar_20[2][211] , \_zy_simnet_tvar_20[2].label[202] );
tran (\_zy_simnet_tvar_20[2][210] , \_zy_simnet_tvar_20[2].label[201] );
tran (\_zy_simnet_tvar_20[2][209] , \_zy_simnet_tvar_20[2].label[200] );
tran (\_zy_simnet_tvar_20[2][208] , \_zy_simnet_tvar_20[2].label[199] );
tran (\_zy_simnet_tvar_20[2][207] , \_zy_simnet_tvar_20[2].label[198] );
tran (\_zy_simnet_tvar_20[2][206] , \_zy_simnet_tvar_20[2].label[197] );
tran (\_zy_simnet_tvar_20[2][205] , \_zy_simnet_tvar_20[2].label[196] );
tran (\_zy_simnet_tvar_20[2][204] , \_zy_simnet_tvar_20[2].label[195] );
tran (\_zy_simnet_tvar_20[2][203] , \_zy_simnet_tvar_20[2].label[194] );
tran (\_zy_simnet_tvar_20[2][202] , \_zy_simnet_tvar_20[2].label[193] );
tran (\_zy_simnet_tvar_20[2][201] , \_zy_simnet_tvar_20[2].label[192] );
tran (\_zy_simnet_tvar_20[2][200] , \_zy_simnet_tvar_20[2].label[191] );
tran (\_zy_simnet_tvar_20[2][199] , \_zy_simnet_tvar_20[2].label[190] );
tran (\_zy_simnet_tvar_20[2][198] , \_zy_simnet_tvar_20[2].label[189] );
tran (\_zy_simnet_tvar_20[2][197] , \_zy_simnet_tvar_20[2].label[188] );
tran (\_zy_simnet_tvar_20[2][196] , \_zy_simnet_tvar_20[2].label[187] );
tran (\_zy_simnet_tvar_20[2][195] , \_zy_simnet_tvar_20[2].label[186] );
tran (\_zy_simnet_tvar_20[2][194] , \_zy_simnet_tvar_20[2].label[185] );
tran (\_zy_simnet_tvar_20[2][193] , \_zy_simnet_tvar_20[2].label[184] );
tran (\_zy_simnet_tvar_20[2][192] , \_zy_simnet_tvar_20[2].label[183] );
tran (\_zy_simnet_tvar_20[2][191] , \_zy_simnet_tvar_20[2].label[182] );
tran (\_zy_simnet_tvar_20[2][190] , \_zy_simnet_tvar_20[2].label[181] );
tran (\_zy_simnet_tvar_20[2][189] , \_zy_simnet_tvar_20[2].label[180] );
tran (\_zy_simnet_tvar_20[2][188] , \_zy_simnet_tvar_20[2].label[179] );
tran (\_zy_simnet_tvar_20[2][187] , \_zy_simnet_tvar_20[2].label[178] );
tran (\_zy_simnet_tvar_20[2][186] , \_zy_simnet_tvar_20[2].label[177] );
tran (\_zy_simnet_tvar_20[2][185] , \_zy_simnet_tvar_20[2].label[176] );
tran (\_zy_simnet_tvar_20[2][184] , \_zy_simnet_tvar_20[2].label[175] );
tran (\_zy_simnet_tvar_20[2][183] , \_zy_simnet_tvar_20[2].label[174] );
tran (\_zy_simnet_tvar_20[2][182] , \_zy_simnet_tvar_20[2].label[173] );
tran (\_zy_simnet_tvar_20[2][181] , \_zy_simnet_tvar_20[2].label[172] );
tran (\_zy_simnet_tvar_20[2][180] , \_zy_simnet_tvar_20[2].label[171] );
tran (\_zy_simnet_tvar_20[2][179] , \_zy_simnet_tvar_20[2].label[170] );
tran (\_zy_simnet_tvar_20[2][178] , \_zy_simnet_tvar_20[2].label[169] );
tran (\_zy_simnet_tvar_20[2][177] , \_zy_simnet_tvar_20[2].label[168] );
tran (\_zy_simnet_tvar_20[2][176] , \_zy_simnet_tvar_20[2].label[167] );
tran (\_zy_simnet_tvar_20[2][175] , \_zy_simnet_tvar_20[2].label[166] );
tran (\_zy_simnet_tvar_20[2][174] , \_zy_simnet_tvar_20[2].label[165] );
tran (\_zy_simnet_tvar_20[2][173] , \_zy_simnet_tvar_20[2].label[164] );
tran (\_zy_simnet_tvar_20[2][172] , \_zy_simnet_tvar_20[2].label[163] );
tran (\_zy_simnet_tvar_20[2][171] , \_zy_simnet_tvar_20[2].label[162] );
tran (\_zy_simnet_tvar_20[2][170] , \_zy_simnet_tvar_20[2].label[161] );
tran (\_zy_simnet_tvar_20[2][169] , \_zy_simnet_tvar_20[2].label[160] );
tran (\_zy_simnet_tvar_20[2][168] , \_zy_simnet_tvar_20[2].label[159] );
tran (\_zy_simnet_tvar_20[2][167] , \_zy_simnet_tvar_20[2].label[158] );
tran (\_zy_simnet_tvar_20[2][166] , \_zy_simnet_tvar_20[2].label[157] );
tran (\_zy_simnet_tvar_20[2][165] , \_zy_simnet_tvar_20[2].label[156] );
tran (\_zy_simnet_tvar_20[2][164] , \_zy_simnet_tvar_20[2].label[155] );
tran (\_zy_simnet_tvar_20[2][163] , \_zy_simnet_tvar_20[2].label[154] );
tran (\_zy_simnet_tvar_20[2][162] , \_zy_simnet_tvar_20[2].label[153] );
tran (\_zy_simnet_tvar_20[2][161] , \_zy_simnet_tvar_20[2].label[152] );
tran (\_zy_simnet_tvar_20[2][160] , \_zy_simnet_tvar_20[2].label[151] );
tran (\_zy_simnet_tvar_20[2][159] , \_zy_simnet_tvar_20[2].label[150] );
tran (\_zy_simnet_tvar_20[2][158] , \_zy_simnet_tvar_20[2].label[149] );
tran (\_zy_simnet_tvar_20[2][157] , \_zy_simnet_tvar_20[2].label[148] );
tran (\_zy_simnet_tvar_20[2][156] , \_zy_simnet_tvar_20[2].label[147] );
tran (\_zy_simnet_tvar_20[2][155] , \_zy_simnet_tvar_20[2].label[146] );
tran (\_zy_simnet_tvar_20[2][154] , \_zy_simnet_tvar_20[2].label[145] );
tran (\_zy_simnet_tvar_20[2][153] , \_zy_simnet_tvar_20[2].label[144] );
tran (\_zy_simnet_tvar_20[2][152] , \_zy_simnet_tvar_20[2].label[143] );
tran (\_zy_simnet_tvar_20[2][151] , \_zy_simnet_tvar_20[2].label[142] );
tran (\_zy_simnet_tvar_20[2][150] , \_zy_simnet_tvar_20[2].label[141] );
tran (\_zy_simnet_tvar_20[2][149] , \_zy_simnet_tvar_20[2].label[140] );
tran (\_zy_simnet_tvar_20[2][148] , \_zy_simnet_tvar_20[2].label[139] );
tran (\_zy_simnet_tvar_20[2][147] , \_zy_simnet_tvar_20[2].label[138] );
tran (\_zy_simnet_tvar_20[2][146] , \_zy_simnet_tvar_20[2].label[137] );
tran (\_zy_simnet_tvar_20[2][145] , \_zy_simnet_tvar_20[2].label[136] );
tran (\_zy_simnet_tvar_20[2][144] , \_zy_simnet_tvar_20[2].label[135] );
tran (\_zy_simnet_tvar_20[2][143] , \_zy_simnet_tvar_20[2].label[134] );
tran (\_zy_simnet_tvar_20[2][142] , \_zy_simnet_tvar_20[2].label[133] );
tran (\_zy_simnet_tvar_20[2][141] , \_zy_simnet_tvar_20[2].label[132] );
tran (\_zy_simnet_tvar_20[2][140] , \_zy_simnet_tvar_20[2].label[131] );
tran (\_zy_simnet_tvar_20[2][139] , \_zy_simnet_tvar_20[2].label[130] );
tran (\_zy_simnet_tvar_20[2][138] , \_zy_simnet_tvar_20[2].label[129] );
tran (\_zy_simnet_tvar_20[2][137] , \_zy_simnet_tvar_20[2].label[128] );
tran (\_zy_simnet_tvar_20[2][136] , \_zy_simnet_tvar_20[2].label[127] );
tran (\_zy_simnet_tvar_20[2][135] , \_zy_simnet_tvar_20[2].label[126] );
tran (\_zy_simnet_tvar_20[2][134] , \_zy_simnet_tvar_20[2].label[125] );
tran (\_zy_simnet_tvar_20[2][133] , \_zy_simnet_tvar_20[2].label[124] );
tran (\_zy_simnet_tvar_20[2][132] , \_zy_simnet_tvar_20[2].label[123] );
tran (\_zy_simnet_tvar_20[2][131] , \_zy_simnet_tvar_20[2].label[122] );
tran (\_zy_simnet_tvar_20[2][130] , \_zy_simnet_tvar_20[2].label[121] );
tran (\_zy_simnet_tvar_20[2][129] , \_zy_simnet_tvar_20[2].label[120] );
tran (\_zy_simnet_tvar_20[2][128] , \_zy_simnet_tvar_20[2].label[119] );
tran (\_zy_simnet_tvar_20[2][127] , \_zy_simnet_tvar_20[2].label[118] );
tran (\_zy_simnet_tvar_20[2][126] , \_zy_simnet_tvar_20[2].label[117] );
tran (\_zy_simnet_tvar_20[2][125] , \_zy_simnet_tvar_20[2].label[116] );
tran (\_zy_simnet_tvar_20[2][124] , \_zy_simnet_tvar_20[2].label[115] );
tran (\_zy_simnet_tvar_20[2][123] , \_zy_simnet_tvar_20[2].label[114] );
tran (\_zy_simnet_tvar_20[2][122] , \_zy_simnet_tvar_20[2].label[113] );
tran (\_zy_simnet_tvar_20[2][121] , \_zy_simnet_tvar_20[2].label[112] );
tran (\_zy_simnet_tvar_20[2][120] , \_zy_simnet_tvar_20[2].label[111] );
tran (\_zy_simnet_tvar_20[2][119] , \_zy_simnet_tvar_20[2].label[110] );
tran (\_zy_simnet_tvar_20[2][118] , \_zy_simnet_tvar_20[2].label[109] );
tran (\_zy_simnet_tvar_20[2][117] , \_zy_simnet_tvar_20[2].label[108] );
tran (\_zy_simnet_tvar_20[2][116] , \_zy_simnet_tvar_20[2].label[107] );
tran (\_zy_simnet_tvar_20[2][115] , \_zy_simnet_tvar_20[2].label[106] );
tran (\_zy_simnet_tvar_20[2][114] , \_zy_simnet_tvar_20[2].label[105] );
tran (\_zy_simnet_tvar_20[2][113] , \_zy_simnet_tvar_20[2].label[104] );
tran (\_zy_simnet_tvar_20[2][112] , \_zy_simnet_tvar_20[2].label[103] );
tran (\_zy_simnet_tvar_20[2][111] , \_zy_simnet_tvar_20[2].label[102] );
tran (\_zy_simnet_tvar_20[2][110] , \_zy_simnet_tvar_20[2].label[101] );
tran (\_zy_simnet_tvar_20[2][109] , \_zy_simnet_tvar_20[2].label[100] );
tran (\_zy_simnet_tvar_20[2][108] , \_zy_simnet_tvar_20[2].label[99] );
tran (\_zy_simnet_tvar_20[2][107] , \_zy_simnet_tvar_20[2].label[98] );
tran (\_zy_simnet_tvar_20[2][106] , \_zy_simnet_tvar_20[2].label[97] );
tran (\_zy_simnet_tvar_20[2][105] , \_zy_simnet_tvar_20[2].label[96] );
tran (\_zy_simnet_tvar_20[2][104] , \_zy_simnet_tvar_20[2].label[95] );
tran (\_zy_simnet_tvar_20[2][103] , \_zy_simnet_tvar_20[2].label[94] );
tran (\_zy_simnet_tvar_20[2][102] , \_zy_simnet_tvar_20[2].label[93] );
tran (\_zy_simnet_tvar_20[2][101] , \_zy_simnet_tvar_20[2].label[92] );
tran (\_zy_simnet_tvar_20[2][100] , \_zy_simnet_tvar_20[2].label[91] );
tran (\_zy_simnet_tvar_20[2][99] , \_zy_simnet_tvar_20[2].label[90] );
tran (\_zy_simnet_tvar_20[2][98] , \_zy_simnet_tvar_20[2].label[89] );
tran (\_zy_simnet_tvar_20[2][97] , \_zy_simnet_tvar_20[2].label[88] );
tran (\_zy_simnet_tvar_20[2][96] , \_zy_simnet_tvar_20[2].label[87] );
tran (\_zy_simnet_tvar_20[2][95] , \_zy_simnet_tvar_20[2].label[86] );
tran (\_zy_simnet_tvar_20[2][94] , \_zy_simnet_tvar_20[2].label[85] );
tran (\_zy_simnet_tvar_20[2][93] , \_zy_simnet_tvar_20[2].label[84] );
tran (\_zy_simnet_tvar_20[2][92] , \_zy_simnet_tvar_20[2].label[83] );
tran (\_zy_simnet_tvar_20[2][91] , \_zy_simnet_tvar_20[2].label[82] );
tran (\_zy_simnet_tvar_20[2][90] , \_zy_simnet_tvar_20[2].label[81] );
tran (\_zy_simnet_tvar_20[2][89] , \_zy_simnet_tvar_20[2].label[80] );
tran (\_zy_simnet_tvar_20[2][88] , \_zy_simnet_tvar_20[2].label[79] );
tran (\_zy_simnet_tvar_20[2][87] , \_zy_simnet_tvar_20[2].label[78] );
tran (\_zy_simnet_tvar_20[2][86] , \_zy_simnet_tvar_20[2].label[77] );
tran (\_zy_simnet_tvar_20[2][85] , \_zy_simnet_tvar_20[2].label[76] );
tran (\_zy_simnet_tvar_20[2][84] , \_zy_simnet_tvar_20[2].label[75] );
tran (\_zy_simnet_tvar_20[2][83] , \_zy_simnet_tvar_20[2].label[74] );
tran (\_zy_simnet_tvar_20[2][82] , \_zy_simnet_tvar_20[2].label[73] );
tran (\_zy_simnet_tvar_20[2][81] , \_zy_simnet_tvar_20[2].label[72] );
tran (\_zy_simnet_tvar_20[2][80] , \_zy_simnet_tvar_20[2].label[71] );
tran (\_zy_simnet_tvar_20[2][79] , \_zy_simnet_tvar_20[2].label[70] );
tran (\_zy_simnet_tvar_20[2][78] , \_zy_simnet_tvar_20[2].label[69] );
tran (\_zy_simnet_tvar_20[2][77] , \_zy_simnet_tvar_20[2].label[68] );
tran (\_zy_simnet_tvar_20[2][76] , \_zy_simnet_tvar_20[2].label[67] );
tran (\_zy_simnet_tvar_20[2][75] , \_zy_simnet_tvar_20[2].label[66] );
tran (\_zy_simnet_tvar_20[2][74] , \_zy_simnet_tvar_20[2].label[65] );
tran (\_zy_simnet_tvar_20[2][73] , \_zy_simnet_tvar_20[2].label[64] );
tran (\_zy_simnet_tvar_20[2][72] , \_zy_simnet_tvar_20[2].label[63] );
tran (\_zy_simnet_tvar_20[2][71] , \_zy_simnet_tvar_20[2].label[62] );
tran (\_zy_simnet_tvar_20[2][70] , \_zy_simnet_tvar_20[2].label[61] );
tran (\_zy_simnet_tvar_20[2][69] , \_zy_simnet_tvar_20[2].label[60] );
tran (\_zy_simnet_tvar_20[2][68] , \_zy_simnet_tvar_20[2].label[59] );
tran (\_zy_simnet_tvar_20[2][67] , \_zy_simnet_tvar_20[2].label[58] );
tran (\_zy_simnet_tvar_20[2][66] , \_zy_simnet_tvar_20[2].label[57] );
tran (\_zy_simnet_tvar_20[2][65] , \_zy_simnet_tvar_20[2].label[56] );
tran (\_zy_simnet_tvar_20[2][64] , \_zy_simnet_tvar_20[2].label[55] );
tran (\_zy_simnet_tvar_20[2][63] , \_zy_simnet_tvar_20[2].label[54] );
tran (\_zy_simnet_tvar_20[2][62] , \_zy_simnet_tvar_20[2].label[53] );
tran (\_zy_simnet_tvar_20[2][61] , \_zy_simnet_tvar_20[2].label[52] );
tran (\_zy_simnet_tvar_20[2][60] , \_zy_simnet_tvar_20[2].label[51] );
tran (\_zy_simnet_tvar_20[2][59] , \_zy_simnet_tvar_20[2].label[50] );
tran (\_zy_simnet_tvar_20[2][58] , \_zy_simnet_tvar_20[2].label[49] );
tran (\_zy_simnet_tvar_20[2][57] , \_zy_simnet_tvar_20[2].label[48] );
tran (\_zy_simnet_tvar_20[2][56] , \_zy_simnet_tvar_20[2].label[47] );
tran (\_zy_simnet_tvar_20[2][55] , \_zy_simnet_tvar_20[2].label[46] );
tran (\_zy_simnet_tvar_20[2][54] , \_zy_simnet_tvar_20[2].label[45] );
tran (\_zy_simnet_tvar_20[2][53] , \_zy_simnet_tvar_20[2].label[44] );
tran (\_zy_simnet_tvar_20[2][52] , \_zy_simnet_tvar_20[2].label[43] );
tran (\_zy_simnet_tvar_20[2][51] , \_zy_simnet_tvar_20[2].label[42] );
tran (\_zy_simnet_tvar_20[2][50] , \_zy_simnet_tvar_20[2].label[41] );
tran (\_zy_simnet_tvar_20[2][49] , \_zy_simnet_tvar_20[2].label[40] );
tran (\_zy_simnet_tvar_20[2][48] , \_zy_simnet_tvar_20[2].label[39] );
tran (\_zy_simnet_tvar_20[2][47] , \_zy_simnet_tvar_20[2].label[38] );
tran (\_zy_simnet_tvar_20[2][46] , \_zy_simnet_tvar_20[2].label[37] );
tran (\_zy_simnet_tvar_20[2][45] , \_zy_simnet_tvar_20[2].label[36] );
tran (\_zy_simnet_tvar_20[2][44] , \_zy_simnet_tvar_20[2].label[35] );
tran (\_zy_simnet_tvar_20[2][43] , \_zy_simnet_tvar_20[2].label[34] );
tran (\_zy_simnet_tvar_20[2][42] , \_zy_simnet_tvar_20[2].label[33] );
tran (\_zy_simnet_tvar_20[2][41] , \_zy_simnet_tvar_20[2].label[32] );
tran (\_zy_simnet_tvar_20[2][40] , \_zy_simnet_tvar_20[2].label[31] );
tran (\_zy_simnet_tvar_20[2][39] , \_zy_simnet_tvar_20[2].label[30] );
tran (\_zy_simnet_tvar_20[2][38] , \_zy_simnet_tvar_20[2].label[29] );
tran (\_zy_simnet_tvar_20[2][37] , \_zy_simnet_tvar_20[2].label[28] );
tran (\_zy_simnet_tvar_20[2][36] , \_zy_simnet_tvar_20[2].label[27] );
tran (\_zy_simnet_tvar_20[2][35] , \_zy_simnet_tvar_20[2].label[26] );
tran (\_zy_simnet_tvar_20[2][34] , \_zy_simnet_tvar_20[2].label[25] );
tran (\_zy_simnet_tvar_20[2][33] , \_zy_simnet_tvar_20[2].label[24] );
tran (\_zy_simnet_tvar_20[2][32] , \_zy_simnet_tvar_20[2].label[23] );
tran (\_zy_simnet_tvar_20[2][31] , \_zy_simnet_tvar_20[2].label[22] );
tran (\_zy_simnet_tvar_20[2][30] , \_zy_simnet_tvar_20[2].label[21] );
tran (\_zy_simnet_tvar_20[2][29] , \_zy_simnet_tvar_20[2].label[20] );
tran (\_zy_simnet_tvar_20[2][28] , \_zy_simnet_tvar_20[2].label[19] );
tran (\_zy_simnet_tvar_20[2][27] , \_zy_simnet_tvar_20[2].label[18] );
tran (\_zy_simnet_tvar_20[2][26] , \_zy_simnet_tvar_20[2].label[17] );
tran (\_zy_simnet_tvar_20[2][25] , \_zy_simnet_tvar_20[2].label[16] );
tran (\_zy_simnet_tvar_20[2][24] , \_zy_simnet_tvar_20[2].label[15] );
tran (\_zy_simnet_tvar_20[2][23] , \_zy_simnet_tvar_20[2].label[14] );
tran (\_zy_simnet_tvar_20[2][22] , \_zy_simnet_tvar_20[2].label[13] );
tran (\_zy_simnet_tvar_20[2][21] , \_zy_simnet_tvar_20[2].label[12] );
tran (\_zy_simnet_tvar_20[2][20] , \_zy_simnet_tvar_20[2].label[11] );
tran (\_zy_simnet_tvar_20[2][19] , \_zy_simnet_tvar_20[2].label[10] );
tran (\_zy_simnet_tvar_20[2][18] , \_zy_simnet_tvar_20[2].label[9] );
tran (\_zy_simnet_tvar_20[2][17] , \_zy_simnet_tvar_20[2].label[8] );
tran (\_zy_simnet_tvar_20[2][16] , \_zy_simnet_tvar_20[2].label[7] );
tran (\_zy_simnet_tvar_20[2][15] , \_zy_simnet_tvar_20[2].label[6] );
tran (\_zy_simnet_tvar_20[2][14] , \_zy_simnet_tvar_20[2].label[5] );
tran (\_zy_simnet_tvar_20[2][13] , \_zy_simnet_tvar_20[2].label[4] );
tran (\_zy_simnet_tvar_20[2][12] , \_zy_simnet_tvar_20[2].label[3] );
tran (\_zy_simnet_tvar_20[2][11] , \_zy_simnet_tvar_20[2].label[2] );
tran (\_zy_simnet_tvar_20[2][10] , \_zy_simnet_tvar_20[2].label[1] );
tran (\_zy_simnet_tvar_20[2][9] , \_zy_simnet_tvar_20[2].label[0] );
tran (\_zy_simnet_tvar_20[2][8] , \_zy_simnet_tvar_20[2].delimiter_valid[0] );
tran (\_zy_simnet_tvar_20[2][7] , \_zy_simnet_tvar_20[2].delimiter[7] );
tran (\_zy_simnet_tvar_20[2][6] , \_zy_simnet_tvar_20[2].delimiter[6] );
tran (\_zy_simnet_tvar_20[2][5] , \_zy_simnet_tvar_20[2].delimiter[5] );
tran (\_zy_simnet_tvar_20[2][4] , \_zy_simnet_tvar_20[2].delimiter[4] );
tran (\_zy_simnet_tvar_20[2][3] , \_zy_simnet_tvar_20[2].delimiter[3] );
tran (\_zy_simnet_tvar_20[2][2] , \_zy_simnet_tvar_20[2].delimiter[2] );
tran (\_zy_simnet_tvar_20[2][1] , \_zy_simnet_tvar_20[2].delimiter[1] );
tran (\_zy_simnet_tvar_20[2][0] , \_zy_simnet_tvar_20[2].delimiter[0] );
tran (\_zy_simnet_tvar_20[1][271] , \_zy_simnet_tvar_20[1].guid_size[0] );
tran (\_zy_simnet_tvar_20[1][270] , \_zy_simnet_tvar_20[1].label_size[5] );
tran (\_zy_simnet_tvar_20[1][269] , \_zy_simnet_tvar_20[1].label_size[4] );
tran (\_zy_simnet_tvar_20[1][268] , \_zy_simnet_tvar_20[1].label_size[3] );
tran (\_zy_simnet_tvar_20[1][267] , \_zy_simnet_tvar_20[1].label_size[2] );
tran (\_zy_simnet_tvar_20[1][266] , \_zy_simnet_tvar_20[1].label_size[1] );
tran (\_zy_simnet_tvar_20[1][265] , \_zy_simnet_tvar_20[1].label_size[0] );
tran (\_zy_simnet_tvar_20[1][264] , \_zy_simnet_tvar_20[1].label[255] );
tran (\_zy_simnet_tvar_20[1][263] , \_zy_simnet_tvar_20[1].label[254] );
tran (\_zy_simnet_tvar_20[1][262] , \_zy_simnet_tvar_20[1].label[253] );
tran (\_zy_simnet_tvar_20[1][261] , \_zy_simnet_tvar_20[1].label[252] );
tran (\_zy_simnet_tvar_20[1][260] , \_zy_simnet_tvar_20[1].label[251] );
tran (\_zy_simnet_tvar_20[1][259] , \_zy_simnet_tvar_20[1].label[250] );
tran (\_zy_simnet_tvar_20[1][258] , \_zy_simnet_tvar_20[1].label[249] );
tran (\_zy_simnet_tvar_20[1][257] , \_zy_simnet_tvar_20[1].label[248] );
tran (\_zy_simnet_tvar_20[1][256] , \_zy_simnet_tvar_20[1].label[247] );
tran (\_zy_simnet_tvar_20[1][255] , \_zy_simnet_tvar_20[1].label[246] );
tran (\_zy_simnet_tvar_20[1][254] , \_zy_simnet_tvar_20[1].label[245] );
tran (\_zy_simnet_tvar_20[1][253] , \_zy_simnet_tvar_20[1].label[244] );
tran (\_zy_simnet_tvar_20[1][252] , \_zy_simnet_tvar_20[1].label[243] );
tran (\_zy_simnet_tvar_20[1][251] , \_zy_simnet_tvar_20[1].label[242] );
tran (\_zy_simnet_tvar_20[1][250] , \_zy_simnet_tvar_20[1].label[241] );
tran (\_zy_simnet_tvar_20[1][249] , \_zy_simnet_tvar_20[1].label[240] );
tran (\_zy_simnet_tvar_20[1][248] , \_zy_simnet_tvar_20[1].label[239] );
tran (\_zy_simnet_tvar_20[1][247] , \_zy_simnet_tvar_20[1].label[238] );
tran (\_zy_simnet_tvar_20[1][246] , \_zy_simnet_tvar_20[1].label[237] );
tran (\_zy_simnet_tvar_20[1][245] , \_zy_simnet_tvar_20[1].label[236] );
tran (\_zy_simnet_tvar_20[1][244] , \_zy_simnet_tvar_20[1].label[235] );
tran (\_zy_simnet_tvar_20[1][243] , \_zy_simnet_tvar_20[1].label[234] );
tran (\_zy_simnet_tvar_20[1][242] , \_zy_simnet_tvar_20[1].label[233] );
tran (\_zy_simnet_tvar_20[1][241] , \_zy_simnet_tvar_20[1].label[232] );
tran (\_zy_simnet_tvar_20[1][240] , \_zy_simnet_tvar_20[1].label[231] );
tran (\_zy_simnet_tvar_20[1][239] , \_zy_simnet_tvar_20[1].label[230] );
tran (\_zy_simnet_tvar_20[1][238] , \_zy_simnet_tvar_20[1].label[229] );
tran (\_zy_simnet_tvar_20[1][237] , \_zy_simnet_tvar_20[1].label[228] );
tran (\_zy_simnet_tvar_20[1][236] , \_zy_simnet_tvar_20[1].label[227] );
tran (\_zy_simnet_tvar_20[1][235] , \_zy_simnet_tvar_20[1].label[226] );
tran (\_zy_simnet_tvar_20[1][234] , \_zy_simnet_tvar_20[1].label[225] );
tran (\_zy_simnet_tvar_20[1][233] , \_zy_simnet_tvar_20[1].label[224] );
tran (\_zy_simnet_tvar_20[1][232] , \_zy_simnet_tvar_20[1].label[223] );
tran (\_zy_simnet_tvar_20[1][231] , \_zy_simnet_tvar_20[1].label[222] );
tran (\_zy_simnet_tvar_20[1][230] , \_zy_simnet_tvar_20[1].label[221] );
tran (\_zy_simnet_tvar_20[1][229] , \_zy_simnet_tvar_20[1].label[220] );
tran (\_zy_simnet_tvar_20[1][228] , \_zy_simnet_tvar_20[1].label[219] );
tran (\_zy_simnet_tvar_20[1][227] , \_zy_simnet_tvar_20[1].label[218] );
tran (\_zy_simnet_tvar_20[1][226] , \_zy_simnet_tvar_20[1].label[217] );
tran (\_zy_simnet_tvar_20[1][225] , \_zy_simnet_tvar_20[1].label[216] );
tran (\_zy_simnet_tvar_20[1][224] , \_zy_simnet_tvar_20[1].label[215] );
tran (\_zy_simnet_tvar_20[1][223] , \_zy_simnet_tvar_20[1].label[214] );
tran (\_zy_simnet_tvar_20[1][222] , \_zy_simnet_tvar_20[1].label[213] );
tran (\_zy_simnet_tvar_20[1][221] , \_zy_simnet_tvar_20[1].label[212] );
tran (\_zy_simnet_tvar_20[1][220] , \_zy_simnet_tvar_20[1].label[211] );
tran (\_zy_simnet_tvar_20[1][219] , \_zy_simnet_tvar_20[1].label[210] );
tran (\_zy_simnet_tvar_20[1][218] , \_zy_simnet_tvar_20[1].label[209] );
tran (\_zy_simnet_tvar_20[1][217] , \_zy_simnet_tvar_20[1].label[208] );
tran (\_zy_simnet_tvar_20[1][216] , \_zy_simnet_tvar_20[1].label[207] );
tran (\_zy_simnet_tvar_20[1][215] , \_zy_simnet_tvar_20[1].label[206] );
tran (\_zy_simnet_tvar_20[1][214] , \_zy_simnet_tvar_20[1].label[205] );
tran (\_zy_simnet_tvar_20[1][213] , \_zy_simnet_tvar_20[1].label[204] );
tran (\_zy_simnet_tvar_20[1][212] , \_zy_simnet_tvar_20[1].label[203] );
tran (\_zy_simnet_tvar_20[1][211] , \_zy_simnet_tvar_20[1].label[202] );
tran (\_zy_simnet_tvar_20[1][210] , \_zy_simnet_tvar_20[1].label[201] );
tran (\_zy_simnet_tvar_20[1][209] , \_zy_simnet_tvar_20[1].label[200] );
tran (\_zy_simnet_tvar_20[1][208] , \_zy_simnet_tvar_20[1].label[199] );
tran (\_zy_simnet_tvar_20[1][207] , \_zy_simnet_tvar_20[1].label[198] );
tran (\_zy_simnet_tvar_20[1][206] , \_zy_simnet_tvar_20[1].label[197] );
tran (\_zy_simnet_tvar_20[1][205] , \_zy_simnet_tvar_20[1].label[196] );
tran (\_zy_simnet_tvar_20[1][204] , \_zy_simnet_tvar_20[1].label[195] );
tran (\_zy_simnet_tvar_20[1][203] , \_zy_simnet_tvar_20[1].label[194] );
tran (\_zy_simnet_tvar_20[1][202] , \_zy_simnet_tvar_20[1].label[193] );
tran (\_zy_simnet_tvar_20[1][201] , \_zy_simnet_tvar_20[1].label[192] );
tran (\_zy_simnet_tvar_20[1][200] , \_zy_simnet_tvar_20[1].label[191] );
tran (\_zy_simnet_tvar_20[1][199] , \_zy_simnet_tvar_20[1].label[190] );
tran (\_zy_simnet_tvar_20[1][198] , \_zy_simnet_tvar_20[1].label[189] );
tran (\_zy_simnet_tvar_20[1][197] , \_zy_simnet_tvar_20[1].label[188] );
tran (\_zy_simnet_tvar_20[1][196] , \_zy_simnet_tvar_20[1].label[187] );
tran (\_zy_simnet_tvar_20[1][195] , \_zy_simnet_tvar_20[1].label[186] );
tran (\_zy_simnet_tvar_20[1][194] , \_zy_simnet_tvar_20[1].label[185] );
tran (\_zy_simnet_tvar_20[1][193] , \_zy_simnet_tvar_20[1].label[184] );
tran (\_zy_simnet_tvar_20[1][192] , \_zy_simnet_tvar_20[1].label[183] );
tran (\_zy_simnet_tvar_20[1][191] , \_zy_simnet_tvar_20[1].label[182] );
tran (\_zy_simnet_tvar_20[1][190] , \_zy_simnet_tvar_20[1].label[181] );
tran (\_zy_simnet_tvar_20[1][189] , \_zy_simnet_tvar_20[1].label[180] );
tran (\_zy_simnet_tvar_20[1][188] , \_zy_simnet_tvar_20[1].label[179] );
tran (\_zy_simnet_tvar_20[1][187] , \_zy_simnet_tvar_20[1].label[178] );
tran (\_zy_simnet_tvar_20[1][186] , \_zy_simnet_tvar_20[1].label[177] );
tran (\_zy_simnet_tvar_20[1][185] , \_zy_simnet_tvar_20[1].label[176] );
tran (\_zy_simnet_tvar_20[1][184] , \_zy_simnet_tvar_20[1].label[175] );
tran (\_zy_simnet_tvar_20[1][183] , \_zy_simnet_tvar_20[1].label[174] );
tran (\_zy_simnet_tvar_20[1][182] , \_zy_simnet_tvar_20[1].label[173] );
tran (\_zy_simnet_tvar_20[1][181] , \_zy_simnet_tvar_20[1].label[172] );
tran (\_zy_simnet_tvar_20[1][180] , \_zy_simnet_tvar_20[1].label[171] );
tran (\_zy_simnet_tvar_20[1][179] , \_zy_simnet_tvar_20[1].label[170] );
tran (\_zy_simnet_tvar_20[1][178] , \_zy_simnet_tvar_20[1].label[169] );
tran (\_zy_simnet_tvar_20[1][177] , \_zy_simnet_tvar_20[1].label[168] );
tran (\_zy_simnet_tvar_20[1][176] , \_zy_simnet_tvar_20[1].label[167] );
tran (\_zy_simnet_tvar_20[1][175] , \_zy_simnet_tvar_20[1].label[166] );
tran (\_zy_simnet_tvar_20[1][174] , \_zy_simnet_tvar_20[1].label[165] );
tran (\_zy_simnet_tvar_20[1][173] , \_zy_simnet_tvar_20[1].label[164] );
tran (\_zy_simnet_tvar_20[1][172] , \_zy_simnet_tvar_20[1].label[163] );
tran (\_zy_simnet_tvar_20[1][171] , \_zy_simnet_tvar_20[1].label[162] );
tran (\_zy_simnet_tvar_20[1][170] , \_zy_simnet_tvar_20[1].label[161] );
tran (\_zy_simnet_tvar_20[1][169] , \_zy_simnet_tvar_20[1].label[160] );
tran (\_zy_simnet_tvar_20[1][168] , \_zy_simnet_tvar_20[1].label[159] );
tran (\_zy_simnet_tvar_20[1][167] , \_zy_simnet_tvar_20[1].label[158] );
tran (\_zy_simnet_tvar_20[1][166] , \_zy_simnet_tvar_20[1].label[157] );
tran (\_zy_simnet_tvar_20[1][165] , \_zy_simnet_tvar_20[1].label[156] );
tran (\_zy_simnet_tvar_20[1][164] , \_zy_simnet_tvar_20[1].label[155] );
tran (\_zy_simnet_tvar_20[1][163] , \_zy_simnet_tvar_20[1].label[154] );
tran (\_zy_simnet_tvar_20[1][162] , \_zy_simnet_tvar_20[1].label[153] );
tran (\_zy_simnet_tvar_20[1][161] , \_zy_simnet_tvar_20[1].label[152] );
tran (\_zy_simnet_tvar_20[1][160] , \_zy_simnet_tvar_20[1].label[151] );
tran (\_zy_simnet_tvar_20[1][159] , \_zy_simnet_tvar_20[1].label[150] );
tran (\_zy_simnet_tvar_20[1][158] , \_zy_simnet_tvar_20[1].label[149] );
tran (\_zy_simnet_tvar_20[1][157] , \_zy_simnet_tvar_20[1].label[148] );
tran (\_zy_simnet_tvar_20[1][156] , \_zy_simnet_tvar_20[1].label[147] );
tran (\_zy_simnet_tvar_20[1][155] , \_zy_simnet_tvar_20[1].label[146] );
tran (\_zy_simnet_tvar_20[1][154] , \_zy_simnet_tvar_20[1].label[145] );
tran (\_zy_simnet_tvar_20[1][153] , \_zy_simnet_tvar_20[1].label[144] );
tran (\_zy_simnet_tvar_20[1][152] , \_zy_simnet_tvar_20[1].label[143] );
tran (\_zy_simnet_tvar_20[1][151] , \_zy_simnet_tvar_20[1].label[142] );
tran (\_zy_simnet_tvar_20[1][150] , \_zy_simnet_tvar_20[1].label[141] );
tran (\_zy_simnet_tvar_20[1][149] , \_zy_simnet_tvar_20[1].label[140] );
tran (\_zy_simnet_tvar_20[1][148] , \_zy_simnet_tvar_20[1].label[139] );
tran (\_zy_simnet_tvar_20[1][147] , \_zy_simnet_tvar_20[1].label[138] );
tran (\_zy_simnet_tvar_20[1][146] , \_zy_simnet_tvar_20[1].label[137] );
tran (\_zy_simnet_tvar_20[1][145] , \_zy_simnet_tvar_20[1].label[136] );
tran (\_zy_simnet_tvar_20[1][144] , \_zy_simnet_tvar_20[1].label[135] );
tran (\_zy_simnet_tvar_20[1][143] , \_zy_simnet_tvar_20[1].label[134] );
tran (\_zy_simnet_tvar_20[1][142] , \_zy_simnet_tvar_20[1].label[133] );
tran (\_zy_simnet_tvar_20[1][141] , \_zy_simnet_tvar_20[1].label[132] );
tran (\_zy_simnet_tvar_20[1][140] , \_zy_simnet_tvar_20[1].label[131] );
tran (\_zy_simnet_tvar_20[1][139] , \_zy_simnet_tvar_20[1].label[130] );
tran (\_zy_simnet_tvar_20[1][138] , \_zy_simnet_tvar_20[1].label[129] );
tran (\_zy_simnet_tvar_20[1][137] , \_zy_simnet_tvar_20[1].label[128] );
tran (\_zy_simnet_tvar_20[1][136] , \_zy_simnet_tvar_20[1].label[127] );
tran (\_zy_simnet_tvar_20[1][135] , \_zy_simnet_tvar_20[1].label[126] );
tran (\_zy_simnet_tvar_20[1][134] , \_zy_simnet_tvar_20[1].label[125] );
tran (\_zy_simnet_tvar_20[1][133] , \_zy_simnet_tvar_20[1].label[124] );
tran (\_zy_simnet_tvar_20[1][132] , \_zy_simnet_tvar_20[1].label[123] );
tran (\_zy_simnet_tvar_20[1][131] , \_zy_simnet_tvar_20[1].label[122] );
tran (\_zy_simnet_tvar_20[1][130] , \_zy_simnet_tvar_20[1].label[121] );
tran (\_zy_simnet_tvar_20[1][129] , \_zy_simnet_tvar_20[1].label[120] );
tran (\_zy_simnet_tvar_20[1][128] , \_zy_simnet_tvar_20[1].label[119] );
tran (\_zy_simnet_tvar_20[1][127] , \_zy_simnet_tvar_20[1].label[118] );
tran (\_zy_simnet_tvar_20[1][126] , \_zy_simnet_tvar_20[1].label[117] );
tran (\_zy_simnet_tvar_20[1][125] , \_zy_simnet_tvar_20[1].label[116] );
tran (\_zy_simnet_tvar_20[1][124] , \_zy_simnet_tvar_20[1].label[115] );
tran (\_zy_simnet_tvar_20[1][123] , \_zy_simnet_tvar_20[1].label[114] );
tran (\_zy_simnet_tvar_20[1][122] , \_zy_simnet_tvar_20[1].label[113] );
tran (\_zy_simnet_tvar_20[1][121] , \_zy_simnet_tvar_20[1].label[112] );
tran (\_zy_simnet_tvar_20[1][120] , \_zy_simnet_tvar_20[1].label[111] );
tran (\_zy_simnet_tvar_20[1][119] , \_zy_simnet_tvar_20[1].label[110] );
tran (\_zy_simnet_tvar_20[1][118] , \_zy_simnet_tvar_20[1].label[109] );
tran (\_zy_simnet_tvar_20[1][117] , \_zy_simnet_tvar_20[1].label[108] );
tran (\_zy_simnet_tvar_20[1][116] , \_zy_simnet_tvar_20[1].label[107] );
tran (\_zy_simnet_tvar_20[1][115] , \_zy_simnet_tvar_20[1].label[106] );
tran (\_zy_simnet_tvar_20[1][114] , \_zy_simnet_tvar_20[1].label[105] );
tran (\_zy_simnet_tvar_20[1][113] , \_zy_simnet_tvar_20[1].label[104] );
tran (\_zy_simnet_tvar_20[1][112] , \_zy_simnet_tvar_20[1].label[103] );
tran (\_zy_simnet_tvar_20[1][111] , \_zy_simnet_tvar_20[1].label[102] );
tran (\_zy_simnet_tvar_20[1][110] , \_zy_simnet_tvar_20[1].label[101] );
tran (\_zy_simnet_tvar_20[1][109] , \_zy_simnet_tvar_20[1].label[100] );
tran (\_zy_simnet_tvar_20[1][108] , \_zy_simnet_tvar_20[1].label[99] );
tran (\_zy_simnet_tvar_20[1][107] , \_zy_simnet_tvar_20[1].label[98] );
tran (\_zy_simnet_tvar_20[1][106] , \_zy_simnet_tvar_20[1].label[97] );
tran (\_zy_simnet_tvar_20[1][105] , \_zy_simnet_tvar_20[1].label[96] );
tran (\_zy_simnet_tvar_20[1][104] , \_zy_simnet_tvar_20[1].label[95] );
tran (\_zy_simnet_tvar_20[1][103] , \_zy_simnet_tvar_20[1].label[94] );
tran (\_zy_simnet_tvar_20[1][102] , \_zy_simnet_tvar_20[1].label[93] );
tran (\_zy_simnet_tvar_20[1][101] , \_zy_simnet_tvar_20[1].label[92] );
tran (\_zy_simnet_tvar_20[1][100] , \_zy_simnet_tvar_20[1].label[91] );
tran (\_zy_simnet_tvar_20[1][99] , \_zy_simnet_tvar_20[1].label[90] );
tran (\_zy_simnet_tvar_20[1][98] , \_zy_simnet_tvar_20[1].label[89] );
tran (\_zy_simnet_tvar_20[1][97] , \_zy_simnet_tvar_20[1].label[88] );
tran (\_zy_simnet_tvar_20[1][96] , \_zy_simnet_tvar_20[1].label[87] );
tran (\_zy_simnet_tvar_20[1][95] , \_zy_simnet_tvar_20[1].label[86] );
tran (\_zy_simnet_tvar_20[1][94] , \_zy_simnet_tvar_20[1].label[85] );
tran (\_zy_simnet_tvar_20[1][93] , \_zy_simnet_tvar_20[1].label[84] );
tran (\_zy_simnet_tvar_20[1][92] , \_zy_simnet_tvar_20[1].label[83] );
tran (\_zy_simnet_tvar_20[1][91] , \_zy_simnet_tvar_20[1].label[82] );
tran (\_zy_simnet_tvar_20[1][90] , \_zy_simnet_tvar_20[1].label[81] );
tran (\_zy_simnet_tvar_20[1][89] , \_zy_simnet_tvar_20[1].label[80] );
tran (\_zy_simnet_tvar_20[1][88] , \_zy_simnet_tvar_20[1].label[79] );
tran (\_zy_simnet_tvar_20[1][87] , \_zy_simnet_tvar_20[1].label[78] );
tran (\_zy_simnet_tvar_20[1][86] , \_zy_simnet_tvar_20[1].label[77] );
tran (\_zy_simnet_tvar_20[1][85] , \_zy_simnet_tvar_20[1].label[76] );
tran (\_zy_simnet_tvar_20[1][84] , \_zy_simnet_tvar_20[1].label[75] );
tran (\_zy_simnet_tvar_20[1][83] , \_zy_simnet_tvar_20[1].label[74] );
tran (\_zy_simnet_tvar_20[1][82] , \_zy_simnet_tvar_20[1].label[73] );
tran (\_zy_simnet_tvar_20[1][81] , \_zy_simnet_tvar_20[1].label[72] );
tran (\_zy_simnet_tvar_20[1][80] , \_zy_simnet_tvar_20[1].label[71] );
tran (\_zy_simnet_tvar_20[1][79] , \_zy_simnet_tvar_20[1].label[70] );
tran (\_zy_simnet_tvar_20[1][78] , \_zy_simnet_tvar_20[1].label[69] );
tran (\_zy_simnet_tvar_20[1][77] , \_zy_simnet_tvar_20[1].label[68] );
tran (\_zy_simnet_tvar_20[1][76] , \_zy_simnet_tvar_20[1].label[67] );
tran (\_zy_simnet_tvar_20[1][75] , \_zy_simnet_tvar_20[1].label[66] );
tran (\_zy_simnet_tvar_20[1][74] , \_zy_simnet_tvar_20[1].label[65] );
tran (\_zy_simnet_tvar_20[1][73] , \_zy_simnet_tvar_20[1].label[64] );
tran (\_zy_simnet_tvar_20[1][72] , \_zy_simnet_tvar_20[1].label[63] );
tran (\_zy_simnet_tvar_20[1][71] , \_zy_simnet_tvar_20[1].label[62] );
tran (\_zy_simnet_tvar_20[1][70] , \_zy_simnet_tvar_20[1].label[61] );
tran (\_zy_simnet_tvar_20[1][69] , \_zy_simnet_tvar_20[1].label[60] );
tran (\_zy_simnet_tvar_20[1][68] , \_zy_simnet_tvar_20[1].label[59] );
tran (\_zy_simnet_tvar_20[1][67] , \_zy_simnet_tvar_20[1].label[58] );
tran (\_zy_simnet_tvar_20[1][66] , \_zy_simnet_tvar_20[1].label[57] );
tran (\_zy_simnet_tvar_20[1][65] , \_zy_simnet_tvar_20[1].label[56] );
tran (\_zy_simnet_tvar_20[1][64] , \_zy_simnet_tvar_20[1].label[55] );
tran (\_zy_simnet_tvar_20[1][63] , \_zy_simnet_tvar_20[1].label[54] );
tran (\_zy_simnet_tvar_20[1][62] , \_zy_simnet_tvar_20[1].label[53] );
tran (\_zy_simnet_tvar_20[1][61] , \_zy_simnet_tvar_20[1].label[52] );
tran (\_zy_simnet_tvar_20[1][60] , \_zy_simnet_tvar_20[1].label[51] );
tran (\_zy_simnet_tvar_20[1][59] , \_zy_simnet_tvar_20[1].label[50] );
tran (\_zy_simnet_tvar_20[1][58] , \_zy_simnet_tvar_20[1].label[49] );
tran (\_zy_simnet_tvar_20[1][57] , \_zy_simnet_tvar_20[1].label[48] );
tran (\_zy_simnet_tvar_20[1][56] , \_zy_simnet_tvar_20[1].label[47] );
tran (\_zy_simnet_tvar_20[1][55] , \_zy_simnet_tvar_20[1].label[46] );
tran (\_zy_simnet_tvar_20[1][54] , \_zy_simnet_tvar_20[1].label[45] );
tran (\_zy_simnet_tvar_20[1][53] , \_zy_simnet_tvar_20[1].label[44] );
tran (\_zy_simnet_tvar_20[1][52] , \_zy_simnet_tvar_20[1].label[43] );
tran (\_zy_simnet_tvar_20[1][51] , \_zy_simnet_tvar_20[1].label[42] );
tran (\_zy_simnet_tvar_20[1][50] , \_zy_simnet_tvar_20[1].label[41] );
tran (\_zy_simnet_tvar_20[1][49] , \_zy_simnet_tvar_20[1].label[40] );
tran (\_zy_simnet_tvar_20[1][48] , \_zy_simnet_tvar_20[1].label[39] );
tran (\_zy_simnet_tvar_20[1][47] , \_zy_simnet_tvar_20[1].label[38] );
tran (\_zy_simnet_tvar_20[1][46] , \_zy_simnet_tvar_20[1].label[37] );
tran (\_zy_simnet_tvar_20[1][45] , \_zy_simnet_tvar_20[1].label[36] );
tran (\_zy_simnet_tvar_20[1][44] , \_zy_simnet_tvar_20[1].label[35] );
tran (\_zy_simnet_tvar_20[1][43] , \_zy_simnet_tvar_20[1].label[34] );
tran (\_zy_simnet_tvar_20[1][42] , \_zy_simnet_tvar_20[1].label[33] );
tran (\_zy_simnet_tvar_20[1][41] , \_zy_simnet_tvar_20[1].label[32] );
tran (\_zy_simnet_tvar_20[1][40] , \_zy_simnet_tvar_20[1].label[31] );
tran (\_zy_simnet_tvar_20[1][39] , \_zy_simnet_tvar_20[1].label[30] );
tran (\_zy_simnet_tvar_20[1][38] , \_zy_simnet_tvar_20[1].label[29] );
tran (\_zy_simnet_tvar_20[1][37] , \_zy_simnet_tvar_20[1].label[28] );
tran (\_zy_simnet_tvar_20[1][36] , \_zy_simnet_tvar_20[1].label[27] );
tran (\_zy_simnet_tvar_20[1][35] , \_zy_simnet_tvar_20[1].label[26] );
tran (\_zy_simnet_tvar_20[1][34] , \_zy_simnet_tvar_20[1].label[25] );
tran (\_zy_simnet_tvar_20[1][33] , \_zy_simnet_tvar_20[1].label[24] );
tran (\_zy_simnet_tvar_20[1][32] , \_zy_simnet_tvar_20[1].label[23] );
tran (\_zy_simnet_tvar_20[1][31] , \_zy_simnet_tvar_20[1].label[22] );
tran (\_zy_simnet_tvar_20[1][30] , \_zy_simnet_tvar_20[1].label[21] );
tran (\_zy_simnet_tvar_20[1][29] , \_zy_simnet_tvar_20[1].label[20] );
tran (\_zy_simnet_tvar_20[1][28] , \_zy_simnet_tvar_20[1].label[19] );
tran (\_zy_simnet_tvar_20[1][27] , \_zy_simnet_tvar_20[1].label[18] );
tran (\_zy_simnet_tvar_20[1][26] , \_zy_simnet_tvar_20[1].label[17] );
tran (\_zy_simnet_tvar_20[1][25] , \_zy_simnet_tvar_20[1].label[16] );
tran (\_zy_simnet_tvar_20[1][24] , \_zy_simnet_tvar_20[1].label[15] );
tran (\_zy_simnet_tvar_20[1][23] , \_zy_simnet_tvar_20[1].label[14] );
tran (\_zy_simnet_tvar_20[1][22] , \_zy_simnet_tvar_20[1].label[13] );
tran (\_zy_simnet_tvar_20[1][21] , \_zy_simnet_tvar_20[1].label[12] );
tran (\_zy_simnet_tvar_20[1][20] , \_zy_simnet_tvar_20[1].label[11] );
tran (\_zy_simnet_tvar_20[1][19] , \_zy_simnet_tvar_20[1].label[10] );
tran (\_zy_simnet_tvar_20[1][18] , \_zy_simnet_tvar_20[1].label[9] );
tran (\_zy_simnet_tvar_20[1][17] , \_zy_simnet_tvar_20[1].label[8] );
tran (\_zy_simnet_tvar_20[1][16] , \_zy_simnet_tvar_20[1].label[7] );
tran (\_zy_simnet_tvar_20[1][15] , \_zy_simnet_tvar_20[1].label[6] );
tran (\_zy_simnet_tvar_20[1][14] , \_zy_simnet_tvar_20[1].label[5] );
tran (\_zy_simnet_tvar_20[1][13] , \_zy_simnet_tvar_20[1].label[4] );
tran (\_zy_simnet_tvar_20[1][12] , \_zy_simnet_tvar_20[1].label[3] );
tran (\_zy_simnet_tvar_20[1][11] , \_zy_simnet_tvar_20[1].label[2] );
tran (\_zy_simnet_tvar_20[1][10] , \_zy_simnet_tvar_20[1].label[1] );
tran (\_zy_simnet_tvar_20[1][9] , \_zy_simnet_tvar_20[1].label[0] );
tran (\_zy_simnet_tvar_20[1][8] , \_zy_simnet_tvar_20[1].delimiter_valid[0] );
tran (\_zy_simnet_tvar_20[1][7] , \_zy_simnet_tvar_20[1].delimiter[7] );
tran (\_zy_simnet_tvar_20[1][6] , \_zy_simnet_tvar_20[1].delimiter[6] );
tran (\_zy_simnet_tvar_20[1][5] , \_zy_simnet_tvar_20[1].delimiter[5] );
tran (\_zy_simnet_tvar_20[1][4] , \_zy_simnet_tvar_20[1].delimiter[4] );
tran (\_zy_simnet_tvar_20[1][3] , \_zy_simnet_tvar_20[1].delimiter[3] );
tran (\_zy_simnet_tvar_20[1][2] , \_zy_simnet_tvar_20[1].delimiter[2] );
tran (\_zy_simnet_tvar_20[1][1] , \_zy_simnet_tvar_20[1].delimiter[1] );
tran (\_zy_simnet_tvar_20[1][0] , \_zy_simnet_tvar_20[1].delimiter[0] );
tran (\_zy_simnet_tvar_20[0][271] , \_zy_simnet_tvar_20[0].guid_size[0] );
tran (\_zy_simnet_tvar_20[0][270] , \_zy_simnet_tvar_20[0].label_size[5] );
tran (\_zy_simnet_tvar_20[0][269] , \_zy_simnet_tvar_20[0].label_size[4] );
tran (\_zy_simnet_tvar_20[0][268] , \_zy_simnet_tvar_20[0].label_size[3] );
tran (\_zy_simnet_tvar_20[0][267] , \_zy_simnet_tvar_20[0].label_size[2] );
tran (\_zy_simnet_tvar_20[0][266] , \_zy_simnet_tvar_20[0].label_size[1] );
tran (\_zy_simnet_tvar_20[0][265] , \_zy_simnet_tvar_20[0].label_size[0] );
tran (\_zy_simnet_tvar_20[0][264] , \_zy_simnet_tvar_20[0].label[255] );
tran (\_zy_simnet_tvar_20[0][263] , \_zy_simnet_tvar_20[0].label[254] );
tran (\_zy_simnet_tvar_20[0][262] , \_zy_simnet_tvar_20[0].label[253] );
tran (\_zy_simnet_tvar_20[0][261] , \_zy_simnet_tvar_20[0].label[252] );
tran (\_zy_simnet_tvar_20[0][260] , \_zy_simnet_tvar_20[0].label[251] );
tran (\_zy_simnet_tvar_20[0][259] , \_zy_simnet_tvar_20[0].label[250] );
tran (\_zy_simnet_tvar_20[0][258] , \_zy_simnet_tvar_20[0].label[249] );
tran (\_zy_simnet_tvar_20[0][257] , \_zy_simnet_tvar_20[0].label[248] );
tran (\_zy_simnet_tvar_20[0][256] , \_zy_simnet_tvar_20[0].label[247] );
tran (\_zy_simnet_tvar_20[0][255] , \_zy_simnet_tvar_20[0].label[246] );
tran (\_zy_simnet_tvar_20[0][254] , \_zy_simnet_tvar_20[0].label[245] );
tran (\_zy_simnet_tvar_20[0][253] , \_zy_simnet_tvar_20[0].label[244] );
tran (\_zy_simnet_tvar_20[0][252] , \_zy_simnet_tvar_20[0].label[243] );
tran (\_zy_simnet_tvar_20[0][251] , \_zy_simnet_tvar_20[0].label[242] );
tran (\_zy_simnet_tvar_20[0][250] , \_zy_simnet_tvar_20[0].label[241] );
tran (\_zy_simnet_tvar_20[0][249] , \_zy_simnet_tvar_20[0].label[240] );
tran (\_zy_simnet_tvar_20[0][248] , \_zy_simnet_tvar_20[0].label[239] );
tran (\_zy_simnet_tvar_20[0][247] , \_zy_simnet_tvar_20[0].label[238] );
tran (\_zy_simnet_tvar_20[0][246] , \_zy_simnet_tvar_20[0].label[237] );
tran (\_zy_simnet_tvar_20[0][245] , \_zy_simnet_tvar_20[0].label[236] );
tran (\_zy_simnet_tvar_20[0][244] , \_zy_simnet_tvar_20[0].label[235] );
tran (\_zy_simnet_tvar_20[0][243] , \_zy_simnet_tvar_20[0].label[234] );
tran (\_zy_simnet_tvar_20[0][242] , \_zy_simnet_tvar_20[0].label[233] );
tran (\_zy_simnet_tvar_20[0][241] , \_zy_simnet_tvar_20[0].label[232] );
tran (\_zy_simnet_tvar_20[0][240] , \_zy_simnet_tvar_20[0].label[231] );
tran (\_zy_simnet_tvar_20[0][239] , \_zy_simnet_tvar_20[0].label[230] );
tran (\_zy_simnet_tvar_20[0][238] , \_zy_simnet_tvar_20[0].label[229] );
tran (\_zy_simnet_tvar_20[0][237] , \_zy_simnet_tvar_20[0].label[228] );
tran (\_zy_simnet_tvar_20[0][236] , \_zy_simnet_tvar_20[0].label[227] );
tran (\_zy_simnet_tvar_20[0][235] , \_zy_simnet_tvar_20[0].label[226] );
tran (\_zy_simnet_tvar_20[0][234] , \_zy_simnet_tvar_20[0].label[225] );
tran (\_zy_simnet_tvar_20[0][233] , \_zy_simnet_tvar_20[0].label[224] );
tran (\_zy_simnet_tvar_20[0][232] , \_zy_simnet_tvar_20[0].label[223] );
tran (\_zy_simnet_tvar_20[0][231] , \_zy_simnet_tvar_20[0].label[222] );
tran (\_zy_simnet_tvar_20[0][230] , \_zy_simnet_tvar_20[0].label[221] );
tran (\_zy_simnet_tvar_20[0][229] , \_zy_simnet_tvar_20[0].label[220] );
tran (\_zy_simnet_tvar_20[0][228] , \_zy_simnet_tvar_20[0].label[219] );
tran (\_zy_simnet_tvar_20[0][227] , \_zy_simnet_tvar_20[0].label[218] );
tran (\_zy_simnet_tvar_20[0][226] , \_zy_simnet_tvar_20[0].label[217] );
tran (\_zy_simnet_tvar_20[0][225] , \_zy_simnet_tvar_20[0].label[216] );
tran (\_zy_simnet_tvar_20[0][224] , \_zy_simnet_tvar_20[0].label[215] );
tran (\_zy_simnet_tvar_20[0][223] , \_zy_simnet_tvar_20[0].label[214] );
tran (\_zy_simnet_tvar_20[0][222] , \_zy_simnet_tvar_20[0].label[213] );
tran (\_zy_simnet_tvar_20[0][221] , \_zy_simnet_tvar_20[0].label[212] );
tran (\_zy_simnet_tvar_20[0][220] , \_zy_simnet_tvar_20[0].label[211] );
tran (\_zy_simnet_tvar_20[0][219] , \_zy_simnet_tvar_20[0].label[210] );
tran (\_zy_simnet_tvar_20[0][218] , \_zy_simnet_tvar_20[0].label[209] );
tran (\_zy_simnet_tvar_20[0][217] , \_zy_simnet_tvar_20[0].label[208] );
tran (\_zy_simnet_tvar_20[0][216] , \_zy_simnet_tvar_20[0].label[207] );
tran (\_zy_simnet_tvar_20[0][215] , \_zy_simnet_tvar_20[0].label[206] );
tran (\_zy_simnet_tvar_20[0][214] , \_zy_simnet_tvar_20[0].label[205] );
tran (\_zy_simnet_tvar_20[0][213] , \_zy_simnet_tvar_20[0].label[204] );
tran (\_zy_simnet_tvar_20[0][212] , \_zy_simnet_tvar_20[0].label[203] );
tran (\_zy_simnet_tvar_20[0][211] , \_zy_simnet_tvar_20[0].label[202] );
tran (\_zy_simnet_tvar_20[0][210] , \_zy_simnet_tvar_20[0].label[201] );
tran (\_zy_simnet_tvar_20[0][209] , \_zy_simnet_tvar_20[0].label[200] );
tran (\_zy_simnet_tvar_20[0][208] , \_zy_simnet_tvar_20[0].label[199] );
tran (\_zy_simnet_tvar_20[0][207] , \_zy_simnet_tvar_20[0].label[198] );
tran (\_zy_simnet_tvar_20[0][206] , \_zy_simnet_tvar_20[0].label[197] );
tran (\_zy_simnet_tvar_20[0][205] , \_zy_simnet_tvar_20[0].label[196] );
tran (\_zy_simnet_tvar_20[0][204] , \_zy_simnet_tvar_20[0].label[195] );
tran (\_zy_simnet_tvar_20[0][203] , \_zy_simnet_tvar_20[0].label[194] );
tran (\_zy_simnet_tvar_20[0][202] , \_zy_simnet_tvar_20[0].label[193] );
tran (\_zy_simnet_tvar_20[0][201] , \_zy_simnet_tvar_20[0].label[192] );
tran (\_zy_simnet_tvar_20[0][200] , \_zy_simnet_tvar_20[0].label[191] );
tran (\_zy_simnet_tvar_20[0][199] , \_zy_simnet_tvar_20[0].label[190] );
tran (\_zy_simnet_tvar_20[0][198] , \_zy_simnet_tvar_20[0].label[189] );
tran (\_zy_simnet_tvar_20[0][197] , \_zy_simnet_tvar_20[0].label[188] );
tran (\_zy_simnet_tvar_20[0][196] , \_zy_simnet_tvar_20[0].label[187] );
tran (\_zy_simnet_tvar_20[0][195] , \_zy_simnet_tvar_20[0].label[186] );
tran (\_zy_simnet_tvar_20[0][194] , \_zy_simnet_tvar_20[0].label[185] );
tran (\_zy_simnet_tvar_20[0][193] , \_zy_simnet_tvar_20[0].label[184] );
tran (\_zy_simnet_tvar_20[0][192] , \_zy_simnet_tvar_20[0].label[183] );
tran (\_zy_simnet_tvar_20[0][191] , \_zy_simnet_tvar_20[0].label[182] );
tran (\_zy_simnet_tvar_20[0][190] , \_zy_simnet_tvar_20[0].label[181] );
tran (\_zy_simnet_tvar_20[0][189] , \_zy_simnet_tvar_20[0].label[180] );
tran (\_zy_simnet_tvar_20[0][188] , \_zy_simnet_tvar_20[0].label[179] );
tran (\_zy_simnet_tvar_20[0][187] , \_zy_simnet_tvar_20[0].label[178] );
tran (\_zy_simnet_tvar_20[0][186] , \_zy_simnet_tvar_20[0].label[177] );
tran (\_zy_simnet_tvar_20[0][185] , \_zy_simnet_tvar_20[0].label[176] );
tran (\_zy_simnet_tvar_20[0][184] , \_zy_simnet_tvar_20[0].label[175] );
tran (\_zy_simnet_tvar_20[0][183] , \_zy_simnet_tvar_20[0].label[174] );
tran (\_zy_simnet_tvar_20[0][182] , \_zy_simnet_tvar_20[0].label[173] );
tran (\_zy_simnet_tvar_20[0][181] , \_zy_simnet_tvar_20[0].label[172] );
tran (\_zy_simnet_tvar_20[0][180] , \_zy_simnet_tvar_20[0].label[171] );
tran (\_zy_simnet_tvar_20[0][179] , \_zy_simnet_tvar_20[0].label[170] );
tran (\_zy_simnet_tvar_20[0][178] , \_zy_simnet_tvar_20[0].label[169] );
tran (\_zy_simnet_tvar_20[0][177] , \_zy_simnet_tvar_20[0].label[168] );
tran (\_zy_simnet_tvar_20[0][176] , \_zy_simnet_tvar_20[0].label[167] );
tran (\_zy_simnet_tvar_20[0][175] , \_zy_simnet_tvar_20[0].label[166] );
tran (\_zy_simnet_tvar_20[0][174] , \_zy_simnet_tvar_20[0].label[165] );
tran (\_zy_simnet_tvar_20[0][173] , \_zy_simnet_tvar_20[0].label[164] );
tran (\_zy_simnet_tvar_20[0][172] , \_zy_simnet_tvar_20[0].label[163] );
tran (\_zy_simnet_tvar_20[0][171] , \_zy_simnet_tvar_20[0].label[162] );
tran (\_zy_simnet_tvar_20[0][170] , \_zy_simnet_tvar_20[0].label[161] );
tran (\_zy_simnet_tvar_20[0][169] , \_zy_simnet_tvar_20[0].label[160] );
tran (\_zy_simnet_tvar_20[0][168] , \_zy_simnet_tvar_20[0].label[159] );
tran (\_zy_simnet_tvar_20[0][167] , \_zy_simnet_tvar_20[0].label[158] );
tran (\_zy_simnet_tvar_20[0][166] , \_zy_simnet_tvar_20[0].label[157] );
tran (\_zy_simnet_tvar_20[0][165] , \_zy_simnet_tvar_20[0].label[156] );
tran (\_zy_simnet_tvar_20[0][164] , \_zy_simnet_tvar_20[0].label[155] );
tran (\_zy_simnet_tvar_20[0][163] , \_zy_simnet_tvar_20[0].label[154] );
tran (\_zy_simnet_tvar_20[0][162] , \_zy_simnet_tvar_20[0].label[153] );
tran (\_zy_simnet_tvar_20[0][161] , \_zy_simnet_tvar_20[0].label[152] );
tran (\_zy_simnet_tvar_20[0][160] , \_zy_simnet_tvar_20[0].label[151] );
tran (\_zy_simnet_tvar_20[0][159] , \_zy_simnet_tvar_20[0].label[150] );
tran (\_zy_simnet_tvar_20[0][158] , \_zy_simnet_tvar_20[0].label[149] );
tran (\_zy_simnet_tvar_20[0][157] , \_zy_simnet_tvar_20[0].label[148] );
tran (\_zy_simnet_tvar_20[0][156] , \_zy_simnet_tvar_20[0].label[147] );
tran (\_zy_simnet_tvar_20[0][155] , \_zy_simnet_tvar_20[0].label[146] );
tran (\_zy_simnet_tvar_20[0][154] , \_zy_simnet_tvar_20[0].label[145] );
tran (\_zy_simnet_tvar_20[0][153] , \_zy_simnet_tvar_20[0].label[144] );
tran (\_zy_simnet_tvar_20[0][152] , \_zy_simnet_tvar_20[0].label[143] );
tran (\_zy_simnet_tvar_20[0][151] , \_zy_simnet_tvar_20[0].label[142] );
tran (\_zy_simnet_tvar_20[0][150] , \_zy_simnet_tvar_20[0].label[141] );
tran (\_zy_simnet_tvar_20[0][149] , \_zy_simnet_tvar_20[0].label[140] );
tran (\_zy_simnet_tvar_20[0][148] , \_zy_simnet_tvar_20[0].label[139] );
tran (\_zy_simnet_tvar_20[0][147] , \_zy_simnet_tvar_20[0].label[138] );
tran (\_zy_simnet_tvar_20[0][146] , \_zy_simnet_tvar_20[0].label[137] );
tran (\_zy_simnet_tvar_20[0][145] , \_zy_simnet_tvar_20[0].label[136] );
tran (\_zy_simnet_tvar_20[0][144] , \_zy_simnet_tvar_20[0].label[135] );
tran (\_zy_simnet_tvar_20[0][143] , \_zy_simnet_tvar_20[0].label[134] );
tran (\_zy_simnet_tvar_20[0][142] , \_zy_simnet_tvar_20[0].label[133] );
tran (\_zy_simnet_tvar_20[0][141] , \_zy_simnet_tvar_20[0].label[132] );
tran (\_zy_simnet_tvar_20[0][140] , \_zy_simnet_tvar_20[0].label[131] );
tran (\_zy_simnet_tvar_20[0][139] , \_zy_simnet_tvar_20[0].label[130] );
tran (\_zy_simnet_tvar_20[0][138] , \_zy_simnet_tvar_20[0].label[129] );
tran (\_zy_simnet_tvar_20[0][137] , \_zy_simnet_tvar_20[0].label[128] );
tran (\_zy_simnet_tvar_20[0][136] , \_zy_simnet_tvar_20[0].label[127] );
tran (\_zy_simnet_tvar_20[0][135] , \_zy_simnet_tvar_20[0].label[126] );
tran (\_zy_simnet_tvar_20[0][134] , \_zy_simnet_tvar_20[0].label[125] );
tran (\_zy_simnet_tvar_20[0][133] , \_zy_simnet_tvar_20[0].label[124] );
tran (\_zy_simnet_tvar_20[0][132] , \_zy_simnet_tvar_20[0].label[123] );
tran (\_zy_simnet_tvar_20[0][131] , \_zy_simnet_tvar_20[0].label[122] );
tran (\_zy_simnet_tvar_20[0][130] , \_zy_simnet_tvar_20[0].label[121] );
tran (\_zy_simnet_tvar_20[0][129] , \_zy_simnet_tvar_20[0].label[120] );
tran (\_zy_simnet_tvar_20[0][128] , \_zy_simnet_tvar_20[0].label[119] );
tran (\_zy_simnet_tvar_20[0][127] , \_zy_simnet_tvar_20[0].label[118] );
tran (\_zy_simnet_tvar_20[0][126] , \_zy_simnet_tvar_20[0].label[117] );
tran (\_zy_simnet_tvar_20[0][125] , \_zy_simnet_tvar_20[0].label[116] );
tran (\_zy_simnet_tvar_20[0][124] , \_zy_simnet_tvar_20[0].label[115] );
tran (\_zy_simnet_tvar_20[0][123] , \_zy_simnet_tvar_20[0].label[114] );
tran (\_zy_simnet_tvar_20[0][122] , \_zy_simnet_tvar_20[0].label[113] );
tran (\_zy_simnet_tvar_20[0][121] , \_zy_simnet_tvar_20[0].label[112] );
tran (\_zy_simnet_tvar_20[0][120] , \_zy_simnet_tvar_20[0].label[111] );
tran (\_zy_simnet_tvar_20[0][119] , \_zy_simnet_tvar_20[0].label[110] );
tran (\_zy_simnet_tvar_20[0][118] , \_zy_simnet_tvar_20[0].label[109] );
tran (\_zy_simnet_tvar_20[0][117] , \_zy_simnet_tvar_20[0].label[108] );
tran (\_zy_simnet_tvar_20[0][116] , \_zy_simnet_tvar_20[0].label[107] );
tran (\_zy_simnet_tvar_20[0][115] , \_zy_simnet_tvar_20[0].label[106] );
tran (\_zy_simnet_tvar_20[0][114] , \_zy_simnet_tvar_20[0].label[105] );
tran (\_zy_simnet_tvar_20[0][113] , \_zy_simnet_tvar_20[0].label[104] );
tran (\_zy_simnet_tvar_20[0][112] , \_zy_simnet_tvar_20[0].label[103] );
tran (\_zy_simnet_tvar_20[0][111] , \_zy_simnet_tvar_20[0].label[102] );
tran (\_zy_simnet_tvar_20[0][110] , \_zy_simnet_tvar_20[0].label[101] );
tran (\_zy_simnet_tvar_20[0][109] , \_zy_simnet_tvar_20[0].label[100] );
tran (\_zy_simnet_tvar_20[0][108] , \_zy_simnet_tvar_20[0].label[99] );
tran (\_zy_simnet_tvar_20[0][107] , \_zy_simnet_tvar_20[0].label[98] );
tran (\_zy_simnet_tvar_20[0][106] , \_zy_simnet_tvar_20[0].label[97] );
tran (\_zy_simnet_tvar_20[0][105] , \_zy_simnet_tvar_20[0].label[96] );
tran (\_zy_simnet_tvar_20[0][104] , \_zy_simnet_tvar_20[0].label[95] );
tran (\_zy_simnet_tvar_20[0][103] , \_zy_simnet_tvar_20[0].label[94] );
tran (\_zy_simnet_tvar_20[0][102] , \_zy_simnet_tvar_20[0].label[93] );
tran (\_zy_simnet_tvar_20[0][101] , \_zy_simnet_tvar_20[0].label[92] );
tran (\_zy_simnet_tvar_20[0][100] , \_zy_simnet_tvar_20[0].label[91] );
tran (\_zy_simnet_tvar_20[0][99] , \_zy_simnet_tvar_20[0].label[90] );
tran (\_zy_simnet_tvar_20[0][98] , \_zy_simnet_tvar_20[0].label[89] );
tran (\_zy_simnet_tvar_20[0][97] , \_zy_simnet_tvar_20[0].label[88] );
tran (\_zy_simnet_tvar_20[0][96] , \_zy_simnet_tvar_20[0].label[87] );
tran (\_zy_simnet_tvar_20[0][95] , \_zy_simnet_tvar_20[0].label[86] );
tran (\_zy_simnet_tvar_20[0][94] , \_zy_simnet_tvar_20[0].label[85] );
tran (\_zy_simnet_tvar_20[0][93] , \_zy_simnet_tvar_20[0].label[84] );
tran (\_zy_simnet_tvar_20[0][92] , \_zy_simnet_tvar_20[0].label[83] );
tran (\_zy_simnet_tvar_20[0][91] , \_zy_simnet_tvar_20[0].label[82] );
tran (\_zy_simnet_tvar_20[0][90] , \_zy_simnet_tvar_20[0].label[81] );
tran (\_zy_simnet_tvar_20[0][89] , \_zy_simnet_tvar_20[0].label[80] );
tran (\_zy_simnet_tvar_20[0][88] , \_zy_simnet_tvar_20[0].label[79] );
tran (\_zy_simnet_tvar_20[0][87] , \_zy_simnet_tvar_20[0].label[78] );
tran (\_zy_simnet_tvar_20[0][86] , \_zy_simnet_tvar_20[0].label[77] );
tran (\_zy_simnet_tvar_20[0][85] , \_zy_simnet_tvar_20[0].label[76] );
tran (\_zy_simnet_tvar_20[0][84] , \_zy_simnet_tvar_20[0].label[75] );
tran (\_zy_simnet_tvar_20[0][83] , \_zy_simnet_tvar_20[0].label[74] );
tran (\_zy_simnet_tvar_20[0][82] , \_zy_simnet_tvar_20[0].label[73] );
tran (\_zy_simnet_tvar_20[0][81] , \_zy_simnet_tvar_20[0].label[72] );
tran (\_zy_simnet_tvar_20[0][80] , \_zy_simnet_tvar_20[0].label[71] );
tran (\_zy_simnet_tvar_20[0][79] , \_zy_simnet_tvar_20[0].label[70] );
tran (\_zy_simnet_tvar_20[0][78] , \_zy_simnet_tvar_20[0].label[69] );
tran (\_zy_simnet_tvar_20[0][77] , \_zy_simnet_tvar_20[0].label[68] );
tran (\_zy_simnet_tvar_20[0][76] , \_zy_simnet_tvar_20[0].label[67] );
tran (\_zy_simnet_tvar_20[0][75] , \_zy_simnet_tvar_20[0].label[66] );
tran (\_zy_simnet_tvar_20[0][74] , \_zy_simnet_tvar_20[0].label[65] );
tran (\_zy_simnet_tvar_20[0][73] , \_zy_simnet_tvar_20[0].label[64] );
tran (\_zy_simnet_tvar_20[0][72] , \_zy_simnet_tvar_20[0].label[63] );
tran (\_zy_simnet_tvar_20[0][71] , \_zy_simnet_tvar_20[0].label[62] );
tran (\_zy_simnet_tvar_20[0][70] , \_zy_simnet_tvar_20[0].label[61] );
tran (\_zy_simnet_tvar_20[0][69] , \_zy_simnet_tvar_20[0].label[60] );
tran (\_zy_simnet_tvar_20[0][68] , \_zy_simnet_tvar_20[0].label[59] );
tran (\_zy_simnet_tvar_20[0][67] , \_zy_simnet_tvar_20[0].label[58] );
tran (\_zy_simnet_tvar_20[0][66] , \_zy_simnet_tvar_20[0].label[57] );
tran (\_zy_simnet_tvar_20[0][65] , \_zy_simnet_tvar_20[0].label[56] );
tran (\_zy_simnet_tvar_20[0][64] , \_zy_simnet_tvar_20[0].label[55] );
tran (\_zy_simnet_tvar_20[0][63] , \_zy_simnet_tvar_20[0].label[54] );
tran (\_zy_simnet_tvar_20[0][62] , \_zy_simnet_tvar_20[0].label[53] );
tran (\_zy_simnet_tvar_20[0][61] , \_zy_simnet_tvar_20[0].label[52] );
tran (\_zy_simnet_tvar_20[0][60] , \_zy_simnet_tvar_20[0].label[51] );
tran (\_zy_simnet_tvar_20[0][59] , \_zy_simnet_tvar_20[0].label[50] );
tran (\_zy_simnet_tvar_20[0][58] , \_zy_simnet_tvar_20[0].label[49] );
tran (\_zy_simnet_tvar_20[0][57] , \_zy_simnet_tvar_20[0].label[48] );
tran (\_zy_simnet_tvar_20[0][56] , \_zy_simnet_tvar_20[0].label[47] );
tran (\_zy_simnet_tvar_20[0][55] , \_zy_simnet_tvar_20[0].label[46] );
tran (\_zy_simnet_tvar_20[0][54] , \_zy_simnet_tvar_20[0].label[45] );
tran (\_zy_simnet_tvar_20[0][53] , \_zy_simnet_tvar_20[0].label[44] );
tran (\_zy_simnet_tvar_20[0][52] , \_zy_simnet_tvar_20[0].label[43] );
tran (\_zy_simnet_tvar_20[0][51] , \_zy_simnet_tvar_20[0].label[42] );
tran (\_zy_simnet_tvar_20[0][50] , \_zy_simnet_tvar_20[0].label[41] );
tran (\_zy_simnet_tvar_20[0][49] , \_zy_simnet_tvar_20[0].label[40] );
tran (\_zy_simnet_tvar_20[0][48] , \_zy_simnet_tvar_20[0].label[39] );
tran (\_zy_simnet_tvar_20[0][47] , \_zy_simnet_tvar_20[0].label[38] );
tran (\_zy_simnet_tvar_20[0][46] , \_zy_simnet_tvar_20[0].label[37] );
tran (\_zy_simnet_tvar_20[0][45] , \_zy_simnet_tvar_20[0].label[36] );
tran (\_zy_simnet_tvar_20[0][44] , \_zy_simnet_tvar_20[0].label[35] );
tran (\_zy_simnet_tvar_20[0][43] , \_zy_simnet_tvar_20[0].label[34] );
tran (\_zy_simnet_tvar_20[0][42] , \_zy_simnet_tvar_20[0].label[33] );
tran (\_zy_simnet_tvar_20[0][41] , \_zy_simnet_tvar_20[0].label[32] );
tran (\_zy_simnet_tvar_20[0][40] , \_zy_simnet_tvar_20[0].label[31] );
tran (\_zy_simnet_tvar_20[0][39] , \_zy_simnet_tvar_20[0].label[30] );
tran (\_zy_simnet_tvar_20[0][38] , \_zy_simnet_tvar_20[0].label[29] );
tran (\_zy_simnet_tvar_20[0][37] , \_zy_simnet_tvar_20[0].label[28] );
tran (\_zy_simnet_tvar_20[0][36] , \_zy_simnet_tvar_20[0].label[27] );
tran (\_zy_simnet_tvar_20[0][35] , \_zy_simnet_tvar_20[0].label[26] );
tran (\_zy_simnet_tvar_20[0][34] , \_zy_simnet_tvar_20[0].label[25] );
tran (\_zy_simnet_tvar_20[0][33] , \_zy_simnet_tvar_20[0].label[24] );
tran (\_zy_simnet_tvar_20[0][32] , \_zy_simnet_tvar_20[0].label[23] );
tran (\_zy_simnet_tvar_20[0][31] , \_zy_simnet_tvar_20[0].label[22] );
tran (\_zy_simnet_tvar_20[0][30] , \_zy_simnet_tvar_20[0].label[21] );
tran (\_zy_simnet_tvar_20[0][29] , \_zy_simnet_tvar_20[0].label[20] );
tran (\_zy_simnet_tvar_20[0][28] , \_zy_simnet_tvar_20[0].label[19] );
tran (\_zy_simnet_tvar_20[0][27] , \_zy_simnet_tvar_20[0].label[18] );
tran (\_zy_simnet_tvar_20[0][26] , \_zy_simnet_tvar_20[0].label[17] );
tran (\_zy_simnet_tvar_20[0][25] , \_zy_simnet_tvar_20[0].label[16] );
tran (\_zy_simnet_tvar_20[0][24] , \_zy_simnet_tvar_20[0].label[15] );
tran (\_zy_simnet_tvar_20[0][23] , \_zy_simnet_tvar_20[0].label[14] );
tran (\_zy_simnet_tvar_20[0][22] , \_zy_simnet_tvar_20[0].label[13] );
tran (\_zy_simnet_tvar_20[0][21] , \_zy_simnet_tvar_20[0].label[12] );
tran (\_zy_simnet_tvar_20[0][20] , \_zy_simnet_tvar_20[0].label[11] );
tran (\_zy_simnet_tvar_20[0][19] , \_zy_simnet_tvar_20[0].label[10] );
tran (\_zy_simnet_tvar_20[0][18] , \_zy_simnet_tvar_20[0].label[9] );
tran (\_zy_simnet_tvar_20[0][17] , \_zy_simnet_tvar_20[0].label[8] );
tran (\_zy_simnet_tvar_20[0][16] , \_zy_simnet_tvar_20[0].label[7] );
tran (\_zy_simnet_tvar_20[0][15] , \_zy_simnet_tvar_20[0].label[6] );
tran (\_zy_simnet_tvar_20[0][14] , \_zy_simnet_tvar_20[0].label[5] );
tran (\_zy_simnet_tvar_20[0][13] , \_zy_simnet_tvar_20[0].label[4] );
tran (\_zy_simnet_tvar_20[0][12] , \_zy_simnet_tvar_20[0].label[3] );
tran (\_zy_simnet_tvar_20[0][11] , \_zy_simnet_tvar_20[0].label[2] );
tran (\_zy_simnet_tvar_20[0][10] , \_zy_simnet_tvar_20[0].label[1] );
tran (\_zy_simnet_tvar_20[0][9] , \_zy_simnet_tvar_20[0].label[0] );
tran (\_zy_simnet_tvar_20[0][8] , \_zy_simnet_tvar_20[0].delimiter_valid[0] );
tran (\_zy_simnet_tvar_20[0][7] , \_zy_simnet_tvar_20[0].delimiter[7] );
tran (\_zy_simnet_tvar_20[0][6] , \_zy_simnet_tvar_20[0].delimiter[6] );
tran (\_zy_simnet_tvar_20[0][5] , \_zy_simnet_tvar_20[0].delimiter[5] );
tran (\_zy_simnet_tvar_20[0][4] , \_zy_simnet_tvar_20[0].delimiter[4] );
tran (\_zy_simnet_tvar_20[0][3] , \_zy_simnet_tvar_20[0].delimiter[3] );
tran (\_zy_simnet_tvar_20[0][2] , \_zy_simnet_tvar_20[0].delimiter[2] );
tran (\_zy_simnet_tvar_20[0][1] , \_zy_simnet_tvar_20[0].delimiter[1] );
tran (\_zy_simnet_tvar_20[0][0] , \_zy_simnet_tvar_20[0].delimiter[0] );
tran (rbus_ring_i[83], \rbus_ring_i.addr [15]);
tran (rbus_ring_i[82], \rbus_ring_i.addr [14]);
tran (rbus_ring_i[81], \rbus_ring_i.addr [13]);
tran (rbus_ring_i[80], \rbus_ring_i.addr [12]);
tran (rbus_ring_i[79], \rbus_ring_i.addr [11]);
tran (rbus_ring_i[78], \rbus_ring_i.addr [10]);
tran (rbus_ring_i[77], \rbus_ring_i.addr [9]);
tran (rbus_ring_i[76], \rbus_ring_i.addr [8]);
tran (rbus_ring_i[75], \rbus_ring_i.addr [7]);
tran (rbus_ring_i[74], \rbus_ring_i.addr [6]);
tran (rbus_ring_i[73], \rbus_ring_i.addr [5]);
tran (rbus_ring_i[72], \rbus_ring_i.addr [4]);
tran (rbus_ring_i[71], \rbus_ring_i.addr [3]);
tran (rbus_ring_i[70], \rbus_ring_i.addr [2]);
tran (rbus_ring_i[69], \rbus_ring_i.addr [1]);
tran (rbus_ring_i[68], \rbus_ring_i.addr [0]);
tran (rbus_ring_i[67], \rbus_ring_i.wr_strb );
tran (rbus_ring_i[66], \rbus_ring_i.wr_data [31]);
tran (rbus_ring_i[65], \rbus_ring_i.wr_data [30]);
tran (rbus_ring_i[64], \rbus_ring_i.wr_data [29]);
tran (rbus_ring_i[63], \rbus_ring_i.wr_data [28]);
tran (rbus_ring_i[62], \rbus_ring_i.wr_data [27]);
tran (rbus_ring_i[61], \rbus_ring_i.wr_data [26]);
tran (rbus_ring_i[60], \rbus_ring_i.wr_data [25]);
tran (rbus_ring_i[59], \rbus_ring_i.wr_data [24]);
tran (rbus_ring_i[58], \rbus_ring_i.wr_data [23]);
tran (rbus_ring_i[57], \rbus_ring_i.wr_data [22]);
tran (rbus_ring_i[56], \rbus_ring_i.wr_data [21]);
tran (rbus_ring_i[55], \rbus_ring_i.wr_data [20]);
tran (rbus_ring_i[54], \rbus_ring_i.wr_data [19]);
tran (rbus_ring_i[53], \rbus_ring_i.wr_data [18]);
tran (rbus_ring_i[52], \rbus_ring_i.wr_data [17]);
tran (rbus_ring_i[51], \rbus_ring_i.wr_data [16]);
tran (rbus_ring_i[50], \rbus_ring_i.wr_data [15]);
tran (rbus_ring_i[49], \rbus_ring_i.wr_data [14]);
tran (rbus_ring_i[48], \rbus_ring_i.wr_data [13]);
tran (rbus_ring_i[47], \rbus_ring_i.wr_data [12]);
tran (rbus_ring_i[46], \rbus_ring_i.wr_data [11]);
tran (rbus_ring_i[45], \rbus_ring_i.wr_data [10]);
tran (rbus_ring_i[44], \rbus_ring_i.wr_data [9]);
tran (rbus_ring_i[43], \rbus_ring_i.wr_data [8]);
tran (rbus_ring_i[42], \rbus_ring_i.wr_data [7]);
tran (rbus_ring_i[41], \rbus_ring_i.wr_data [6]);
tran (rbus_ring_i[40], \rbus_ring_i.wr_data [5]);
tran (rbus_ring_i[39], \rbus_ring_i.wr_data [4]);
tran (rbus_ring_i[38], \rbus_ring_i.wr_data [3]);
tran (rbus_ring_i[37], \rbus_ring_i.wr_data [2]);
tran (rbus_ring_i[36], \rbus_ring_i.wr_data [1]);
tran (rbus_ring_i[35], \rbus_ring_i.wr_data [0]);
tran (rbus_ring_i[34], \rbus_ring_i.rd_strb );
tran (rbus_ring_o[83], \rbus_ring_o.addr [15]);
tran (rbus_ring_o[82], \rbus_ring_o.addr [14]);
tran (rbus_ring_o[81], \rbus_ring_o.addr [13]);
tran (rbus_ring_o[80], \rbus_ring_o.addr [12]);
tran (rbus_ring_o[79], \rbus_ring_o.addr [11]);
tran (rbus_ring_o[78], \rbus_ring_o.addr [10]);
tran (rbus_ring_o[77], \rbus_ring_o.addr [9]);
tran (rbus_ring_o[76], \rbus_ring_o.addr [8]);
tran (rbus_ring_o[75], \rbus_ring_o.addr [7]);
tran (rbus_ring_o[74], \rbus_ring_o.addr [6]);
tran (rbus_ring_o[73], \rbus_ring_o.addr [5]);
tran (rbus_ring_o[72], \rbus_ring_o.addr [4]);
tran (rbus_ring_o[71], \rbus_ring_o.addr [3]);
tran (rbus_ring_o[70], \rbus_ring_o.addr [2]);
tran (rbus_ring_o[69], \rbus_ring_o.addr [1]);
tran (rbus_ring_o[68], \rbus_ring_o.addr [0]);
tran (rbus_ring_o[67], \rbus_ring_o.wr_strb );
tran (rbus_ring_o[66], \rbus_ring_o.wr_data [31]);
tran (rbus_ring_o[65], \rbus_ring_o.wr_data [30]);
tran (rbus_ring_o[64], \rbus_ring_o.wr_data [29]);
tran (rbus_ring_o[63], \rbus_ring_o.wr_data [28]);
tran (rbus_ring_o[62], \rbus_ring_o.wr_data [27]);
tran (rbus_ring_o[61], \rbus_ring_o.wr_data [26]);
tran (rbus_ring_o[60], \rbus_ring_o.wr_data [25]);
tran (rbus_ring_o[59], \rbus_ring_o.wr_data [24]);
tran (rbus_ring_o[58], \rbus_ring_o.wr_data [23]);
tran (rbus_ring_o[57], \rbus_ring_o.wr_data [22]);
tran (rbus_ring_o[56], \rbus_ring_o.wr_data [21]);
tran (rbus_ring_o[55], \rbus_ring_o.wr_data [20]);
tran (rbus_ring_o[54], \rbus_ring_o.wr_data [19]);
tran (rbus_ring_o[53], \rbus_ring_o.wr_data [18]);
tran (rbus_ring_o[52], \rbus_ring_o.wr_data [17]);
tran (rbus_ring_o[51], \rbus_ring_o.wr_data [16]);
tran (rbus_ring_o[50], \rbus_ring_o.wr_data [15]);
tran (rbus_ring_o[49], \rbus_ring_o.wr_data [14]);
tran (rbus_ring_o[48], \rbus_ring_o.wr_data [13]);
tran (rbus_ring_o[47], \rbus_ring_o.wr_data [12]);
tran (rbus_ring_o[46], \rbus_ring_o.wr_data [11]);
tran (rbus_ring_o[45], \rbus_ring_o.wr_data [10]);
tran (rbus_ring_o[44], \rbus_ring_o.wr_data [9]);
tran (rbus_ring_o[43], \rbus_ring_o.wr_data [8]);
tran (rbus_ring_o[42], \rbus_ring_o.wr_data [7]);
tran (rbus_ring_o[41], \rbus_ring_o.wr_data [6]);
tran (rbus_ring_o[40], \rbus_ring_o.wr_data [5]);
tran (rbus_ring_o[39], \rbus_ring_o.wr_data [4]);
tran (rbus_ring_o[38], \rbus_ring_o.wr_data [3]);
tran (rbus_ring_o[37], \rbus_ring_o.wr_data [2]);
tran (rbus_ring_o[36], \rbus_ring_o.wr_data [1]);
tran (rbus_ring_o[35], \rbus_ring_o.wr_data [0]);
tran (rbus_ring_o[34], \rbus_ring_o.rd_strb );
tran (rbus_ring_o[33], \rbus_ring_o.rd_data [31]);
tran (rbus_ring_o[32], \rbus_ring_o.rd_data [30]);
tran (rbus_ring_o[31], \rbus_ring_o.rd_data [29]);
tran (rbus_ring_o[30], \rbus_ring_o.rd_data [28]);
tran (rbus_ring_o[29], \rbus_ring_o.rd_data [27]);
tran (rbus_ring_o[28], \rbus_ring_o.rd_data [26]);
tran (rbus_ring_o[27], \rbus_ring_o.rd_data [25]);
tran (rbus_ring_o[26], \rbus_ring_o.rd_data [24]);
tran (rbus_ring_o[25], \rbus_ring_o.rd_data [23]);
tran (rbus_ring_o[24], \rbus_ring_o.rd_data [22]);
tran (rbus_ring_o[23], \rbus_ring_o.rd_data [21]);
tran (rbus_ring_o[22], \rbus_ring_o.rd_data [20]);
tran (rbus_ring_o[21], \rbus_ring_o.rd_data [19]);
tran (rbus_ring_o[20], \rbus_ring_o.rd_data [18]);
tran (rbus_ring_o[19], \rbus_ring_o.rd_data [17]);
tran (rbus_ring_o[18], \rbus_ring_o.rd_data [16]);
tran (rbus_ring_o[17], \rbus_ring_o.rd_data [15]);
tran (rbus_ring_o[16], \rbus_ring_o.rd_data [14]);
tran (rbus_ring_o[15], \rbus_ring_o.rd_data [13]);
tran (rbus_ring_o[14], \rbus_ring_o.rd_data [12]);
tran (rbus_ring_o[13], \rbus_ring_o.rd_data [11]);
tran (rbus_ring_o[12], \rbus_ring_o.rd_data [10]);
tran (rbus_ring_o[11], \rbus_ring_o.rd_data [9]);
tran (rbus_ring_o[10], \rbus_ring_o.rd_data [8]);
tran (rbus_ring_o[9], \rbus_ring_o.rd_data [7]);
tran (rbus_ring_o[8], \rbus_ring_o.rd_data [6]);
tran (rbus_ring_o[7], \rbus_ring_o.rd_data [5]);
tran (rbus_ring_o[6], \rbus_ring_o.rd_data [4]);
tran (rbus_ring_o[5], \rbus_ring_o.rd_data [3]);
tran (rbus_ring_o[4], \rbus_ring_o.rd_data [2]);
tran (rbus_ring_o[3], \rbus_ring_o.rd_data [1]);
tran (rbus_ring_o[2], \rbus_ring_o.rd_data [0]);
tran (rbus_ring_o[1], \rbus_ring_o.ack );
tran (rbus_ring_o[0], \rbus_ring_o.err_ack );
tran (kme_cceip0_ob_out[82], \kme_cceip0_ob_out.tvalid );
tran (kme_cceip0_ob_out[81], \kme_cceip0_ob_out.tlast );
tran (kme_cceip0_ob_out[80], \kme_cceip0_ob_out.tid [0]);
tran (kme_cceip0_ob_out[79], \kme_cceip0_ob_out.tstrb [7]);
tran (kme_cceip0_ob_out[78], \kme_cceip0_ob_out.tstrb [6]);
tran (kme_cceip0_ob_out[77], \kme_cceip0_ob_out.tstrb [5]);
tran (kme_cceip0_ob_out[76], \kme_cceip0_ob_out.tstrb [4]);
tran (kme_cceip0_ob_out[75], \kme_cceip0_ob_out.tstrb [3]);
tran (kme_cceip0_ob_out[74], \kme_cceip0_ob_out.tstrb [2]);
tran (kme_cceip0_ob_out[73], \kme_cceip0_ob_out.tstrb [1]);
tran (kme_cceip0_ob_out[72], \kme_cceip0_ob_out.tstrb [0]);
tran (kme_cceip0_ob_out[71], \kme_cceip0_ob_out.tuser [7]);
tran (kme_cceip0_ob_out[70], \kme_cceip0_ob_out.tuser [6]);
tran (kme_cceip0_ob_out[69], \kme_cceip0_ob_out.tuser [5]);
tran (kme_cceip0_ob_out[68], \kme_cceip0_ob_out.tuser [4]);
tran (kme_cceip0_ob_out[67], \kme_cceip0_ob_out.tuser [3]);
tran (kme_cceip0_ob_out[66], \kme_cceip0_ob_out.tuser [2]);
tran (kme_cceip0_ob_out[65], \kme_cceip0_ob_out.tuser [1]);
tran (kme_cceip0_ob_out[64], \kme_cceip0_ob_out.tuser [0]);
tran (kme_cceip0_ob_out[63], \kme_cceip0_ob_out.tdata [63]);
tran (kme_cceip0_ob_out[62], \kme_cceip0_ob_out.tdata [62]);
tran (kme_cceip0_ob_out[61], \kme_cceip0_ob_out.tdata [61]);
tran (kme_cceip0_ob_out[60], \kme_cceip0_ob_out.tdata [60]);
tran (kme_cceip0_ob_out[59], \kme_cceip0_ob_out.tdata [59]);
tran (kme_cceip0_ob_out[58], \kme_cceip0_ob_out.tdata [58]);
tran (kme_cceip0_ob_out[57], \kme_cceip0_ob_out.tdata [57]);
tran (kme_cceip0_ob_out[56], \kme_cceip0_ob_out.tdata [56]);
tran (kme_cceip0_ob_out[55], \kme_cceip0_ob_out.tdata [55]);
tran (kme_cceip0_ob_out[54], \kme_cceip0_ob_out.tdata [54]);
tran (kme_cceip0_ob_out[53], \kme_cceip0_ob_out.tdata [53]);
tran (kme_cceip0_ob_out[52], \kme_cceip0_ob_out.tdata [52]);
tran (kme_cceip0_ob_out[51], \kme_cceip0_ob_out.tdata [51]);
tran (kme_cceip0_ob_out[50], \kme_cceip0_ob_out.tdata [50]);
tran (kme_cceip0_ob_out[49], \kme_cceip0_ob_out.tdata [49]);
tran (kme_cceip0_ob_out[48], \kme_cceip0_ob_out.tdata [48]);
tran (kme_cceip0_ob_out[47], \kme_cceip0_ob_out.tdata [47]);
tran (kme_cceip0_ob_out[46], \kme_cceip0_ob_out.tdata [46]);
tran (kme_cceip0_ob_out[45], \kme_cceip0_ob_out.tdata [45]);
tran (kme_cceip0_ob_out[44], \kme_cceip0_ob_out.tdata [44]);
tran (kme_cceip0_ob_out[43], \kme_cceip0_ob_out.tdata [43]);
tran (kme_cceip0_ob_out[42], \kme_cceip0_ob_out.tdata [42]);
tran (kme_cceip0_ob_out[41], \kme_cceip0_ob_out.tdata [41]);
tran (kme_cceip0_ob_out[40], \kme_cceip0_ob_out.tdata [40]);
tran (kme_cceip0_ob_out[39], \kme_cceip0_ob_out.tdata [39]);
tran (kme_cceip0_ob_out[38], \kme_cceip0_ob_out.tdata [38]);
tran (kme_cceip0_ob_out[37], \kme_cceip0_ob_out.tdata [37]);
tran (kme_cceip0_ob_out[36], \kme_cceip0_ob_out.tdata [36]);
tran (kme_cceip0_ob_out[35], \kme_cceip0_ob_out.tdata [35]);
tran (kme_cceip0_ob_out[34], \kme_cceip0_ob_out.tdata [34]);
tran (kme_cceip0_ob_out[33], \kme_cceip0_ob_out.tdata [33]);
tran (kme_cceip0_ob_out[32], \kme_cceip0_ob_out.tdata [32]);
tran (kme_cceip0_ob_out[31], \kme_cceip0_ob_out.tdata [31]);
tran (kme_cceip0_ob_out[30], \kme_cceip0_ob_out.tdata [30]);
tran (kme_cceip0_ob_out[29], \kme_cceip0_ob_out.tdata [29]);
tran (kme_cceip0_ob_out[28], \kme_cceip0_ob_out.tdata [28]);
tran (kme_cceip0_ob_out[27], \kme_cceip0_ob_out.tdata [27]);
tran (kme_cceip0_ob_out[26], \kme_cceip0_ob_out.tdata [26]);
tran (kme_cceip0_ob_out[25], \kme_cceip0_ob_out.tdata [25]);
tran (kme_cceip0_ob_out[24], \kme_cceip0_ob_out.tdata [24]);
tran (kme_cceip0_ob_out[23], \kme_cceip0_ob_out.tdata [23]);
tran (kme_cceip0_ob_out[22], \kme_cceip0_ob_out.tdata [22]);
tran (kme_cceip0_ob_out[21], \kme_cceip0_ob_out.tdata [21]);
tran (kme_cceip0_ob_out[20], \kme_cceip0_ob_out.tdata [20]);
tran (kme_cceip0_ob_out[19], \kme_cceip0_ob_out.tdata [19]);
tran (kme_cceip0_ob_out[18], \kme_cceip0_ob_out.tdata [18]);
tran (kme_cceip0_ob_out[17], \kme_cceip0_ob_out.tdata [17]);
tran (kme_cceip0_ob_out[16], \kme_cceip0_ob_out.tdata [16]);
tran (kme_cceip0_ob_out[15], \kme_cceip0_ob_out.tdata [15]);
tran (kme_cceip0_ob_out[14], \kme_cceip0_ob_out.tdata [14]);
tran (kme_cceip0_ob_out[13], \kme_cceip0_ob_out.tdata [13]);
tran (kme_cceip0_ob_out[12], \kme_cceip0_ob_out.tdata [12]);
tran (kme_cceip0_ob_out[11], \kme_cceip0_ob_out.tdata [11]);
tran (kme_cceip0_ob_out[10], \kme_cceip0_ob_out.tdata [10]);
tran (kme_cceip0_ob_out[9], \kme_cceip0_ob_out.tdata [9]);
tran (kme_cceip0_ob_out[8], \kme_cceip0_ob_out.tdata [8]);
tran (kme_cceip0_ob_out[7], \kme_cceip0_ob_out.tdata [7]);
tran (kme_cceip0_ob_out[6], \kme_cceip0_ob_out.tdata [6]);
tran (kme_cceip0_ob_out[5], \kme_cceip0_ob_out.tdata [5]);
tran (kme_cceip0_ob_out[4], \kme_cceip0_ob_out.tdata [4]);
tran (kme_cceip0_ob_out[3], \kme_cceip0_ob_out.tdata [3]);
tran (kme_cceip0_ob_out[2], \kme_cceip0_ob_out.tdata [2]);
tran (kme_cceip0_ob_out[1], \kme_cceip0_ob_out.tdata [1]);
tran (kme_cceip0_ob_out[0], \kme_cceip0_ob_out.tdata [0]);
tran (kme_cceip0_ob_in_mod[0], \kme_cceip0_ob_in_mod.tready );
tran (kme_cceip1_ob_out[82], \kme_cceip1_ob_out.tvalid );
tran (kme_cceip1_ob_out[81], \kme_cceip1_ob_out.tlast );
tran (kme_cceip1_ob_out[80], \kme_cceip1_ob_out.tid [0]);
tran (kme_cceip1_ob_out[79], \kme_cceip1_ob_out.tstrb [7]);
tran (kme_cceip1_ob_out[78], \kme_cceip1_ob_out.tstrb [6]);
tran (kme_cceip1_ob_out[77], \kme_cceip1_ob_out.tstrb [5]);
tran (kme_cceip1_ob_out[76], \kme_cceip1_ob_out.tstrb [4]);
tran (kme_cceip1_ob_out[75], \kme_cceip1_ob_out.tstrb [3]);
tran (kme_cceip1_ob_out[74], \kme_cceip1_ob_out.tstrb [2]);
tran (kme_cceip1_ob_out[73], \kme_cceip1_ob_out.tstrb [1]);
tran (kme_cceip1_ob_out[72], \kme_cceip1_ob_out.tstrb [0]);
tran (kme_cceip1_ob_out[71], \kme_cceip1_ob_out.tuser [7]);
tran (kme_cceip1_ob_out[70], \kme_cceip1_ob_out.tuser [6]);
tran (kme_cceip1_ob_out[69], \kme_cceip1_ob_out.tuser [5]);
tran (kme_cceip1_ob_out[68], \kme_cceip1_ob_out.tuser [4]);
tran (kme_cceip1_ob_out[67], \kme_cceip1_ob_out.tuser [3]);
tran (kme_cceip1_ob_out[66], \kme_cceip1_ob_out.tuser [2]);
tran (kme_cceip1_ob_out[65], \kme_cceip1_ob_out.tuser [1]);
tran (kme_cceip1_ob_out[64], \kme_cceip1_ob_out.tuser [0]);
tran (kme_cceip1_ob_out[63], \kme_cceip1_ob_out.tdata [63]);
tran (kme_cceip1_ob_out[62], \kme_cceip1_ob_out.tdata [62]);
tran (kme_cceip1_ob_out[61], \kme_cceip1_ob_out.tdata [61]);
tran (kme_cceip1_ob_out[60], \kme_cceip1_ob_out.tdata [60]);
tran (kme_cceip1_ob_out[59], \kme_cceip1_ob_out.tdata [59]);
tran (kme_cceip1_ob_out[58], \kme_cceip1_ob_out.tdata [58]);
tran (kme_cceip1_ob_out[57], \kme_cceip1_ob_out.tdata [57]);
tran (kme_cceip1_ob_out[56], \kme_cceip1_ob_out.tdata [56]);
tran (kme_cceip1_ob_out[55], \kme_cceip1_ob_out.tdata [55]);
tran (kme_cceip1_ob_out[54], \kme_cceip1_ob_out.tdata [54]);
tran (kme_cceip1_ob_out[53], \kme_cceip1_ob_out.tdata [53]);
tran (kme_cceip1_ob_out[52], \kme_cceip1_ob_out.tdata [52]);
tran (kme_cceip1_ob_out[51], \kme_cceip1_ob_out.tdata [51]);
tran (kme_cceip1_ob_out[50], \kme_cceip1_ob_out.tdata [50]);
tran (kme_cceip1_ob_out[49], \kme_cceip1_ob_out.tdata [49]);
tran (kme_cceip1_ob_out[48], \kme_cceip1_ob_out.tdata [48]);
tran (kme_cceip1_ob_out[47], \kme_cceip1_ob_out.tdata [47]);
tran (kme_cceip1_ob_out[46], \kme_cceip1_ob_out.tdata [46]);
tran (kme_cceip1_ob_out[45], \kme_cceip1_ob_out.tdata [45]);
tran (kme_cceip1_ob_out[44], \kme_cceip1_ob_out.tdata [44]);
tran (kme_cceip1_ob_out[43], \kme_cceip1_ob_out.tdata [43]);
tran (kme_cceip1_ob_out[42], \kme_cceip1_ob_out.tdata [42]);
tran (kme_cceip1_ob_out[41], \kme_cceip1_ob_out.tdata [41]);
tran (kme_cceip1_ob_out[40], \kme_cceip1_ob_out.tdata [40]);
tran (kme_cceip1_ob_out[39], \kme_cceip1_ob_out.tdata [39]);
tran (kme_cceip1_ob_out[38], \kme_cceip1_ob_out.tdata [38]);
tran (kme_cceip1_ob_out[37], \kme_cceip1_ob_out.tdata [37]);
tran (kme_cceip1_ob_out[36], \kme_cceip1_ob_out.tdata [36]);
tran (kme_cceip1_ob_out[35], \kme_cceip1_ob_out.tdata [35]);
tran (kme_cceip1_ob_out[34], \kme_cceip1_ob_out.tdata [34]);
tran (kme_cceip1_ob_out[33], \kme_cceip1_ob_out.tdata [33]);
tran (kme_cceip1_ob_out[32], \kme_cceip1_ob_out.tdata [32]);
tran (kme_cceip1_ob_out[31], \kme_cceip1_ob_out.tdata [31]);
tran (kme_cceip1_ob_out[30], \kme_cceip1_ob_out.tdata [30]);
tran (kme_cceip1_ob_out[29], \kme_cceip1_ob_out.tdata [29]);
tran (kme_cceip1_ob_out[28], \kme_cceip1_ob_out.tdata [28]);
tran (kme_cceip1_ob_out[27], \kme_cceip1_ob_out.tdata [27]);
tran (kme_cceip1_ob_out[26], \kme_cceip1_ob_out.tdata [26]);
tran (kme_cceip1_ob_out[25], \kme_cceip1_ob_out.tdata [25]);
tran (kme_cceip1_ob_out[24], \kme_cceip1_ob_out.tdata [24]);
tran (kme_cceip1_ob_out[23], \kme_cceip1_ob_out.tdata [23]);
tran (kme_cceip1_ob_out[22], \kme_cceip1_ob_out.tdata [22]);
tran (kme_cceip1_ob_out[21], \kme_cceip1_ob_out.tdata [21]);
tran (kme_cceip1_ob_out[20], \kme_cceip1_ob_out.tdata [20]);
tran (kme_cceip1_ob_out[19], \kme_cceip1_ob_out.tdata [19]);
tran (kme_cceip1_ob_out[18], \kme_cceip1_ob_out.tdata [18]);
tran (kme_cceip1_ob_out[17], \kme_cceip1_ob_out.tdata [17]);
tran (kme_cceip1_ob_out[16], \kme_cceip1_ob_out.tdata [16]);
tran (kme_cceip1_ob_out[15], \kme_cceip1_ob_out.tdata [15]);
tran (kme_cceip1_ob_out[14], \kme_cceip1_ob_out.tdata [14]);
tran (kme_cceip1_ob_out[13], \kme_cceip1_ob_out.tdata [13]);
tran (kme_cceip1_ob_out[12], \kme_cceip1_ob_out.tdata [12]);
tran (kme_cceip1_ob_out[11], \kme_cceip1_ob_out.tdata [11]);
tran (kme_cceip1_ob_out[10], \kme_cceip1_ob_out.tdata [10]);
tran (kme_cceip1_ob_out[9], \kme_cceip1_ob_out.tdata [9]);
tran (kme_cceip1_ob_out[8], \kme_cceip1_ob_out.tdata [8]);
tran (kme_cceip1_ob_out[7], \kme_cceip1_ob_out.tdata [7]);
tran (kme_cceip1_ob_out[6], \kme_cceip1_ob_out.tdata [6]);
tran (kme_cceip1_ob_out[5], \kme_cceip1_ob_out.tdata [5]);
tran (kme_cceip1_ob_out[4], \kme_cceip1_ob_out.tdata [4]);
tran (kme_cceip1_ob_out[3], \kme_cceip1_ob_out.tdata [3]);
tran (kme_cceip1_ob_out[2], \kme_cceip1_ob_out.tdata [2]);
tran (kme_cceip1_ob_out[1], \kme_cceip1_ob_out.tdata [1]);
tran (kme_cceip1_ob_out[0], \kme_cceip1_ob_out.tdata [0]);
tran (kme_cceip1_ob_in_mod[0], \kme_cceip1_ob_in_mod.tready );
tran (kme_cceip2_ob_out[82], \kme_cceip2_ob_out.tvalid );
tran (kme_cceip2_ob_out[81], \kme_cceip2_ob_out.tlast );
tran (kme_cceip2_ob_out[80], \kme_cceip2_ob_out.tid [0]);
tran (kme_cceip2_ob_out[79], \kme_cceip2_ob_out.tstrb [7]);
tran (kme_cceip2_ob_out[78], \kme_cceip2_ob_out.tstrb [6]);
tran (kme_cceip2_ob_out[77], \kme_cceip2_ob_out.tstrb [5]);
tran (kme_cceip2_ob_out[76], \kme_cceip2_ob_out.tstrb [4]);
tran (kme_cceip2_ob_out[75], \kme_cceip2_ob_out.tstrb [3]);
tran (kme_cceip2_ob_out[74], \kme_cceip2_ob_out.tstrb [2]);
tran (kme_cceip2_ob_out[73], \kme_cceip2_ob_out.tstrb [1]);
tran (kme_cceip2_ob_out[72], \kme_cceip2_ob_out.tstrb [0]);
tran (kme_cceip2_ob_out[71], \kme_cceip2_ob_out.tuser [7]);
tran (kme_cceip2_ob_out[70], \kme_cceip2_ob_out.tuser [6]);
tran (kme_cceip2_ob_out[69], \kme_cceip2_ob_out.tuser [5]);
tran (kme_cceip2_ob_out[68], \kme_cceip2_ob_out.tuser [4]);
tran (kme_cceip2_ob_out[67], \kme_cceip2_ob_out.tuser [3]);
tran (kme_cceip2_ob_out[66], \kme_cceip2_ob_out.tuser [2]);
tran (kme_cceip2_ob_out[65], \kme_cceip2_ob_out.tuser [1]);
tran (kme_cceip2_ob_out[64], \kme_cceip2_ob_out.tuser [0]);
tran (kme_cceip2_ob_out[63], \kme_cceip2_ob_out.tdata [63]);
tran (kme_cceip2_ob_out[62], \kme_cceip2_ob_out.tdata [62]);
tran (kme_cceip2_ob_out[61], \kme_cceip2_ob_out.tdata [61]);
tran (kme_cceip2_ob_out[60], \kme_cceip2_ob_out.tdata [60]);
tran (kme_cceip2_ob_out[59], \kme_cceip2_ob_out.tdata [59]);
tran (kme_cceip2_ob_out[58], \kme_cceip2_ob_out.tdata [58]);
tran (kme_cceip2_ob_out[57], \kme_cceip2_ob_out.tdata [57]);
tran (kme_cceip2_ob_out[56], \kme_cceip2_ob_out.tdata [56]);
tran (kme_cceip2_ob_out[55], \kme_cceip2_ob_out.tdata [55]);
tran (kme_cceip2_ob_out[54], \kme_cceip2_ob_out.tdata [54]);
tran (kme_cceip2_ob_out[53], \kme_cceip2_ob_out.tdata [53]);
tran (kme_cceip2_ob_out[52], \kme_cceip2_ob_out.tdata [52]);
tran (kme_cceip2_ob_out[51], \kme_cceip2_ob_out.tdata [51]);
tran (kme_cceip2_ob_out[50], \kme_cceip2_ob_out.tdata [50]);
tran (kme_cceip2_ob_out[49], \kme_cceip2_ob_out.tdata [49]);
tran (kme_cceip2_ob_out[48], \kme_cceip2_ob_out.tdata [48]);
tran (kme_cceip2_ob_out[47], \kme_cceip2_ob_out.tdata [47]);
tran (kme_cceip2_ob_out[46], \kme_cceip2_ob_out.tdata [46]);
tran (kme_cceip2_ob_out[45], \kme_cceip2_ob_out.tdata [45]);
tran (kme_cceip2_ob_out[44], \kme_cceip2_ob_out.tdata [44]);
tran (kme_cceip2_ob_out[43], \kme_cceip2_ob_out.tdata [43]);
tran (kme_cceip2_ob_out[42], \kme_cceip2_ob_out.tdata [42]);
tran (kme_cceip2_ob_out[41], \kme_cceip2_ob_out.tdata [41]);
tran (kme_cceip2_ob_out[40], \kme_cceip2_ob_out.tdata [40]);
tran (kme_cceip2_ob_out[39], \kme_cceip2_ob_out.tdata [39]);
tran (kme_cceip2_ob_out[38], \kme_cceip2_ob_out.tdata [38]);
tran (kme_cceip2_ob_out[37], \kme_cceip2_ob_out.tdata [37]);
tran (kme_cceip2_ob_out[36], \kme_cceip2_ob_out.tdata [36]);
tran (kme_cceip2_ob_out[35], \kme_cceip2_ob_out.tdata [35]);
tran (kme_cceip2_ob_out[34], \kme_cceip2_ob_out.tdata [34]);
tran (kme_cceip2_ob_out[33], \kme_cceip2_ob_out.tdata [33]);
tran (kme_cceip2_ob_out[32], \kme_cceip2_ob_out.tdata [32]);
tran (kme_cceip2_ob_out[31], \kme_cceip2_ob_out.tdata [31]);
tran (kme_cceip2_ob_out[30], \kme_cceip2_ob_out.tdata [30]);
tran (kme_cceip2_ob_out[29], \kme_cceip2_ob_out.tdata [29]);
tran (kme_cceip2_ob_out[28], \kme_cceip2_ob_out.tdata [28]);
tran (kme_cceip2_ob_out[27], \kme_cceip2_ob_out.tdata [27]);
tran (kme_cceip2_ob_out[26], \kme_cceip2_ob_out.tdata [26]);
tran (kme_cceip2_ob_out[25], \kme_cceip2_ob_out.tdata [25]);
tran (kme_cceip2_ob_out[24], \kme_cceip2_ob_out.tdata [24]);
tran (kme_cceip2_ob_out[23], \kme_cceip2_ob_out.tdata [23]);
tran (kme_cceip2_ob_out[22], \kme_cceip2_ob_out.tdata [22]);
tran (kme_cceip2_ob_out[21], \kme_cceip2_ob_out.tdata [21]);
tran (kme_cceip2_ob_out[20], \kme_cceip2_ob_out.tdata [20]);
tran (kme_cceip2_ob_out[19], \kme_cceip2_ob_out.tdata [19]);
tran (kme_cceip2_ob_out[18], \kme_cceip2_ob_out.tdata [18]);
tran (kme_cceip2_ob_out[17], \kme_cceip2_ob_out.tdata [17]);
tran (kme_cceip2_ob_out[16], \kme_cceip2_ob_out.tdata [16]);
tran (kme_cceip2_ob_out[15], \kme_cceip2_ob_out.tdata [15]);
tran (kme_cceip2_ob_out[14], \kme_cceip2_ob_out.tdata [14]);
tran (kme_cceip2_ob_out[13], \kme_cceip2_ob_out.tdata [13]);
tran (kme_cceip2_ob_out[12], \kme_cceip2_ob_out.tdata [12]);
tran (kme_cceip2_ob_out[11], \kme_cceip2_ob_out.tdata [11]);
tran (kme_cceip2_ob_out[10], \kme_cceip2_ob_out.tdata [10]);
tran (kme_cceip2_ob_out[9], \kme_cceip2_ob_out.tdata [9]);
tran (kme_cceip2_ob_out[8], \kme_cceip2_ob_out.tdata [8]);
tran (kme_cceip2_ob_out[7], \kme_cceip2_ob_out.tdata [7]);
tran (kme_cceip2_ob_out[6], \kme_cceip2_ob_out.tdata [6]);
tran (kme_cceip2_ob_out[5], \kme_cceip2_ob_out.tdata [5]);
tran (kme_cceip2_ob_out[4], \kme_cceip2_ob_out.tdata [4]);
tran (kme_cceip2_ob_out[3], \kme_cceip2_ob_out.tdata [3]);
tran (kme_cceip2_ob_out[2], \kme_cceip2_ob_out.tdata [2]);
tran (kme_cceip2_ob_out[1], \kme_cceip2_ob_out.tdata [1]);
tran (kme_cceip2_ob_out[0], \kme_cceip2_ob_out.tdata [0]);
tran (kme_cceip2_ob_in_mod[0], \kme_cceip2_ob_in_mod.tready );
tran (kme_cceip3_ob_out[82], \kme_cceip3_ob_out.tvalid );
tran (kme_cceip3_ob_out[81], \kme_cceip3_ob_out.tlast );
tran (kme_cceip3_ob_out[80], \kme_cceip3_ob_out.tid [0]);
tran (kme_cceip3_ob_out[79], \kme_cceip3_ob_out.tstrb [7]);
tran (kme_cceip3_ob_out[78], \kme_cceip3_ob_out.tstrb [6]);
tran (kme_cceip3_ob_out[77], \kme_cceip3_ob_out.tstrb [5]);
tran (kme_cceip3_ob_out[76], \kme_cceip3_ob_out.tstrb [4]);
tran (kme_cceip3_ob_out[75], \kme_cceip3_ob_out.tstrb [3]);
tran (kme_cceip3_ob_out[74], \kme_cceip3_ob_out.tstrb [2]);
tran (kme_cceip3_ob_out[73], \kme_cceip3_ob_out.tstrb [1]);
tran (kme_cceip3_ob_out[72], \kme_cceip3_ob_out.tstrb [0]);
tran (kme_cceip3_ob_out[71], \kme_cceip3_ob_out.tuser [7]);
tran (kme_cceip3_ob_out[70], \kme_cceip3_ob_out.tuser [6]);
tran (kme_cceip3_ob_out[69], \kme_cceip3_ob_out.tuser [5]);
tran (kme_cceip3_ob_out[68], \kme_cceip3_ob_out.tuser [4]);
tran (kme_cceip3_ob_out[67], \kme_cceip3_ob_out.tuser [3]);
tran (kme_cceip3_ob_out[66], \kme_cceip3_ob_out.tuser [2]);
tran (kme_cceip3_ob_out[65], \kme_cceip3_ob_out.tuser [1]);
tran (kme_cceip3_ob_out[64], \kme_cceip3_ob_out.tuser [0]);
tran (kme_cceip3_ob_out[63], \kme_cceip3_ob_out.tdata [63]);
tran (kme_cceip3_ob_out[62], \kme_cceip3_ob_out.tdata [62]);
tran (kme_cceip3_ob_out[61], \kme_cceip3_ob_out.tdata [61]);
tran (kme_cceip3_ob_out[60], \kme_cceip3_ob_out.tdata [60]);
tran (kme_cceip3_ob_out[59], \kme_cceip3_ob_out.tdata [59]);
tran (kme_cceip3_ob_out[58], \kme_cceip3_ob_out.tdata [58]);
tran (kme_cceip3_ob_out[57], \kme_cceip3_ob_out.tdata [57]);
tran (kme_cceip3_ob_out[56], \kme_cceip3_ob_out.tdata [56]);
tran (kme_cceip3_ob_out[55], \kme_cceip3_ob_out.tdata [55]);
tran (kme_cceip3_ob_out[54], \kme_cceip3_ob_out.tdata [54]);
tran (kme_cceip3_ob_out[53], \kme_cceip3_ob_out.tdata [53]);
tran (kme_cceip3_ob_out[52], \kme_cceip3_ob_out.tdata [52]);
tran (kme_cceip3_ob_out[51], \kme_cceip3_ob_out.tdata [51]);
tran (kme_cceip3_ob_out[50], \kme_cceip3_ob_out.tdata [50]);
tran (kme_cceip3_ob_out[49], \kme_cceip3_ob_out.tdata [49]);
tran (kme_cceip3_ob_out[48], \kme_cceip3_ob_out.tdata [48]);
tran (kme_cceip3_ob_out[47], \kme_cceip3_ob_out.tdata [47]);
tran (kme_cceip3_ob_out[46], \kme_cceip3_ob_out.tdata [46]);
tran (kme_cceip3_ob_out[45], \kme_cceip3_ob_out.tdata [45]);
tran (kme_cceip3_ob_out[44], \kme_cceip3_ob_out.tdata [44]);
tran (kme_cceip3_ob_out[43], \kme_cceip3_ob_out.tdata [43]);
tran (kme_cceip3_ob_out[42], \kme_cceip3_ob_out.tdata [42]);
tran (kme_cceip3_ob_out[41], \kme_cceip3_ob_out.tdata [41]);
tran (kme_cceip3_ob_out[40], \kme_cceip3_ob_out.tdata [40]);
tran (kme_cceip3_ob_out[39], \kme_cceip3_ob_out.tdata [39]);
tran (kme_cceip3_ob_out[38], \kme_cceip3_ob_out.tdata [38]);
tran (kme_cceip3_ob_out[37], \kme_cceip3_ob_out.tdata [37]);
tran (kme_cceip3_ob_out[36], \kme_cceip3_ob_out.tdata [36]);
tran (kme_cceip3_ob_out[35], \kme_cceip3_ob_out.tdata [35]);
tran (kme_cceip3_ob_out[34], \kme_cceip3_ob_out.tdata [34]);
tran (kme_cceip3_ob_out[33], \kme_cceip3_ob_out.tdata [33]);
tran (kme_cceip3_ob_out[32], \kme_cceip3_ob_out.tdata [32]);
tran (kme_cceip3_ob_out[31], \kme_cceip3_ob_out.tdata [31]);
tran (kme_cceip3_ob_out[30], \kme_cceip3_ob_out.tdata [30]);
tran (kme_cceip3_ob_out[29], \kme_cceip3_ob_out.tdata [29]);
tran (kme_cceip3_ob_out[28], \kme_cceip3_ob_out.tdata [28]);
tran (kme_cceip3_ob_out[27], \kme_cceip3_ob_out.tdata [27]);
tran (kme_cceip3_ob_out[26], \kme_cceip3_ob_out.tdata [26]);
tran (kme_cceip3_ob_out[25], \kme_cceip3_ob_out.tdata [25]);
tran (kme_cceip3_ob_out[24], \kme_cceip3_ob_out.tdata [24]);
tran (kme_cceip3_ob_out[23], \kme_cceip3_ob_out.tdata [23]);
tran (kme_cceip3_ob_out[22], \kme_cceip3_ob_out.tdata [22]);
tran (kme_cceip3_ob_out[21], \kme_cceip3_ob_out.tdata [21]);
tran (kme_cceip3_ob_out[20], \kme_cceip3_ob_out.tdata [20]);
tran (kme_cceip3_ob_out[19], \kme_cceip3_ob_out.tdata [19]);
tran (kme_cceip3_ob_out[18], \kme_cceip3_ob_out.tdata [18]);
tran (kme_cceip3_ob_out[17], \kme_cceip3_ob_out.tdata [17]);
tran (kme_cceip3_ob_out[16], \kme_cceip3_ob_out.tdata [16]);
tran (kme_cceip3_ob_out[15], \kme_cceip3_ob_out.tdata [15]);
tran (kme_cceip3_ob_out[14], \kme_cceip3_ob_out.tdata [14]);
tran (kme_cceip3_ob_out[13], \kme_cceip3_ob_out.tdata [13]);
tran (kme_cceip3_ob_out[12], \kme_cceip3_ob_out.tdata [12]);
tran (kme_cceip3_ob_out[11], \kme_cceip3_ob_out.tdata [11]);
tran (kme_cceip3_ob_out[10], \kme_cceip3_ob_out.tdata [10]);
tran (kme_cceip3_ob_out[9], \kme_cceip3_ob_out.tdata [9]);
tran (kme_cceip3_ob_out[8], \kme_cceip3_ob_out.tdata [8]);
tran (kme_cceip3_ob_out[7], \kme_cceip3_ob_out.tdata [7]);
tran (kme_cceip3_ob_out[6], \kme_cceip3_ob_out.tdata [6]);
tran (kme_cceip3_ob_out[5], \kme_cceip3_ob_out.tdata [5]);
tran (kme_cceip3_ob_out[4], \kme_cceip3_ob_out.tdata [4]);
tran (kme_cceip3_ob_out[3], \kme_cceip3_ob_out.tdata [3]);
tran (kme_cceip3_ob_out[2], \kme_cceip3_ob_out.tdata [2]);
tran (kme_cceip3_ob_out[1], \kme_cceip3_ob_out.tdata [1]);
tran (kme_cceip3_ob_out[0], \kme_cceip3_ob_out.tdata [0]);
tran (kme_cceip3_ob_in_mod[0], \kme_cceip3_ob_in_mod.tready );
tran (kme_cddip0_ob_out[82], \kme_cddip0_ob_out.tvalid );
tran (kme_cddip0_ob_out[81], \kme_cddip0_ob_out.tlast );
tran (kme_cddip0_ob_out[80], \kme_cddip0_ob_out.tid [0]);
tran (kme_cddip0_ob_out[79], \kme_cddip0_ob_out.tstrb [7]);
tran (kme_cddip0_ob_out[78], \kme_cddip0_ob_out.tstrb [6]);
tran (kme_cddip0_ob_out[77], \kme_cddip0_ob_out.tstrb [5]);
tran (kme_cddip0_ob_out[76], \kme_cddip0_ob_out.tstrb [4]);
tran (kme_cddip0_ob_out[75], \kme_cddip0_ob_out.tstrb [3]);
tran (kme_cddip0_ob_out[74], \kme_cddip0_ob_out.tstrb [2]);
tran (kme_cddip0_ob_out[73], \kme_cddip0_ob_out.tstrb [1]);
tran (kme_cddip0_ob_out[72], \kme_cddip0_ob_out.tstrb [0]);
tran (kme_cddip0_ob_out[71], \kme_cddip0_ob_out.tuser [7]);
tran (kme_cddip0_ob_out[70], \kme_cddip0_ob_out.tuser [6]);
tran (kme_cddip0_ob_out[69], \kme_cddip0_ob_out.tuser [5]);
tran (kme_cddip0_ob_out[68], \kme_cddip0_ob_out.tuser [4]);
tran (kme_cddip0_ob_out[67], \kme_cddip0_ob_out.tuser [3]);
tran (kme_cddip0_ob_out[66], \kme_cddip0_ob_out.tuser [2]);
tran (kme_cddip0_ob_out[65], \kme_cddip0_ob_out.tuser [1]);
tran (kme_cddip0_ob_out[64], \kme_cddip0_ob_out.tuser [0]);
tran (kme_cddip0_ob_out[63], \kme_cddip0_ob_out.tdata [63]);
tran (kme_cddip0_ob_out[62], \kme_cddip0_ob_out.tdata [62]);
tran (kme_cddip0_ob_out[61], \kme_cddip0_ob_out.tdata [61]);
tran (kme_cddip0_ob_out[60], \kme_cddip0_ob_out.tdata [60]);
tran (kme_cddip0_ob_out[59], \kme_cddip0_ob_out.tdata [59]);
tran (kme_cddip0_ob_out[58], \kme_cddip0_ob_out.tdata [58]);
tran (kme_cddip0_ob_out[57], \kme_cddip0_ob_out.tdata [57]);
tran (kme_cddip0_ob_out[56], \kme_cddip0_ob_out.tdata [56]);
tran (kme_cddip0_ob_out[55], \kme_cddip0_ob_out.tdata [55]);
tran (kme_cddip0_ob_out[54], \kme_cddip0_ob_out.tdata [54]);
tran (kme_cddip0_ob_out[53], \kme_cddip0_ob_out.tdata [53]);
tran (kme_cddip0_ob_out[52], \kme_cddip0_ob_out.tdata [52]);
tran (kme_cddip0_ob_out[51], \kme_cddip0_ob_out.tdata [51]);
tran (kme_cddip0_ob_out[50], \kme_cddip0_ob_out.tdata [50]);
tran (kme_cddip0_ob_out[49], \kme_cddip0_ob_out.tdata [49]);
tran (kme_cddip0_ob_out[48], \kme_cddip0_ob_out.tdata [48]);
tran (kme_cddip0_ob_out[47], \kme_cddip0_ob_out.tdata [47]);
tran (kme_cddip0_ob_out[46], \kme_cddip0_ob_out.tdata [46]);
tran (kme_cddip0_ob_out[45], \kme_cddip0_ob_out.tdata [45]);
tran (kme_cddip0_ob_out[44], \kme_cddip0_ob_out.tdata [44]);
tran (kme_cddip0_ob_out[43], \kme_cddip0_ob_out.tdata [43]);
tran (kme_cddip0_ob_out[42], \kme_cddip0_ob_out.tdata [42]);
tran (kme_cddip0_ob_out[41], \kme_cddip0_ob_out.tdata [41]);
tran (kme_cddip0_ob_out[40], \kme_cddip0_ob_out.tdata [40]);
tran (kme_cddip0_ob_out[39], \kme_cddip0_ob_out.tdata [39]);
tran (kme_cddip0_ob_out[38], \kme_cddip0_ob_out.tdata [38]);
tran (kme_cddip0_ob_out[37], \kme_cddip0_ob_out.tdata [37]);
tran (kme_cddip0_ob_out[36], \kme_cddip0_ob_out.tdata [36]);
tran (kme_cddip0_ob_out[35], \kme_cddip0_ob_out.tdata [35]);
tran (kme_cddip0_ob_out[34], \kme_cddip0_ob_out.tdata [34]);
tran (kme_cddip0_ob_out[33], \kme_cddip0_ob_out.tdata [33]);
tran (kme_cddip0_ob_out[32], \kme_cddip0_ob_out.tdata [32]);
tran (kme_cddip0_ob_out[31], \kme_cddip0_ob_out.tdata [31]);
tran (kme_cddip0_ob_out[30], \kme_cddip0_ob_out.tdata [30]);
tran (kme_cddip0_ob_out[29], \kme_cddip0_ob_out.tdata [29]);
tran (kme_cddip0_ob_out[28], \kme_cddip0_ob_out.tdata [28]);
tran (kme_cddip0_ob_out[27], \kme_cddip0_ob_out.tdata [27]);
tran (kme_cddip0_ob_out[26], \kme_cddip0_ob_out.tdata [26]);
tran (kme_cddip0_ob_out[25], \kme_cddip0_ob_out.tdata [25]);
tran (kme_cddip0_ob_out[24], \kme_cddip0_ob_out.tdata [24]);
tran (kme_cddip0_ob_out[23], \kme_cddip0_ob_out.tdata [23]);
tran (kme_cddip0_ob_out[22], \kme_cddip0_ob_out.tdata [22]);
tran (kme_cddip0_ob_out[21], \kme_cddip0_ob_out.tdata [21]);
tran (kme_cddip0_ob_out[20], \kme_cddip0_ob_out.tdata [20]);
tran (kme_cddip0_ob_out[19], \kme_cddip0_ob_out.tdata [19]);
tran (kme_cddip0_ob_out[18], \kme_cddip0_ob_out.tdata [18]);
tran (kme_cddip0_ob_out[17], \kme_cddip0_ob_out.tdata [17]);
tran (kme_cddip0_ob_out[16], \kme_cddip0_ob_out.tdata [16]);
tran (kme_cddip0_ob_out[15], \kme_cddip0_ob_out.tdata [15]);
tran (kme_cddip0_ob_out[14], \kme_cddip0_ob_out.tdata [14]);
tran (kme_cddip0_ob_out[13], \kme_cddip0_ob_out.tdata [13]);
tran (kme_cddip0_ob_out[12], \kme_cddip0_ob_out.tdata [12]);
tran (kme_cddip0_ob_out[11], \kme_cddip0_ob_out.tdata [11]);
tran (kme_cddip0_ob_out[10], \kme_cddip0_ob_out.tdata [10]);
tran (kme_cddip0_ob_out[9], \kme_cddip0_ob_out.tdata [9]);
tran (kme_cddip0_ob_out[8], \kme_cddip0_ob_out.tdata [8]);
tran (kme_cddip0_ob_out[7], \kme_cddip0_ob_out.tdata [7]);
tran (kme_cddip0_ob_out[6], \kme_cddip0_ob_out.tdata [6]);
tran (kme_cddip0_ob_out[5], \kme_cddip0_ob_out.tdata [5]);
tran (kme_cddip0_ob_out[4], \kme_cddip0_ob_out.tdata [4]);
tran (kme_cddip0_ob_out[3], \kme_cddip0_ob_out.tdata [3]);
tran (kme_cddip0_ob_out[2], \kme_cddip0_ob_out.tdata [2]);
tran (kme_cddip0_ob_out[1], \kme_cddip0_ob_out.tdata [1]);
tran (kme_cddip0_ob_out[0], \kme_cddip0_ob_out.tdata [0]);
tran (kme_cddip0_ob_in_mod[0], \kme_cddip0_ob_in_mod.tready );
tran (kme_cddip1_ob_out[82], \kme_cddip1_ob_out.tvalid );
tran (kme_cddip1_ob_out[81], \kme_cddip1_ob_out.tlast );
tran (kme_cddip1_ob_out[80], \kme_cddip1_ob_out.tid [0]);
tran (kme_cddip1_ob_out[79], \kme_cddip1_ob_out.tstrb [7]);
tran (kme_cddip1_ob_out[78], \kme_cddip1_ob_out.tstrb [6]);
tran (kme_cddip1_ob_out[77], \kme_cddip1_ob_out.tstrb [5]);
tran (kme_cddip1_ob_out[76], \kme_cddip1_ob_out.tstrb [4]);
tran (kme_cddip1_ob_out[75], \kme_cddip1_ob_out.tstrb [3]);
tran (kme_cddip1_ob_out[74], \kme_cddip1_ob_out.tstrb [2]);
tran (kme_cddip1_ob_out[73], \kme_cddip1_ob_out.tstrb [1]);
tran (kme_cddip1_ob_out[72], \kme_cddip1_ob_out.tstrb [0]);
tran (kme_cddip1_ob_out[71], \kme_cddip1_ob_out.tuser [7]);
tran (kme_cddip1_ob_out[70], \kme_cddip1_ob_out.tuser [6]);
tran (kme_cddip1_ob_out[69], \kme_cddip1_ob_out.tuser [5]);
tran (kme_cddip1_ob_out[68], \kme_cddip1_ob_out.tuser [4]);
tran (kme_cddip1_ob_out[67], \kme_cddip1_ob_out.tuser [3]);
tran (kme_cddip1_ob_out[66], \kme_cddip1_ob_out.tuser [2]);
tran (kme_cddip1_ob_out[65], \kme_cddip1_ob_out.tuser [1]);
tran (kme_cddip1_ob_out[64], \kme_cddip1_ob_out.tuser [0]);
tran (kme_cddip1_ob_out[63], \kme_cddip1_ob_out.tdata [63]);
tran (kme_cddip1_ob_out[62], \kme_cddip1_ob_out.tdata [62]);
tran (kme_cddip1_ob_out[61], \kme_cddip1_ob_out.tdata [61]);
tran (kme_cddip1_ob_out[60], \kme_cddip1_ob_out.tdata [60]);
tran (kme_cddip1_ob_out[59], \kme_cddip1_ob_out.tdata [59]);
tran (kme_cddip1_ob_out[58], \kme_cddip1_ob_out.tdata [58]);
tran (kme_cddip1_ob_out[57], \kme_cddip1_ob_out.tdata [57]);
tran (kme_cddip1_ob_out[56], \kme_cddip1_ob_out.tdata [56]);
tran (kme_cddip1_ob_out[55], \kme_cddip1_ob_out.tdata [55]);
tran (kme_cddip1_ob_out[54], \kme_cddip1_ob_out.tdata [54]);
tran (kme_cddip1_ob_out[53], \kme_cddip1_ob_out.tdata [53]);
tran (kme_cddip1_ob_out[52], \kme_cddip1_ob_out.tdata [52]);
tran (kme_cddip1_ob_out[51], \kme_cddip1_ob_out.tdata [51]);
tran (kme_cddip1_ob_out[50], \kme_cddip1_ob_out.tdata [50]);
tran (kme_cddip1_ob_out[49], \kme_cddip1_ob_out.tdata [49]);
tran (kme_cddip1_ob_out[48], \kme_cddip1_ob_out.tdata [48]);
tran (kme_cddip1_ob_out[47], \kme_cddip1_ob_out.tdata [47]);
tran (kme_cddip1_ob_out[46], \kme_cddip1_ob_out.tdata [46]);
tran (kme_cddip1_ob_out[45], \kme_cddip1_ob_out.tdata [45]);
tran (kme_cddip1_ob_out[44], \kme_cddip1_ob_out.tdata [44]);
tran (kme_cddip1_ob_out[43], \kme_cddip1_ob_out.tdata [43]);
tran (kme_cddip1_ob_out[42], \kme_cddip1_ob_out.tdata [42]);
tran (kme_cddip1_ob_out[41], \kme_cddip1_ob_out.tdata [41]);
tran (kme_cddip1_ob_out[40], \kme_cddip1_ob_out.tdata [40]);
tran (kme_cddip1_ob_out[39], \kme_cddip1_ob_out.tdata [39]);
tran (kme_cddip1_ob_out[38], \kme_cddip1_ob_out.tdata [38]);
tran (kme_cddip1_ob_out[37], \kme_cddip1_ob_out.tdata [37]);
tran (kme_cddip1_ob_out[36], \kme_cddip1_ob_out.tdata [36]);
tran (kme_cddip1_ob_out[35], \kme_cddip1_ob_out.tdata [35]);
tran (kme_cddip1_ob_out[34], \kme_cddip1_ob_out.tdata [34]);
tran (kme_cddip1_ob_out[33], \kme_cddip1_ob_out.tdata [33]);
tran (kme_cddip1_ob_out[32], \kme_cddip1_ob_out.tdata [32]);
tran (kme_cddip1_ob_out[31], \kme_cddip1_ob_out.tdata [31]);
tran (kme_cddip1_ob_out[30], \kme_cddip1_ob_out.tdata [30]);
tran (kme_cddip1_ob_out[29], \kme_cddip1_ob_out.tdata [29]);
tran (kme_cddip1_ob_out[28], \kme_cddip1_ob_out.tdata [28]);
tran (kme_cddip1_ob_out[27], \kme_cddip1_ob_out.tdata [27]);
tran (kme_cddip1_ob_out[26], \kme_cddip1_ob_out.tdata [26]);
tran (kme_cddip1_ob_out[25], \kme_cddip1_ob_out.tdata [25]);
tran (kme_cddip1_ob_out[24], \kme_cddip1_ob_out.tdata [24]);
tran (kme_cddip1_ob_out[23], \kme_cddip1_ob_out.tdata [23]);
tran (kme_cddip1_ob_out[22], \kme_cddip1_ob_out.tdata [22]);
tran (kme_cddip1_ob_out[21], \kme_cddip1_ob_out.tdata [21]);
tran (kme_cddip1_ob_out[20], \kme_cddip1_ob_out.tdata [20]);
tran (kme_cddip1_ob_out[19], \kme_cddip1_ob_out.tdata [19]);
tran (kme_cddip1_ob_out[18], \kme_cddip1_ob_out.tdata [18]);
tran (kme_cddip1_ob_out[17], \kme_cddip1_ob_out.tdata [17]);
tran (kme_cddip1_ob_out[16], \kme_cddip1_ob_out.tdata [16]);
tran (kme_cddip1_ob_out[15], \kme_cddip1_ob_out.tdata [15]);
tran (kme_cddip1_ob_out[14], \kme_cddip1_ob_out.tdata [14]);
tran (kme_cddip1_ob_out[13], \kme_cddip1_ob_out.tdata [13]);
tran (kme_cddip1_ob_out[12], \kme_cddip1_ob_out.tdata [12]);
tran (kme_cddip1_ob_out[11], \kme_cddip1_ob_out.tdata [11]);
tran (kme_cddip1_ob_out[10], \kme_cddip1_ob_out.tdata [10]);
tran (kme_cddip1_ob_out[9], \kme_cddip1_ob_out.tdata [9]);
tran (kme_cddip1_ob_out[8], \kme_cddip1_ob_out.tdata [8]);
tran (kme_cddip1_ob_out[7], \kme_cddip1_ob_out.tdata [7]);
tran (kme_cddip1_ob_out[6], \kme_cddip1_ob_out.tdata [6]);
tran (kme_cddip1_ob_out[5], \kme_cddip1_ob_out.tdata [5]);
tran (kme_cddip1_ob_out[4], \kme_cddip1_ob_out.tdata [4]);
tran (kme_cddip1_ob_out[3], \kme_cddip1_ob_out.tdata [3]);
tran (kme_cddip1_ob_out[2], \kme_cddip1_ob_out.tdata [2]);
tran (kme_cddip1_ob_out[1], \kme_cddip1_ob_out.tdata [1]);
tran (kme_cddip1_ob_out[0], \kme_cddip1_ob_out.tdata [0]);
tran (kme_cddip1_ob_in_mod[0], \kme_cddip1_ob_in_mod.tready );
tran (kme_cddip2_ob_out[82], \kme_cddip2_ob_out.tvalid );
tran (kme_cddip2_ob_out[81], \kme_cddip2_ob_out.tlast );
tran (kme_cddip2_ob_out[80], \kme_cddip2_ob_out.tid [0]);
tran (kme_cddip2_ob_out[79], \kme_cddip2_ob_out.tstrb [7]);
tran (kme_cddip2_ob_out[78], \kme_cddip2_ob_out.tstrb [6]);
tran (kme_cddip2_ob_out[77], \kme_cddip2_ob_out.tstrb [5]);
tran (kme_cddip2_ob_out[76], \kme_cddip2_ob_out.tstrb [4]);
tran (kme_cddip2_ob_out[75], \kme_cddip2_ob_out.tstrb [3]);
tran (kme_cddip2_ob_out[74], \kme_cddip2_ob_out.tstrb [2]);
tran (kme_cddip2_ob_out[73], \kme_cddip2_ob_out.tstrb [1]);
tran (kme_cddip2_ob_out[72], \kme_cddip2_ob_out.tstrb [0]);
tran (kme_cddip2_ob_out[71], \kme_cddip2_ob_out.tuser [7]);
tran (kme_cddip2_ob_out[70], \kme_cddip2_ob_out.tuser [6]);
tran (kme_cddip2_ob_out[69], \kme_cddip2_ob_out.tuser [5]);
tran (kme_cddip2_ob_out[68], \kme_cddip2_ob_out.tuser [4]);
tran (kme_cddip2_ob_out[67], \kme_cddip2_ob_out.tuser [3]);
tran (kme_cddip2_ob_out[66], \kme_cddip2_ob_out.tuser [2]);
tran (kme_cddip2_ob_out[65], \kme_cddip2_ob_out.tuser [1]);
tran (kme_cddip2_ob_out[64], \kme_cddip2_ob_out.tuser [0]);
tran (kme_cddip2_ob_out[63], \kme_cddip2_ob_out.tdata [63]);
tran (kme_cddip2_ob_out[62], \kme_cddip2_ob_out.tdata [62]);
tran (kme_cddip2_ob_out[61], \kme_cddip2_ob_out.tdata [61]);
tran (kme_cddip2_ob_out[60], \kme_cddip2_ob_out.tdata [60]);
tran (kme_cddip2_ob_out[59], \kme_cddip2_ob_out.tdata [59]);
tran (kme_cddip2_ob_out[58], \kme_cddip2_ob_out.tdata [58]);
tran (kme_cddip2_ob_out[57], \kme_cddip2_ob_out.tdata [57]);
tran (kme_cddip2_ob_out[56], \kme_cddip2_ob_out.tdata [56]);
tran (kme_cddip2_ob_out[55], \kme_cddip2_ob_out.tdata [55]);
tran (kme_cddip2_ob_out[54], \kme_cddip2_ob_out.tdata [54]);
tran (kme_cddip2_ob_out[53], \kme_cddip2_ob_out.tdata [53]);
tran (kme_cddip2_ob_out[52], \kme_cddip2_ob_out.tdata [52]);
tran (kme_cddip2_ob_out[51], \kme_cddip2_ob_out.tdata [51]);
tran (kme_cddip2_ob_out[50], \kme_cddip2_ob_out.tdata [50]);
tran (kme_cddip2_ob_out[49], \kme_cddip2_ob_out.tdata [49]);
tran (kme_cddip2_ob_out[48], \kme_cddip2_ob_out.tdata [48]);
tran (kme_cddip2_ob_out[47], \kme_cddip2_ob_out.tdata [47]);
tran (kme_cddip2_ob_out[46], \kme_cddip2_ob_out.tdata [46]);
tran (kme_cddip2_ob_out[45], \kme_cddip2_ob_out.tdata [45]);
tran (kme_cddip2_ob_out[44], \kme_cddip2_ob_out.tdata [44]);
tran (kme_cddip2_ob_out[43], \kme_cddip2_ob_out.tdata [43]);
tran (kme_cddip2_ob_out[42], \kme_cddip2_ob_out.tdata [42]);
tran (kme_cddip2_ob_out[41], \kme_cddip2_ob_out.tdata [41]);
tran (kme_cddip2_ob_out[40], \kme_cddip2_ob_out.tdata [40]);
tran (kme_cddip2_ob_out[39], \kme_cddip2_ob_out.tdata [39]);
tran (kme_cddip2_ob_out[38], \kme_cddip2_ob_out.tdata [38]);
tran (kme_cddip2_ob_out[37], \kme_cddip2_ob_out.tdata [37]);
tran (kme_cddip2_ob_out[36], \kme_cddip2_ob_out.tdata [36]);
tran (kme_cddip2_ob_out[35], \kme_cddip2_ob_out.tdata [35]);
tran (kme_cddip2_ob_out[34], \kme_cddip2_ob_out.tdata [34]);
tran (kme_cddip2_ob_out[33], \kme_cddip2_ob_out.tdata [33]);
tran (kme_cddip2_ob_out[32], \kme_cddip2_ob_out.tdata [32]);
tran (kme_cddip2_ob_out[31], \kme_cddip2_ob_out.tdata [31]);
tran (kme_cddip2_ob_out[30], \kme_cddip2_ob_out.tdata [30]);
tran (kme_cddip2_ob_out[29], \kme_cddip2_ob_out.tdata [29]);
tran (kme_cddip2_ob_out[28], \kme_cddip2_ob_out.tdata [28]);
tran (kme_cddip2_ob_out[27], \kme_cddip2_ob_out.tdata [27]);
tran (kme_cddip2_ob_out[26], \kme_cddip2_ob_out.tdata [26]);
tran (kme_cddip2_ob_out[25], \kme_cddip2_ob_out.tdata [25]);
tran (kme_cddip2_ob_out[24], \kme_cddip2_ob_out.tdata [24]);
tran (kme_cddip2_ob_out[23], \kme_cddip2_ob_out.tdata [23]);
tran (kme_cddip2_ob_out[22], \kme_cddip2_ob_out.tdata [22]);
tran (kme_cddip2_ob_out[21], \kme_cddip2_ob_out.tdata [21]);
tran (kme_cddip2_ob_out[20], \kme_cddip2_ob_out.tdata [20]);
tran (kme_cddip2_ob_out[19], \kme_cddip2_ob_out.tdata [19]);
tran (kme_cddip2_ob_out[18], \kme_cddip2_ob_out.tdata [18]);
tran (kme_cddip2_ob_out[17], \kme_cddip2_ob_out.tdata [17]);
tran (kme_cddip2_ob_out[16], \kme_cddip2_ob_out.tdata [16]);
tran (kme_cddip2_ob_out[15], \kme_cddip2_ob_out.tdata [15]);
tran (kme_cddip2_ob_out[14], \kme_cddip2_ob_out.tdata [14]);
tran (kme_cddip2_ob_out[13], \kme_cddip2_ob_out.tdata [13]);
tran (kme_cddip2_ob_out[12], \kme_cddip2_ob_out.tdata [12]);
tran (kme_cddip2_ob_out[11], \kme_cddip2_ob_out.tdata [11]);
tran (kme_cddip2_ob_out[10], \kme_cddip2_ob_out.tdata [10]);
tran (kme_cddip2_ob_out[9], \kme_cddip2_ob_out.tdata [9]);
tran (kme_cddip2_ob_out[8], \kme_cddip2_ob_out.tdata [8]);
tran (kme_cddip2_ob_out[7], \kme_cddip2_ob_out.tdata [7]);
tran (kme_cddip2_ob_out[6], \kme_cddip2_ob_out.tdata [6]);
tran (kme_cddip2_ob_out[5], \kme_cddip2_ob_out.tdata [5]);
tran (kme_cddip2_ob_out[4], \kme_cddip2_ob_out.tdata [4]);
tran (kme_cddip2_ob_out[3], \kme_cddip2_ob_out.tdata [3]);
tran (kme_cddip2_ob_out[2], \kme_cddip2_ob_out.tdata [2]);
tran (kme_cddip2_ob_out[1], \kme_cddip2_ob_out.tdata [1]);
tran (kme_cddip2_ob_out[0], \kme_cddip2_ob_out.tdata [0]);
tran (kme_cddip2_ob_in_mod[0], \kme_cddip2_ob_in_mod.tready );
tran (kme_cddip3_ob_out[82], \kme_cddip3_ob_out.tvalid );
tran (kme_cddip3_ob_out[81], \kme_cddip3_ob_out.tlast );
tran (kme_cddip3_ob_out[80], \kme_cddip3_ob_out.tid [0]);
tran (kme_cddip3_ob_out[79], \kme_cddip3_ob_out.tstrb [7]);
tran (kme_cddip3_ob_out[78], \kme_cddip3_ob_out.tstrb [6]);
tran (kme_cddip3_ob_out[77], \kme_cddip3_ob_out.tstrb [5]);
tran (kme_cddip3_ob_out[76], \kme_cddip3_ob_out.tstrb [4]);
tran (kme_cddip3_ob_out[75], \kme_cddip3_ob_out.tstrb [3]);
tran (kme_cddip3_ob_out[74], \kme_cddip3_ob_out.tstrb [2]);
tran (kme_cddip3_ob_out[73], \kme_cddip3_ob_out.tstrb [1]);
tran (kme_cddip3_ob_out[72], \kme_cddip3_ob_out.tstrb [0]);
tran (kme_cddip3_ob_out[71], \kme_cddip3_ob_out.tuser [7]);
tran (kme_cddip3_ob_out[70], \kme_cddip3_ob_out.tuser [6]);
tran (kme_cddip3_ob_out[69], \kme_cddip3_ob_out.tuser [5]);
tran (kme_cddip3_ob_out[68], \kme_cddip3_ob_out.tuser [4]);
tran (kme_cddip3_ob_out[67], \kme_cddip3_ob_out.tuser [3]);
tran (kme_cddip3_ob_out[66], \kme_cddip3_ob_out.tuser [2]);
tran (kme_cddip3_ob_out[65], \kme_cddip3_ob_out.tuser [1]);
tran (kme_cddip3_ob_out[64], \kme_cddip3_ob_out.tuser [0]);
tran (kme_cddip3_ob_out[63], \kme_cddip3_ob_out.tdata [63]);
tran (kme_cddip3_ob_out[62], \kme_cddip3_ob_out.tdata [62]);
tran (kme_cddip3_ob_out[61], \kme_cddip3_ob_out.tdata [61]);
tran (kme_cddip3_ob_out[60], \kme_cddip3_ob_out.tdata [60]);
tran (kme_cddip3_ob_out[59], \kme_cddip3_ob_out.tdata [59]);
tran (kme_cddip3_ob_out[58], \kme_cddip3_ob_out.tdata [58]);
tran (kme_cddip3_ob_out[57], \kme_cddip3_ob_out.tdata [57]);
tran (kme_cddip3_ob_out[56], \kme_cddip3_ob_out.tdata [56]);
tran (kme_cddip3_ob_out[55], \kme_cddip3_ob_out.tdata [55]);
tran (kme_cddip3_ob_out[54], \kme_cddip3_ob_out.tdata [54]);
tran (kme_cddip3_ob_out[53], \kme_cddip3_ob_out.tdata [53]);
tran (kme_cddip3_ob_out[52], \kme_cddip3_ob_out.tdata [52]);
tran (kme_cddip3_ob_out[51], \kme_cddip3_ob_out.tdata [51]);
tran (kme_cddip3_ob_out[50], \kme_cddip3_ob_out.tdata [50]);
tran (kme_cddip3_ob_out[49], \kme_cddip3_ob_out.tdata [49]);
tran (kme_cddip3_ob_out[48], \kme_cddip3_ob_out.tdata [48]);
tran (kme_cddip3_ob_out[47], \kme_cddip3_ob_out.tdata [47]);
tran (kme_cddip3_ob_out[46], \kme_cddip3_ob_out.tdata [46]);
tran (kme_cddip3_ob_out[45], \kme_cddip3_ob_out.tdata [45]);
tran (kme_cddip3_ob_out[44], \kme_cddip3_ob_out.tdata [44]);
tran (kme_cddip3_ob_out[43], \kme_cddip3_ob_out.tdata [43]);
tran (kme_cddip3_ob_out[42], \kme_cddip3_ob_out.tdata [42]);
tran (kme_cddip3_ob_out[41], \kme_cddip3_ob_out.tdata [41]);
tran (kme_cddip3_ob_out[40], \kme_cddip3_ob_out.tdata [40]);
tran (kme_cddip3_ob_out[39], \kme_cddip3_ob_out.tdata [39]);
tran (kme_cddip3_ob_out[38], \kme_cddip3_ob_out.tdata [38]);
tran (kme_cddip3_ob_out[37], \kme_cddip3_ob_out.tdata [37]);
tran (kme_cddip3_ob_out[36], \kme_cddip3_ob_out.tdata [36]);
tran (kme_cddip3_ob_out[35], \kme_cddip3_ob_out.tdata [35]);
tran (kme_cddip3_ob_out[34], \kme_cddip3_ob_out.tdata [34]);
tran (kme_cddip3_ob_out[33], \kme_cddip3_ob_out.tdata [33]);
tran (kme_cddip3_ob_out[32], \kme_cddip3_ob_out.tdata [32]);
tran (kme_cddip3_ob_out[31], \kme_cddip3_ob_out.tdata [31]);
tran (kme_cddip3_ob_out[30], \kme_cddip3_ob_out.tdata [30]);
tran (kme_cddip3_ob_out[29], \kme_cddip3_ob_out.tdata [29]);
tran (kme_cddip3_ob_out[28], \kme_cddip3_ob_out.tdata [28]);
tran (kme_cddip3_ob_out[27], \kme_cddip3_ob_out.tdata [27]);
tran (kme_cddip3_ob_out[26], \kme_cddip3_ob_out.tdata [26]);
tran (kme_cddip3_ob_out[25], \kme_cddip3_ob_out.tdata [25]);
tran (kme_cddip3_ob_out[24], \kme_cddip3_ob_out.tdata [24]);
tran (kme_cddip3_ob_out[23], \kme_cddip3_ob_out.tdata [23]);
tran (kme_cddip3_ob_out[22], \kme_cddip3_ob_out.tdata [22]);
tran (kme_cddip3_ob_out[21], \kme_cddip3_ob_out.tdata [21]);
tran (kme_cddip3_ob_out[20], \kme_cddip3_ob_out.tdata [20]);
tran (kme_cddip3_ob_out[19], \kme_cddip3_ob_out.tdata [19]);
tran (kme_cddip3_ob_out[18], \kme_cddip3_ob_out.tdata [18]);
tran (kme_cddip3_ob_out[17], \kme_cddip3_ob_out.tdata [17]);
tran (kme_cddip3_ob_out[16], \kme_cddip3_ob_out.tdata [16]);
tran (kme_cddip3_ob_out[15], \kme_cddip3_ob_out.tdata [15]);
tran (kme_cddip3_ob_out[14], \kme_cddip3_ob_out.tdata [14]);
tran (kme_cddip3_ob_out[13], \kme_cddip3_ob_out.tdata [13]);
tran (kme_cddip3_ob_out[12], \kme_cddip3_ob_out.tdata [12]);
tran (kme_cddip3_ob_out[11], \kme_cddip3_ob_out.tdata [11]);
tran (kme_cddip3_ob_out[10], \kme_cddip3_ob_out.tdata [10]);
tran (kme_cddip3_ob_out[9], \kme_cddip3_ob_out.tdata [9]);
tran (kme_cddip3_ob_out[8], \kme_cddip3_ob_out.tdata [8]);
tran (kme_cddip3_ob_out[7], \kme_cddip3_ob_out.tdata [7]);
tran (kme_cddip3_ob_out[6], \kme_cddip3_ob_out.tdata [6]);
tran (kme_cddip3_ob_out[5], \kme_cddip3_ob_out.tdata [5]);
tran (kme_cddip3_ob_out[4], \kme_cddip3_ob_out.tdata [4]);
tran (kme_cddip3_ob_out[3], \kme_cddip3_ob_out.tdata [3]);
tran (kme_cddip3_ob_out[2], \kme_cddip3_ob_out.tdata [2]);
tran (kme_cddip3_ob_out[1], \kme_cddip3_ob_out.tdata [1]);
tran (kme_cddip3_ob_out[0], \kme_cddip3_ob_out.tdata [0]);
tran (kme_cddip3_ob_in_mod[0], \kme_cddip3_ob_in_mod.tready );
tran (kim_dout[37], \kim_dout.valid [0]);
tran (kim_dout[36], \kim_dout.label_index [2]);
tran (kim_dout[35], \kim_dout.label_index [1]);
tran (kim_dout[34], \kim_dout.label_index [0]);
tran (kim_dout[33], \kim_dout.ckv_length [1]);
tran (kim_dout[32], \kim_dout.ckv_length [0]);
tran (kim_dout[31], \kim_dout.ckv_pointer [14]);
tran (kim_dout[30], \kim_dout.ckv_pointer [13]);
tran (kim_dout[29], \kim_dout.ckv_pointer [12]);
tran (kim_dout[28], \kim_dout.ckv_pointer [11]);
tran (kim_dout[27], \kim_dout.ckv_pointer [10]);
tran (kim_dout[26], \kim_dout.ckv_pointer [9]);
tran (kim_dout[25], \kim_dout.ckv_pointer [8]);
tran (kim_dout[24], \kim_dout.ckv_pointer [7]);
tran (kim_dout[23], \kim_dout.ckv_pointer [6]);
tran (kim_dout[22], \kim_dout.ckv_pointer [5]);
tran (kim_dout[21], \kim_dout.ckv_pointer [4]);
tran (kim_dout[20], \kim_dout.ckv_pointer [3]);
tran (kim_dout[19], \kim_dout.ckv_pointer [2]);
tran (kim_dout[18], \kim_dout.ckv_pointer [1]);
tran (kim_dout[17], \kim_dout.ckv_pointer [0]);
tran (kim_dout[16], \kim_dout.pf_num [3]);
tran (kim_dout[15], \kim_dout.pf_num [2]);
tran (kim_dout[14], \kim_dout.pf_num [1]);
tran (kim_dout[13], \kim_dout.pf_num [0]);
tran (kim_dout[12], \kim_dout.vf_num [11]);
tran (kim_dout[11], \kim_dout.vf_num [10]);
tran (kim_dout[10], \kim_dout.vf_num [9]);
tran (kim_dout[9], \kim_dout.vf_num [8]);
tran (kim_dout[8], \kim_dout.vf_num [7]);
tran (kim_dout[7], \kim_dout.vf_num [6]);
tran (kim_dout[6], \kim_dout.vf_num [5]);
tran (kim_dout[5], \kim_dout.vf_num [4]);
tran (kim_dout[4], \kim_dout.vf_num [3]);
tran (kim_dout[3], \kim_dout.vf_num [2]);
tran (kim_dout[2], \kim_dout.vf_num [1]);
tran (kim_dout[1], \kim_dout.vf_num [0]);
tran (kim_dout[0], \kim_dout.vf_valid [0]);
tran (\labels[7][271] , \labels[7].guid_size[0] );
tran (\labels[7][270] , \labels[7].label_size[5] );
tran (\labels[7][269] , \labels[7].label_size[4] );
tran (\labels[7][268] , \labels[7].label_size[3] );
tran (\labels[7][267] , \labels[7].label_size[2] );
tran (\labels[7][266] , \labels[7].label_size[1] );
tran (\labels[7][265] , \labels[7].label_size[0] );
tran (\labels[7][264] , \labels[7].label[255] );
tran (\labels[7][263] , \labels[7].label[254] );
tran (\labels[7][262] , \labels[7].label[253] );
tran (\labels[7][261] , \labels[7].label[252] );
tran (\labels[7][260] , \labels[7].label[251] );
tran (\labels[7][259] , \labels[7].label[250] );
tran (\labels[7][258] , \labels[7].label[249] );
tran (\labels[7][257] , \labels[7].label[248] );
tran (\labels[7][256] , \labels[7].label[247] );
tran (\labels[7][255] , \labels[7].label[246] );
tran (\labels[7][254] , \labels[7].label[245] );
tran (\labels[7][253] , \labels[7].label[244] );
tran (\labels[7][252] , \labels[7].label[243] );
tran (\labels[7][251] , \labels[7].label[242] );
tran (\labels[7][250] , \labels[7].label[241] );
tran (\labels[7][249] , \labels[7].label[240] );
tran (\labels[7][248] , \labels[7].label[239] );
tran (\labels[7][247] , \labels[7].label[238] );
tran (\labels[7][246] , \labels[7].label[237] );
tran (\labels[7][245] , \labels[7].label[236] );
tran (\labels[7][244] , \labels[7].label[235] );
tran (\labels[7][243] , \labels[7].label[234] );
tran (\labels[7][242] , \labels[7].label[233] );
tran (\labels[7][241] , \labels[7].label[232] );
tran (\labels[7][240] , \labels[7].label[231] );
tran (\labels[7][239] , \labels[7].label[230] );
tran (\labels[7][238] , \labels[7].label[229] );
tran (\labels[7][237] , \labels[7].label[228] );
tran (\labels[7][236] , \labels[7].label[227] );
tran (\labels[7][235] , \labels[7].label[226] );
tran (\labels[7][234] , \labels[7].label[225] );
tran (\labels[7][233] , \labels[7].label[224] );
tran (\labels[7][232] , \labels[7].label[223] );
tran (\labels[7][231] , \labels[7].label[222] );
tran (\labels[7][230] , \labels[7].label[221] );
tran (\labels[7][229] , \labels[7].label[220] );
tran (\labels[7][228] , \labels[7].label[219] );
tran (\labels[7][227] , \labels[7].label[218] );
tran (\labels[7][226] , \labels[7].label[217] );
tran (\labels[7][225] , \labels[7].label[216] );
tran (\labels[7][224] , \labels[7].label[215] );
tran (\labels[7][223] , \labels[7].label[214] );
tran (\labels[7][222] , \labels[7].label[213] );
tran (\labels[7][221] , \labels[7].label[212] );
tran (\labels[7][220] , \labels[7].label[211] );
tran (\labels[7][219] , \labels[7].label[210] );
tran (\labels[7][218] , \labels[7].label[209] );
tran (\labels[7][217] , \labels[7].label[208] );
tran (\labels[7][216] , \labels[7].label[207] );
tran (\labels[7][215] , \labels[7].label[206] );
tran (\labels[7][214] , \labels[7].label[205] );
tran (\labels[7][213] , \labels[7].label[204] );
tran (\labels[7][212] , \labels[7].label[203] );
tran (\labels[7][211] , \labels[7].label[202] );
tran (\labels[7][210] , \labels[7].label[201] );
tran (\labels[7][209] , \labels[7].label[200] );
tran (\labels[7][208] , \labels[7].label[199] );
tran (\labels[7][207] , \labels[7].label[198] );
tran (\labels[7][206] , \labels[7].label[197] );
tran (\labels[7][205] , \labels[7].label[196] );
tran (\labels[7][204] , \labels[7].label[195] );
tran (\labels[7][203] , \labels[7].label[194] );
tran (\labels[7][202] , \labels[7].label[193] );
tran (\labels[7][201] , \labels[7].label[192] );
tran (\labels[7][200] , \labels[7].label[191] );
tran (\labels[7][199] , \labels[7].label[190] );
tran (\labels[7][198] , \labels[7].label[189] );
tran (\labels[7][197] , \labels[7].label[188] );
tran (\labels[7][196] , \labels[7].label[187] );
tran (\labels[7][195] , \labels[7].label[186] );
tran (\labels[7][194] , \labels[7].label[185] );
tran (\labels[7][193] , \labels[7].label[184] );
tran (\labels[7][192] , \labels[7].label[183] );
tran (\labels[7][191] , \labels[7].label[182] );
tran (\labels[7][190] , \labels[7].label[181] );
tran (\labels[7][189] , \labels[7].label[180] );
tran (\labels[7][188] , \labels[7].label[179] );
tran (\labels[7][187] , \labels[7].label[178] );
tran (\labels[7][186] , \labels[7].label[177] );
tran (\labels[7][185] , \labels[7].label[176] );
tran (\labels[7][184] , \labels[7].label[175] );
tran (\labels[7][183] , \labels[7].label[174] );
tran (\labels[7][182] , \labels[7].label[173] );
tran (\labels[7][181] , \labels[7].label[172] );
tran (\labels[7][180] , \labels[7].label[171] );
tran (\labels[7][179] , \labels[7].label[170] );
tran (\labels[7][178] , \labels[7].label[169] );
tran (\labels[7][177] , \labels[7].label[168] );
tran (\labels[7][176] , \labels[7].label[167] );
tran (\labels[7][175] , \labels[7].label[166] );
tran (\labels[7][174] , \labels[7].label[165] );
tran (\labels[7][173] , \labels[7].label[164] );
tran (\labels[7][172] , \labels[7].label[163] );
tran (\labels[7][171] , \labels[7].label[162] );
tran (\labels[7][170] , \labels[7].label[161] );
tran (\labels[7][169] , \labels[7].label[160] );
tran (\labels[7][168] , \labels[7].label[159] );
tran (\labels[7][167] , \labels[7].label[158] );
tran (\labels[7][166] , \labels[7].label[157] );
tran (\labels[7][165] , \labels[7].label[156] );
tran (\labels[7][164] , \labels[7].label[155] );
tran (\labels[7][163] , \labels[7].label[154] );
tran (\labels[7][162] , \labels[7].label[153] );
tran (\labels[7][161] , \labels[7].label[152] );
tran (\labels[7][160] , \labels[7].label[151] );
tran (\labels[7][159] , \labels[7].label[150] );
tran (\labels[7][158] , \labels[7].label[149] );
tran (\labels[7][157] , \labels[7].label[148] );
tran (\labels[7][156] , \labels[7].label[147] );
tran (\labels[7][155] , \labels[7].label[146] );
tran (\labels[7][154] , \labels[7].label[145] );
tran (\labels[7][153] , \labels[7].label[144] );
tran (\labels[7][152] , \labels[7].label[143] );
tran (\labels[7][151] , \labels[7].label[142] );
tran (\labels[7][150] , \labels[7].label[141] );
tran (\labels[7][149] , \labels[7].label[140] );
tran (\labels[7][148] , \labels[7].label[139] );
tran (\labels[7][147] , \labels[7].label[138] );
tran (\labels[7][146] , \labels[7].label[137] );
tran (\labels[7][145] , \labels[7].label[136] );
tran (\labels[7][144] , \labels[7].label[135] );
tran (\labels[7][143] , \labels[7].label[134] );
tran (\labels[7][142] , \labels[7].label[133] );
tran (\labels[7][141] , \labels[7].label[132] );
tran (\labels[7][140] , \labels[7].label[131] );
tran (\labels[7][139] , \labels[7].label[130] );
tran (\labels[7][138] , \labels[7].label[129] );
tran (\labels[7][137] , \labels[7].label[128] );
tran (\labels[7][136] , \labels[7].label[127] );
tran (\labels[7][135] , \labels[7].label[126] );
tran (\labels[7][134] , \labels[7].label[125] );
tran (\labels[7][133] , \labels[7].label[124] );
tran (\labels[7][132] , \labels[7].label[123] );
tran (\labels[7][131] , \labels[7].label[122] );
tran (\labels[7][130] , \labels[7].label[121] );
tran (\labels[7][129] , \labels[7].label[120] );
tran (\labels[7][128] , \labels[7].label[119] );
tran (\labels[7][127] , \labels[7].label[118] );
tran (\labels[7][126] , \labels[7].label[117] );
tran (\labels[7][125] , \labels[7].label[116] );
tran (\labels[7][124] , \labels[7].label[115] );
tran (\labels[7][123] , \labels[7].label[114] );
tran (\labels[7][122] , \labels[7].label[113] );
tran (\labels[7][121] , \labels[7].label[112] );
tran (\labels[7][120] , \labels[7].label[111] );
tran (\labels[7][119] , \labels[7].label[110] );
tran (\labels[7][118] , \labels[7].label[109] );
tran (\labels[7][117] , \labels[7].label[108] );
tran (\labels[7][116] , \labels[7].label[107] );
tran (\labels[7][115] , \labels[7].label[106] );
tran (\labels[7][114] , \labels[7].label[105] );
tran (\labels[7][113] , \labels[7].label[104] );
tran (\labels[7][112] , \labels[7].label[103] );
tran (\labels[7][111] , \labels[7].label[102] );
tran (\labels[7][110] , \labels[7].label[101] );
tran (\labels[7][109] , \labels[7].label[100] );
tran (\labels[7][108] , \labels[7].label[99] );
tran (\labels[7][107] , \labels[7].label[98] );
tran (\labels[7][106] , \labels[7].label[97] );
tran (\labels[7][105] , \labels[7].label[96] );
tran (\labels[7][104] , \labels[7].label[95] );
tran (\labels[7][103] , \labels[7].label[94] );
tran (\labels[7][102] , \labels[7].label[93] );
tran (\labels[7][101] , \labels[7].label[92] );
tran (\labels[7][100] , \labels[7].label[91] );
tran (\labels[7][99] , \labels[7].label[90] );
tran (\labels[7][98] , \labels[7].label[89] );
tran (\labels[7][97] , \labels[7].label[88] );
tran (\labels[7][96] , \labels[7].label[87] );
tran (\labels[7][95] , \labels[7].label[86] );
tran (\labels[7][94] , \labels[7].label[85] );
tran (\labels[7][93] , \labels[7].label[84] );
tran (\labels[7][92] , \labels[7].label[83] );
tran (\labels[7][91] , \labels[7].label[82] );
tran (\labels[7][90] , \labels[7].label[81] );
tran (\labels[7][89] , \labels[7].label[80] );
tran (\labels[7][88] , \labels[7].label[79] );
tran (\labels[7][87] , \labels[7].label[78] );
tran (\labels[7][86] , \labels[7].label[77] );
tran (\labels[7][85] , \labels[7].label[76] );
tran (\labels[7][84] , \labels[7].label[75] );
tran (\labels[7][83] , \labels[7].label[74] );
tran (\labels[7][82] , \labels[7].label[73] );
tran (\labels[7][81] , \labels[7].label[72] );
tran (\labels[7][80] , \labels[7].label[71] );
tran (\labels[7][79] , \labels[7].label[70] );
tran (\labels[7][78] , \labels[7].label[69] );
tran (\labels[7][77] , \labels[7].label[68] );
tran (\labels[7][76] , \labels[7].label[67] );
tran (\labels[7][75] , \labels[7].label[66] );
tran (\labels[7][74] , \labels[7].label[65] );
tran (\labels[7][73] , \labels[7].label[64] );
tran (\labels[7][72] , \labels[7].label[63] );
tran (\labels[7][71] , \labels[7].label[62] );
tran (\labels[7][70] , \labels[7].label[61] );
tran (\labels[7][69] , \labels[7].label[60] );
tran (\labels[7][68] , \labels[7].label[59] );
tran (\labels[7][67] , \labels[7].label[58] );
tran (\labels[7][66] , \labels[7].label[57] );
tran (\labels[7][65] , \labels[7].label[56] );
tran (\labels[7][64] , \labels[7].label[55] );
tran (\labels[7][63] , \labels[7].label[54] );
tran (\labels[7][62] , \labels[7].label[53] );
tran (\labels[7][61] , \labels[7].label[52] );
tran (\labels[7][60] , \labels[7].label[51] );
tran (\labels[7][59] , \labels[7].label[50] );
tran (\labels[7][58] , \labels[7].label[49] );
tran (\labels[7][57] , \labels[7].label[48] );
tran (\labels[7][56] , \labels[7].label[47] );
tran (\labels[7][55] , \labels[7].label[46] );
tran (\labels[7][54] , \labels[7].label[45] );
tran (\labels[7][53] , \labels[7].label[44] );
tran (\labels[7][52] , \labels[7].label[43] );
tran (\labels[7][51] , \labels[7].label[42] );
tran (\labels[7][50] , \labels[7].label[41] );
tran (\labels[7][49] , \labels[7].label[40] );
tran (\labels[7][48] , \labels[7].label[39] );
tran (\labels[7][47] , \labels[7].label[38] );
tran (\labels[7][46] , \labels[7].label[37] );
tran (\labels[7][45] , \labels[7].label[36] );
tran (\labels[7][44] , \labels[7].label[35] );
tran (\labels[7][43] , \labels[7].label[34] );
tran (\labels[7][42] , \labels[7].label[33] );
tran (\labels[7][41] , \labels[7].label[32] );
tran (\labels[7][40] , \labels[7].label[31] );
tran (\labels[7][39] , \labels[7].label[30] );
tran (\labels[7][38] , \labels[7].label[29] );
tran (\labels[7][37] , \labels[7].label[28] );
tran (\labels[7][36] , \labels[7].label[27] );
tran (\labels[7][35] , \labels[7].label[26] );
tran (\labels[7][34] , \labels[7].label[25] );
tran (\labels[7][33] , \labels[7].label[24] );
tran (\labels[7][32] , \labels[7].label[23] );
tran (\labels[7][31] , \labels[7].label[22] );
tran (\labels[7][30] , \labels[7].label[21] );
tran (\labels[7][29] , \labels[7].label[20] );
tran (\labels[7][28] , \labels[7].label[19] );
tran (\labels[7][27] , \labels[7].label[18] );
tran (\labels[7][26] , \labels[7].label[17] );
tran (\labels[7][25] , \labels[7].label[16] );
tran (\labels[7][24] , \labels[7].label[15] );
tran (\labels[7][23] , \labels[7].label[14] );
tran (\labels[7][22] , \labels[7].label[13] );
tran (\labels[7][21] , \labels[7].label[12] );
tran (\labels[7][20] , \labels[7].label[11] );
tran (\labels[7][19] , \labels[7].label[10] );
tran (\labels[7][18] , \labels[7].label[9] );
tran (\labels[7][17] , \labels[7].label[8] );
tran (\labels[7][16] , \labels[7].label[7] );
tran (\labels[7][15] , \labels[7].label[6] );
tran (\labels[7][14] , \labels[7].label[5] );
tran (\labels[7][13] , \labels[7].label[4] );
tran (\labels[7][12] , \labels[7].label[3] );
tran (\labels[7][11] , \labels[7].label[2] );
tran (\labels[7][10] , \labels[7].label[1] );
tran (\labels[7][9] , \labels[7].label[0] );
tran (\labels[7][8] , \labels[7].delimiter_valid[0] );
tran (\labels[7][7] , \labels[7].delimiter[7] );
tran (\labels[7][6] , \labels[7].delimiter[6] );
tran (\labels[7][5] , \labels[7].delimiter[5] );
tran (\labels[7][4] , \labels[7].delimiter[4] );
tran (\labels[7][3] , \labels[7].delimiter[3] );
tran (\labels[7][2] , \labels[7].delimiter[2] );
tran (\labels[7][1] , \labels[7].delimiter[1] );
tran (\labels[7][0] , \labels[7].delimiter[0] );
tran (\labels[6][271] , \labels[6].guid_size[0] );
tran (\labels[6][270] , \labels[6].label_size[5] );
tran (\labels[6][269] , \labels[6].label_size[4] );
tran (\labels[6][268] , \labels[6].label_size[3] );
tran (\labels[6][267] , \labels[6].label_size[2] );
tran (\labels[6][266] , \labels[6].label_size[1] );
tran (\labels[6][265] , \labels[6].label_size[0] );
tran (\labels[6][264] , \labels[6].label[255] );
tran (\labels[6][263] , \labels[6].label[254] );
tran (\labels[6][262] , \labels[6].label[253] );
tran (\labels[6][261] , \labels[6].label[252] );
tran (\labels[6][260] , \labels[6].label[251] );
tran (\labels[6][259] , \labels[6].label[250] );
tran (\labels[6][258] , \labels[6].label[249] );
tran (\labels[6][257] , \labels[6].label[248] );
tran (\labels[6][256] , \labels[6].label[247] );
tran (\labels[6][255] , \labels[6].label[246] );
tran (\labels[6][254] , \labels[6].label[245] );
tran (\labels[6][253] , \labels[6].label[244] );
tran (\labels[6][252] , \labels[6].label[243] );
tran (\labels[6][251] , \labels[6].label[242] );
tran (\labels[6][250] , \labels[6].label[241] );
tran (\labels[6][249] , \labels[6].label[240] );
tran (\labels[6][248] , \labels[6].label[239] );
tran (\labels[6][247] , \labels[6].label[238] );
tran (\labels[6][246] , \labels[6].label[237] );
tran (\labels[6][245] , \labels[6].label[236] );
tran (\labels[6][244] , \labels[6].label[235] );
tran (\labels[6][243] , \labels[6].label[234] );
tran (\labels[6][242] , \labels[6].label[233] );
tran (\labels[6][241] , \labels[6].label[232] );
tran (\labels[6][240] , \labels[6].label[231] );
tran (\labels[6][239] , \labels[6].label[230] );
tran (\labels[6][238] , \labels[6].label[229] );
tran (\labels[6][237] , \labels[6].label[228] );
tran (\labels[6][236] , \labels[6].label[227] );
tran (\labels[6][235] , \labels[6].label[226] );
tran (\labels[6][234] , \labels[6].label[225] );
tran (\labels[6][233] , \labels[6].label[224] );
tran (\labels[6][232] , \labels[6].label[223] );
tran (\labels[6][231] , \labels[6].label[222] );
tran (\labels[6][230] , \labels[6].label[221] );
tran (\labels[6][229] , \labels[6].label[220] );
tran (\labels[6][228] , \labels[6].label[219] );
tran (\labels[6][227] , \labels[6].label[218] );
tran (\labels[6][226] , \labels[6].label[217] );
tran (\labels[6][225] , \labels[6].label[216] );
tran (\labels[6][224] , \labels[6].label[215] );
tran (\labels[6][223] , \labels[6].label[214] );
tran (\labels[6][222] , \labels[6].label[213] );
tran (\labels[6][221] , \labels[6].label[212] );
tran (\labels[6][220] , \labels[6].label[211] );
tran (\labels[6][219] , \labels[6].label[210] );
tran (\labels[6][218] , \labels[6].label[209] );
tran (\labels[6][217] , \labels[6].label[208] );
tran (\labels[6][216] , \labels[6].label[207] );
tran (\labels[6][215] , \labels[6].label[206] );
tran (\labels[6][214] , \labels[6].label[205] );
tran (\labels[6][213] , \labels[6].label[204] );
tran (\labels[6][212] , \labels[6].label[203] );
tran (\labels[6][211] , \labels[6].label[202] );
tran (\labels[6][210] , \labels[6].label[201] );
tran (\labels[6][209] , \labels[6].label[200] );
tran (\labels[6][208] , \labels[6].label[199] );
tran (\labels[6][207] , \labels[6].label[198] );
tran (\labels[6][206] , \labels[6].label[197] );
tran (\labels[6][205] , \labels[6].label[196] );
tran (\labels[6][204] , \labels[6].label[195] );
tran (\labels[6][203] , \labels[6].label[194] );
tran (\labels[6][202] , \labels[6].label[193] );
tran (\labels[6][201] , \labels[6].label[192] );
tran (\labels[6][200] , \labels[6].label[191] );
tran (\labels[6][199] , \labels[6].label[190] );
tran (\labels[6][198] , \labels[6].label[189] );
tran (\labels[6][197] , \labels[6].label[188] );
tran (\labels[6][196] , \labels[6].label[187] );
tran (\labels[6][195] , \labels[6].label[186] );
tran (\labels[6][194] , \labels[6].label[185] );
tran (\labels[6][193] , \labels[6].label[184] );
tran (\labels[6][192] , \labels[6].label[183] );
tran (\labels[6][191] , \labels[6].label[182] );
tran (\labels[6][190] , \labels[6].label[181] );
tran (\labels[6][189] , \labels[6].label[180] );
tran (\labels[6][188] , \labels[6].label[179] );
tran (\labels[6][187] , \labels[6].label[178] );
tran (\labels[6][186] , \labels[6].label[177] );
tran (\labels[6][185] , \labels[6].label[176] );
tran (\labels[6][184] , \labels[6].label[175] );
tran (\labels[6][183] , \labels[6].label[174] );
tran (\labels[6][182] , \labels[6].label[173] );
tran (\labels[6][181] , \labels[6].label[172] );
tran (\labels[6][180] , \labels[6].label[171] );
tran (\labels[6][179] , \labels[6].label[170] );
tran (\labels[6][178] , \labels[6].label[169] );
tran (\labels[6][177] , \labels[6].label[168] );
tran (\labels[6][176] , \labels[6].label[167] );
tran (\labels[6][175] , \labels[6].label[166] );
tran (\labels[6][174] , \labels[6].label[165] );
tran (\labels[6][173] , \labels[6].label[164] );
tran (\labels[6][172] , \labels[6].label[163] );
tran (\labels[6][171] , \labels[6].label[162] );
tran (\labels[6][170] , \labels[6].label[161] );
tran (\labels[6][169] , \labels[6].label[160] );
tran (\labels[6][168] , \labels[6].label[159] );
tran (\labels[6][167] , \labels[6].label[158] );
tran (\labels[6][166] , \labels[6].label[157] );
tran (\labels[6][165] , \labels[6].label[156] );
tran (\labels[6][164] , \labels[6].label[155] );
tran (\labels[6][163] , \labels[6].label[154] );
tran (\labels[6][162] , \labels[6].label[153] );
tran (\labels[6][161] , \labels[6].label[152] );
tran (\labels[6][160] , \labels[6].label[151] );
tran (\labels[6][159] , \labels[6].label[150] );
tran (\labels[6][158] , \labels[6].label[149] );
tran (\labels[6][157] , \labels[6].label[148] );
tran (\labels[6][156] , \labels[6].label[147] );
tran (\labels[6][155] , \labels[6].label[146] );
tran (\labels[6][154] , \labels[6].label[145] );
tran (\labels[6][153] , \labels[6].label[144] );
tran (\labels[6][152] , \labels[6].label[143] );
tran (\labels[6][151] , \labels[6].label[142] );
tran (\labels[6][150] , \labels[6].label[141] );
tran (\labels[6][149] , \labels[6].label[140] );
tran (\labels[6][148] , \labels[6].label[139] );
tran (\labels[6][147] , \labels[6].label[138] );
tran (\labels[6][146] , \labels[6].label[137] );
tran (\labels[6][145] , \labels[6].label[136] );
tran (\labels[6][144] , \labels[6].label[135] );
tran (\labels[6][143] , \labels[6].label[134] );
tran (\labels[6][142] , \labels[6].label[133] );
tran (\labels[6][141] , \labels[6].label[132] );
tran (\labels[6][140] , \labels[6].label[131] );
tran (\labels[6][139] , \labels[6].label[130] );
tran (\labels[6][138] , \labels[6].label[129] );
tran (\labels[6][137] , \labels[6].label[128] );
tran (\labels[6][136] , \labels[6].label[127] );
tran (\labels[6][135] , \labels[6].label[126] );
tran (\labels[6][134] , \labels[6].label[125] );
tran (\labels[6][133] , \labels[6].label[124] );
tran (\labels[6][132] , \labels[6].label[123] );
tran (\labels[6][131] , \labels[6].label[122] );
tran (\labels[6][130] , \labels[6].label[121] );
tran (\labels[6][129] , \labels[6].label[120] );
tran (\labels[6][128] , \labels[6].label[119] );
tran (\labels[6][127] , \labels[6].label[118] );
tran (\labels[6][126] , \labels[6].label[117] );
tran (\labels[6][125] , \labels[6].label[116] );
tran (\labels[6][124] , \labels[6].label[115] );
tran (\labels[6][123] , \labels[6].label[114] );
tran (\labels[6][122] , \labels[6].label[113] );
tran (\labels[6][121] , \labels[6].label[112] );
tran (\labels[6][120] , \labels[6].label[111] );
tran (\labels[6][119] , \labels[6].label[110] );
tran (\labels[6][118] , \labels[6].label[109] );
tran (\labels[6][117] , \labels[6].label[108] );
tran (\labels[6][116] , \labels[6].label[107] );
tran (\labels[6][115] , \labels[6].label[106] );
tran (\labels[6][114] , \labels[6].label[105] );
tran (\labels[6][113] , \labels[6].label[104] );
tran (\labels[6][112] , \labels[6].label[103] );
tran (\labels[6][111] , \labels[6].label[102] );
tran (\labels[6][110] , \labels[6].label[101] );
tran (\labels[6][109] , \labels[6].label[100] );
tran (\labels[6][108] , \labels[6].label[99] );
tran (\labels[6][107] , \labels[6].label[98] );
tran (\labels[6][106] , \labels[6].label[97] );
tran (\labels[6][105] , \labels[6].label[96] );
tran (\labels[6][104] , \labels[6].label[95] );
tran (\labels[6][103] , \labels[6].label[94] );
tran (\labels[6][102] , \labels[6].label[93] );
tran (\labels[6][101] , \labels[6].label[92] );
tran (\labels[6][100] , \labels[6].label[91] );
tran (\labels[6][99] , \labels[6].label[90] );
tran (\labels[6][98] , \labels[6].label[89] );
tran (\labels[6][97] , \labels[6].label[88] );
tran (\labels[6][96] , \labels[6].label[87] );
tran (\labels[6][95] , \labels[6].label[86] );
tran (\labels[6][94] , \labels[6].label[85] );
tran (\labels[6][93] , \labels[6].label[84] );
tran (\labels[6][92] , \labels[6].label[83] );
tran (\labels[6][91] , \labels[6].label[82] );
tran (\labels[6][90] , \labels[6].label[81] );
tran (\labels[6][89] , \labels[6].label[80] );
tran (\labels[6][88] , \labels[6].label[79] );
tran (\labels[6][87] , \labels[6].label[78] );
tran (\labels[6][86] , \labels[6].label[77] );
tran (\labels[6][85] , \labels[6].label[76] );
tran (\labels[6][84] , \labels[6].label[75] );
tran (\labels[6][83] , \labels[6].label[74] );
tran (\labels[6][82] , \labels[6].label[73] );
tran (\labels[6][81] , \labels[6].label[72] );
tran (\labels[6][80] , \labels[6].label[71] );
tran (\labels[6][79] , \labels[6].label[70] );
tran (\labels[6][78] , \labels[6].label[69] );
tran (\labels[6][77] , \labels[6].label[68] );
tran (\labels[6][76] , \labels[6].label[67] );
tran (\labels[6][75] , \labels[6].label[66] );
tran (\labels[6][74] , \labels[6].label[65] );
tran (\labels[6][73] , \labels[6].label[64] );
tran (\labels[6][72] , \labels[6].label[63] );
tran (\labels[6][71] , \labels[6].label[62] );
tran (\labels[6][70] , \labels[6].label[61] );
tran (\labels[6][69] , \labels[6].label[60] );
tran (\labels[6][68] , \labels[6].label[59] );
tran (\labels[6][67] , \labels[6].label[58] );
tran (\labels[6][66] , \labels[6].label[57] );
tran (\labels[6][65] , \labels[6].label[56] );
tran (\labels[6][64] , \labels[6].label[55] );
tran (\labels[6][63] , \labels[6].label[54] );
tran (\labels[6][62] , \labels[6].label[53] );
tran (\labels[6][61] , \labels[6].label[52] );
tran (\labels[6][60] , \labels[6].label[51] );
tran (\labels[6][59] , \labels[6].label[50] );
tran (\labels[6][58] , \labels[6].label[49] );
tran (\labels[6][57] , \labels[6].label[48] );
tran (\labels[6][56] , \labels[6].label[47] );
tran (\labels[6][55] , \labels[6].label[46] );
tran (\labels[6][54] , \labels[6].label[45] );
tran (\labels[6][53] , \labels[6].label[44] );
tran (\labels[6][52] , \labels[6].label[43] );
tran (\labels[6][51] , \labels[6].label[42] );
tran (\labels[6][50] , \labels[6].label[41] );
tran (\labels[6][49] , \labels[6].label[40] );
tran (\labels[6][48] , \labels[6].label[39] );
tran (\labels[6][47] , \labels[6].label[38] );
tran (\labels[6][46] , \labels[6].label[37] );
tran (\labels[6][45] , \labels[6].label[36] );
tran (\labels[6][44] , \labels[6].label[35] );
tran (\labels[6][43] , \labels[6].label[34] );
tran (\labels[6][42] , \labels[6].label[33] );
tran (\labels[6][41] , \labels[6].label[32] );
tran (\labels[6][40] , \labels[6].label[31] );
tran (\labels[6][39] , \labels[6].label[30] );
tran (\labels[6][38] , \labels[6].label[29] );
tran (\labels[6][37] , \labels[6].label[28] );
tran (\labels[6][36] , \labels[6].label[27] );
tran (\labels[6][35] , \labels[6].label[26] );
tran (\labels[6][34] , \labels[6].label[25] );
tran (\labels[6][33] , \labels[6].label[24] );
tran (\labels[6][32] , \labels[6].label[23] );
tran (\labels[6][31] , \labels[6].label[22] );
tran (\labels[6][30] , \labels[6].label[21] );
tran (\labels[6][29] , \labels[6].label[20] );
tran (\labels[6][28] , \labels[6].label[19] );
tran (\labels[6][27] , \labels[6].label[18] );
tran (\labels[6][26] , \labels[6].label[17] );
tran (\labels[6][25] , \labels[6].label[16] );
tran (\labels[6][24] , \labels[6].label[15] );
tran (\labels[6][23] , \labels[6].label[14] );
tran (\labels[6][22] , \labels[6].label[13] );
tran (\labels[6][21] , \labels[6].label[12] );
tran (\labels[6][20] , \labels[6].label[11] );
tran (\labels[6][19] , \labels[6].label[10] );
tran (\labels[6][18] , \labels[6].label[9] );
tran (\labels[6][17] , \labels[6].label[8] );
tran (\labels[6][16] , \labels[6].label[7] );
tran (\labels[6][15] , \labels[6].label[6] );
tran (\labels[6][14] , \labels[6].label[5] );
tran (\labels[6][13] , \labels[6].label[4] );
tran (\labels[6][12] , \labels[6].label[3] );
tran (\labels[6][11] , \labels[6].label[2] );
tran (\labels[6][10] , \labels[6].label[1] );
tran (\labels[6][9] , \labels[6].label[0] );
tran (\labels[6][8] , \labels[6].delimiter_valid[0] );
tran (\labels[6][7] , \labels[6].delimiter[7] );
tran (\labels[6][6] , \labels[6].delimiter[6] );
tran (\labels[6][5] , \labels[6].delimiter[5] );
tran (\labels[6][4] , \labels[6].delimiter[4] );
tran (\labels[6][3] , \labels[6].delimiter[3] );
tran (\labels[6][2] , \labels[6].delimiter[2] );
tran (\labels[6][1] , \labels[6].delimiter[1] );
tran (\labels[6][0] , \labels[6].delimiter[0] );
tran (\labels[5][271] , \labels[5].guid_size[0] );
tran (\labels[5][270] , \labels[5].label_size[5] );
tran (\labels[5][269] , \labels[5].label_size[4] );
tran (\labels[5][268] , \labels[5].label_size[3] );
tran (\labels[5][267] , \labels[5].label_size[2] );
tran (\labels[5][266] , \labels[5].label_size[1] );
tran (\labels[5][265] , \labels[5].label_size[0] );
tran (\labels[5][264] , \labels[5].label[255] );
tran (\labels[5][263] , \labels[5].label[254] );
tran (\labels[5][262] , \labels[5].label[253] );
tran (\labels[5][261] , \labels[5].label[252] );
tran (\labels[5][260] , \labels[5].label[251] );
tran (\labels[5][259] , \labels[5].label[250] );
tran (\labels[5][258] , \labels[5].label[249] );
tran (\labels[5][257] , \labels[5].label[248] );
tran (\labels[5][256] , \labels[5].label[247] );
tran (\labels[5][255] , \labels[5].label[246] );
tran (\labels[5][254] , \labels[5].label[245] );
tran (\labels[5][253] , \labels[5].label[244] );
tran (\labels[5][252] , \labels[5].label[243] );
tran (\labels[5][251] , \labels[5].label[242] );
tran (\labels[5][250] , \labels[5].label[241] );
tran (\labels[5][249] , \labels[5].label[240] );
tran (\labels[5][248] , \labels[5].label[239] );
tran (\labels[5][247] , \labels[5].label[238] );
tran (\labels[5][246] , \labels[5].label[237] );
tran (\labels[5][245] , \labels[5].label[236] );
tran (\labels[5][244] , \labels[5].label[235] );
tran (\labels[5][243] , \labels[5].label[234] );
tran (\labels[5][242] , \labels[5].label[233] );
tran (\labels[5][241] , \labels[5].label[232] );
tran (\labels[5][240] , \labels[5].label[231] );
tran (\labels[5][239] , \labels[5].label[230] );
tran (\labels[5][238] , \labels[5].label[229] );
tran (\labels[5][237] , \labels[5].label[228] );
tran (\labels[5][236] , \labels[5].label[227] );
tran (\labels[5][235] , \labels[5].label[226] );
tran (\labels[5][234] , \labels[5].label[225] );
tran (\labels[5][233] , \labels[5].label[224] );
tran (\labels[5][232] , \labels[5].label[223] );
tran (\labels[5][231] , \labels[5].label[222] );
tran (\labels[5][230] , \labels[5].label[221] );
tran (\labels[5][229] , \labels[5].label[220] );
tran (\labels[5][228] , \labels[5].label[219] );
tran (\labels[5][227] , \labels[5].label[218] );
tran (\labels[5][226] , \labels[5].label[217] );
tran (\labels[5][225] , \labels[5].label[216] );
tran (\labels[5][224] , \labels[5].label[215] );
tran (\labels[5][223] , \labels[5].label[214] );
tran (\labels[5][222] , \labels[5].label[213] );
tran (\labels[5][221] , \labels[5].label[212] );
tran (\labels[5][220] , \labels[5].label[211] );
tran (\labels[5][219] , \labels[5].label[210] );
tran (\labels[5][218] , \labels[5].label[209] );
tran (\labels[5][217] , \labels[5].label[208] );
tran (\labels[5][216] , \labels[5].label[207] );
tran (\labels[5][215] , \labels[5].label[206] );
tran (\labels[5][214] , \labels[5].label[205] );
tran (\labels[5][213] , \labels[5].label[204] );
tran (\labels[5][212] , \labels[5].label[203] );
tran (\labels[5][211] , \labels[5].label[202] );
tran (\labels[5][210] , \labels[5].label[201] );
tran (\labels[5][209] , \labels[5].label[200] );
tran (\labels[5][208] , \labels[5].label[199] );
tran (\labels[5][207] , \labels[5].label[198] );
tran (\labels[5][206] , \labels[5].label[197] );
tran (\labels[5][205] , \labels[5].label[196] );
tran (\labels[5][204] , \labels[5].label[195] );
tran (\labels[5][203] , \labels[5].label[194] );
tran (\labels[5][202] , \labels[5].label[193] );
tran (\labels[5][201] , \labels[5].label[192] );
tran (\labels[5][200] , \labels[5].label[191] );
tran (\labels[5][199] , \labels[5].label[190] );
tran (\labels[5][198] , \labels[5].label[189] );
tran (\labels[5][197] , \labels[5].label[188] );
tran (\labels[5][196] , \labels[5].label[187] );
tran (\labels[5][195] , \labels[5].label[186] );
tran (\labels[5][194] , \labels[5].label[185] );
tran (\labels[5][193] , \labels[5].label[184] );
tran (\labels[5][192] , \labels[5].label[183] );
tran (\labels[5][191] , \labels[5].label[182] );
tran (\labels[5][190] , \labels[5].label[181] );
tran (\labels[5][189] , \labels[5].label[180] );
tran (\labels[5][188] , \labels[5].label[179] );
tran (\labels[5][187] , \labels[5].label[178] );
tran (\labels[5][186] , \labels[5].label[177] );
tran (\labels[5][185] , \labels[5].label[176] );
tran (\labels[5][184] , \labels[5].label[175] );
tran (\labels[5][183] , \labels[5].label[174] );
tran (\labels[5][182] , \labels[5].label[173] );
tran (\labels[5][181] , \labels[5].label[172] );
tran (\labels[5][180] , \labels[5].label[171] );
tran (\labels[5][179] , \labels[5].label[170] );
tran (\labels[5][178] , \labels[5].label[169] );
tran (\labels[5][177] , \labels[5].label[168] );
tran (\labels[5][176] , \labels[5].label[167] );
tran (\labels[5][175] , \labels[5].label[166] );
tran (\labels[5][174] , \labels[5].label[165] );
tran (\labels[5][173] , \labels[5].label[164] );
tran (\labels[5][172] , \labels[5].label[163] );
tran (\labels[5][171] , \labels[5].label[162] );
tran (\labels[5][170] , \labels[5].label[161] );
tran (\labels[5][169] , \labels[5].label[160] );
tran (\labels[5][168] , \labels[5].label[159] );
tran (\labels[5][167] , \labels[5].label[158] );
tran (\labels[5][166] , \labels[5].label[157] );
tran (\labels[5][165] , \labels[5].label[156] );
tran (\labels[5][164] , \labels[5].label[155] );
tran (\labels[5][163] , \labels[5].label[154] );
tran (\labels[5][162] , \labels[5].label[153] );
tran (\labels[5][161] , \labels[5].label[152] );
tran (\labels[5][160] , \labels[5].label[151] );
tran (\labels[5][159] , \labels[5].label[150] );
tran (\labels[5][158] , \labels[5].label[149] );
tran (\labels[5][157] , \labels[5].label[148] );
tran (\labels[5][156] , \labels[5].label[147] );
tran (\labels[5][155] , \labels[5].label[146] );
tran (\labels[5][154] , \labels[5].label[145] );
tran (\labels[5][153] , \labels[5].label[144] );
tran (\labels[5][152] , \labels[5].label[143] );
tran (\labels[5][151] , \labels[5].label[142] );
tran (\labels[5][150] , \labels[5].label[141] );
tran (\labels[5][149] , \labels[5].label[140] );
tran (\labels[5][148] , \labels[5].label[139] );
tran (\labels[5][147] , \labels[5].label[138] );
tran (\labels[5][146] , \labels[5].label[137] );
tran (\labels[5][145] , \labels[5].label[136] );
tran (\labels[5][144] , \labels[5].label[135] );
tran (\labels[5][143] , \labels[5].label[134] );
tran (\labels[5][142] , \labels[5].label[133] );
tran (\labels[5][141] , \labels[5].label[132] );
tran (\labels[5][140] , \labels[5].label[131] );
tran (\labels[5][139] , \labels[5].label[130] );
tran (\labels[5][138] , \labels[5].label[129] );
tran (\labels[5][137] , \labels[5].label[128] );
tran (\labels[5][136] , \labels[5].label[127] );
tran (\labels[5][135] , \labels[5].label[126] );
tran (\labels[5][134] , \labels[5].label[125] );
tran (\labels[5][133] , \labels[5].label[124] );
tran (\labels[5][132] , \labels[5].label[123] );
tran (\labels[5][131] , \labels[5].label[122] );
tran (\labels[5][130] , \labels[5].label[121] );
tran (\labels[5][129] , \labels[5].label[120] );
tran (\labels[5][128] , \labels[5].label[119] );
tran (\labels[5][127] , \labels[5].label[118] );
tran (\labels[5][126] , \labels[5].label[117] );
tran (\labels[5][125] , \labels[5].label[116] );
tran (\labels[5][124] , \labels[5].label[115] );
tran (\labels[5][123] , \labels[5].label[114] );
tran (\labels[5][122] , \labels[5].label[113] );
tran (\labels[5][121] , \labels[5].label[112] );
tran (\labels[5][120] , \labels[5].label[111] );
tran (\labels[5][119] , \labels[5].label[110] );
tran (\labels[5][118] , \labels[5].label[109] );
tran (\labels[5][117] , \labels[5].label[108] );
tran (\labels[5][116] , \labels[5].label[107] );
tran (\labels[5][115] , \labels[5].label[106] );
tran (\labels[5][114] , \labels[5].label[105] );
tran (\labels[5][113] , \labels[5].label[104] );
tran (\labels[5][112] , \labels[5].label[103] );
tran (\labels[5][111] , \labels[5].label[102] );
tran (\labels[5][110] , \labels[5].label[101] );
tran (\labels[5][109] , \labels[5].label[100] );
tran (\labels[5][108] , \labels[5].label[99] );
tran (\labels[5][107] , \labels[5].label[98] );
tran (\labels[5][106] , \labels[5].label[97] );
tran (\labels[5][105] , \labels[5].label[96] );
tran (\labels[5][104] , \labels[5].label[95] );
tran (\labels[5][103] , \labels[5].label[94] );
tran (\labels[5][102] , \labels[5].label[93] );
tran (\labels[5][101] , \labels[5].label[92] );
tran (\labels[5][100] , \labels[5].label[91] );
tran (\labels[5][99] , \labels[5].label[90] );
tran (\labels[5][98] , \labels[5].label[89] );
tran (\labels[5][97] , \labels[5].label[88] );
tran (\labels[5][96] , \labels[5].label[87] );
tran (\labels[5][95] , \labels[5].label[86] );
tran (\labels[5][94] , \labels[5].label[85] );
tran (\labels[5][93] , \labels[5].label[84] );
tran (\labels[5][92] , \labels[5].label[83] );
tran (\labels[5][91] , \labels[5].label[82] );
tran (\labels[5][90] , \labels[5].label[81] );
tran (\labels[5][89] , \labels[5].label[80] );
tran (\labels[5][88] , \labels[5].label[79] );
tran (\labels[5][87] , \labels[5].label[78] );
tran (\labels[5][86] , \labels[5].label[77] );
tran (\labels[5][85] , \labels[5].label[76] );
tran (\labels[5][84] , \labels[5].label[75] );
tran (\labels[5][83] , \labels[5].label[74] );
tran (\labels[5][82] , \labels[5].label[73] );
tran (\labels[5][81] , \labels[5].label[72] );
tran (\labels[5][80] , \labels[5].label[71] );
tran (\labels[5][79] , \labels[5].label[70] );
tran (\labels[5][78] , \labels[5].label[69] );
tran (\labels[5][77] , \labels[5].label[68] );
tran (\labels[5][76] , \labels[5].label[67] );
tran (\labels[5][75] , \labels[5].label[66] );
tran (\labels[5][74] , \labels[5].label[65] );
tran (\labels[5][73] , \labels[5].label[64] );
tran (\labels[5][72] , \labels[5].label[63] );
tran (\labels[5][71] , \labels[5].label[62] );
tran (\labels[5][70] , \labels[5].label[61] );
tran (\labels[5][69] , \labels[5].label[60] );
tran (\labels[5][68] , \labels[5].label[59] );
tran (\labels[5][67] , \labels[5].label[58] );
tran (\labels[5][66] , \labels[5].label[57] );
tran (\labels[5][65] , \labels[5].label[56] );
tran (\labels[5][64] , \labels[5].label[55] );
tran (\labels[5][63] , \labels[5].label[54] );
tran (\labels[5][62] , \labels[5].label[53] );
tran (\labels[5][61] , \labels[5].label[52] );
tran (\labels[5][60] , \labels[5].label[51] );
tran (\labels[5][59] , \labels[5].label[50] );
tran (\labels[5][58] , \labels[5].label[49] );
tran (\labels[5][57] , \labels[5].label[48] );
tran (\labels[5][56] , \labels[5].label[47] );
tran (\labels[5][55] , \labels[5].label[46] );
tran (\labels[5][54] , \labels[5].label[45] );
tran (\labels[5][53] , \labels[5].label[44] );
tran (\labels[5][52] , \labels[5].label[43] );
tran (\labels[5][51] , \labels[5].label[42] );
tran (\labels[5][50] , \labels[5].label[41] );
tran (\labels[5][49] , \labels[5].label[40] );
tran (\labels[5][48] , \labels[5].label[39] );
tran (\labels[5][47] , \labels[5].label[38] );
tran (\labels[5][46] , \labels[5].label[37] );
tran (\labels[5][45] , \labels[5].label[36] );
tran (\labels[5][44] , \labels[5].label[35] );
tran (\labels[5][43] , \labels[5].label[34] );
tran (\labels[5][42] , \labels[5].label[33] );
tran (\labels[5][41] , \labels[5].label[32] );
tran (\labels[5][40] , \labels[5].label[31] );
tran (\labels[5][39] , \labels[5].label[30] );
tran (\labels[5][38] , \labels[5].label[29] );
tran (\labels[5][37] , \labels[5].label[28] );
tran (\labels[5][36] , \labels[5].label[27] );
tran (\labels[5][35] , \labels[5].label[26] );
tran (\labels[5][34] , \labels[5].label[25] );
tran (\labels[5][33] , \labels[5].label[24] );
tran (\labels[5][32] , \labels[5].label[23] );
tran (\labels[5][31] , \labels[5].label[22] );
tran (\labels[5][30] , \labels[5].label[21] );
tran (\labels[5][29] , \labels[5].label[20] );
tran (\labels[5][28] , \labels[5].label[19] );
tran (\labels[5][27] , \labels[5].label[18] );
tran (\labels[5][26] , \labels[5].label[17] );
tran (\labels[5][25] , \labels[5].label[16] );
tran (\labels[5][24] , \labels[5].label[15] );
tran (\labels[5][23] , \labels[5].label[14] );
tran (\labels[5][22] , \labels[5].label[13] );
tran (\labels[5][21] , \labels[5].label[12] );
tran (\labels[5][20] , \labels[5].label[11] );
tran (\labels[5][19] , \labels[5].label[10] );
tran (\labels[5][18] , \labels[5].label[9] );
tran (\labels[5][17] , \labels[5].label[8] );
tran (\labels[5][16] , \labels[5].label[7] );
tran (\labels[5][15] , \labels[5].label[6] );
tran (\labels[5][14] , \labels[5].label[5] );
tran (\labels[5][13] , \labels[5].label[4] );
tran (\labels[5][12] , \labels[5].label[3] );
tran (\labels[5][11] , \labels[5].label[2] );
tran (\labels[5][10] , \labels[5].label[1] );
tran (\labels[5][9] , \labels[5].label[0] );
tran (\labels[5][8] , \labels[5].delimiter_valid[0] );
tran (\labels[5][7] , \labels[5].delimiter[7] );
tran (\labels[5][6] , \labels[5].delimiter[6] );
tran (\labels[5][5] , \labels[5].delimiter[5] );
tran (\labels[5][4] , \labels[5].delimiter[4] );
tran (\labels[5][3] , \labels[5].delimiter[3] );
tran (\labels[5][2] , \labels[5].delimiter[2] );
tran (\labels[5][1] , \labels[5].delimiter[1] );
tran (\labels[5][0] , \labels[5].delimiter[0] );
tran (\labels[4][271] , \labels[4].guid_size[0] );
tran (\labels[4][270] , \labels[4].label_size[5] );
tran (\labels[4][269] , \labels[4].label_size[4] );
tran (\labels[4][268] , \labels[4].label_size[3] );
tran (\labels[4][267] , \labels[4].label_size[2] );
tran (\labels[4][266] , \labels[4].label_size[1] );
tran (\labels[4][265] , \labels[4].label_size[0] );
tran (\labels[4][264] , \labels[4].label[255] );
tran (\labels[4][263] , \labels[4].label[254] );
tran (\labels[4][262] , \labels[4].label[253] );
tran (\labels[4][261] , \labels[4].label[252] );
tran (\labels[4][260] , \labels[4].label[251] );
tran (\labels[4][259] , \labels[4].label[250] );
tran (\labels[4][258] , \labels[4].label[249] );
tran (\labels[4][257] , \labels[4].label[248] );
tran (\labels[4][256] , \labels[4].label[247] );
tran (\labels[4][255] , \labels[4].label[246] );
tran (\labels[4][254] , \labels[4].label[245] );
tran (\labels[4][253] , \labels[4].label[244] );
tran (\labels[4][252] , \labels[4].label[243] );
tran (\labels[4][251] , \labels[4].label[242] );
tran (\labels[4][250] , \labels[4].label[241] );
tran (\labels[4][249] , \labels[4].label[240] );
tran (\labels[4][248] , \labels[4].label[239] );
tran (\labels[4][247] , \labels[4].label[238] );
tran (\labels[4][246] , \labels[4].label[237] );
tran (\labels[4][245] , \labels[4].label[236] );
tran (\labels[4][244] , \labels[4].label[235] );
tran (\labels[4][243] , \labels[4].label[234] );
tran (\labels[4][242] , \labels[4].label[233] );
tran (\labels[4][241] , \labels[4].label[232] );
tran (\labels[4][240] , \labels[4].label[231] );
tran (\labels[4][239] , \labels[4].label[230] );
tran (\labels[4][238] , \labels[4].label[229] );
tran (\labels[4][237] , \labels[4].label[228] );
tran (\labels[4][236] , \labels[4].label[227] );
tran (\labels[4][235] , \labels[4].label[226] );
tran (\labels[4][234] , \labels[4].label[225] );
tran (\labels[4][233] , \labels[4].label[224] );
tran (\labels[4][232] , \labels[4].label[223] );
tran (\labels[4][231] , \labels[4].label[222] );
tran (\labels[4][230] , \labels[4].label[221] );
tran (\labels[4][229] , \labels[4].label[220] );
tran (\labels[4][228] , \labels[4].label[219] );
tran (\labels[4][227] , \labels[4].label[218] );
tran (\labels[4][226] , \labels[4].label[217] );
tran (\labels[4][225] , \labels[4].label[216] );
tran (\labels[4][224] , \labels[4].label[215] );
tran (\labels[4][223] , \labels[4].label[214] );
tran (\labels[4][222] , \labels[4].label[213] );
tran (\labels[4][221] , \labels[4].label[212] );
tran (\labels[4][220] , \labels[4].label[211] );
tran (\labels[4][219] , \labels[4].label[210] );
tran (\labels[4][218] , \labels[4].label[209] );
tran (\labels[4][217] , \labels[4].label[208] );
tran (\labels[4][216] , \labels[4].label[207] );
tran (\labels[4][215] , \labels[4].label[206] );
tran (\labels[4][214] , \labels[4].label[205] );
tran (\labels[4][213] , \labels[4].label[204] );
tran (\labels[4][212] , \labels[4].label[203] );
tran (\labels[4][211] , \labels[4].label[202] );
tran (\labels[4][210] , \labels[4].label[201] );
tran (\labels[4][209] , \labels[4].label[200] );
tran (\labels[4][208] , \labels[4].label[199] );
tran (\labels[4][207] , \labels[4].label[198] );
tran (\labels[4][206] , \labels[4].label[197] );
tran (\labels[4][205] , \labels[4].label[196] );
tran (\labels[4][204] , \labels[4].label[195] );
tran (\labels[4][203] , \labels[4].label[194] );
tran (\labels[4][202] , \labels[4].label[193] );
tran (\labels[4][201] , \labels[4].label[192] );
tran (\labels[4][200] , \labels[4].label[191] );
tran (\labels[4][199] , \labels[4].label[190] );
tran (\labels[4][198] , \labels[4].label[189] );
tran (\labels[4][197] , \labels[4].label[188] );
tran (\labels[4][196] , \labels[4].label[187] );
tran (\labels[4][195] , \labels[4].label[186] );
tran (\labels[4][194] , \labels[4].label[185] );
tran (\labels[4][193] , \labels[4].label[184] );
tran (\labels[4][192] , \labels[4].label[183] );
tran (\labels[4][191] , \labels[4].label[182] );
tran (\labels[4][190] , \labels[4].label[181] );
tran (\labels[4][189] , \labels[4].label[180] );
tran (\labels[4][188] , \labels[4].label[179] );
tran (\labels[4][187] , \labels[4].label[178] );
tran (\labels[4][186] , \labels[4].label[177] );
tran (\labels[4][185] , \labels[4].label[176] );
tran (\labels[4][184] , \labels[4].label[175] );
tran (\labels[4][183] , \labels[4].label[174] );
tran (\labels[4][182] , \labels[4].label[173] );
tran (\labels[4][181] , \labels[4].label[172] );
tran (\labels[4][180] , \labels[4].label[171] );
tran (\labels[4][179] , \labels[4].label[170] );
tran (\labels[4][178] , \labels[4].label[169] );
tran (\labels[4][177] , \labels[4].label[168] );
tran (\labels[4][176] , \labels[4].label[167] );
tran (\labels[4][175] , \labels[4].label[166] );
tran (\labels[4][174] , \labels[4].label[165] );
tran (\labels[4][173] , \labels[4].label[164] );
tran (\labels[4][172] , \labels[4].label[163] );
tran (\labels[4][171] , \labels[4].label[162] );
tran (\labels[4][170] , \labels[4].label[161] );
tran (\labels[4][169] , \labels[4].label[160] );
tran (\labels[4][168] , \labels[4].label[159] );
tran (\labels[4][167] , \labels[4].label[158] );
tran (\labels[4][166] , \labels[4].label[157] );
tran (\labels[4][165] , \labels[4].label[156] );
tran (\labels[4][164] , \labels[4].label[155] );
tran (\labels[4][163] , \labels[4].label[154] );
tran (\labels[4][162] , \labels[4].label[153] );
tran (\labels[4][161] , \labels[4].label[152] );
tran (\labels[4][160] , \labels[4].label[151] );
tran (\labels[4][159] , \labels[4].label[150] );
tran (\labels[4][158] , \labels[4].label[149] );
tran (\labels[4][157] , \labels[4].label[148] );
tran (\labels[4][156] , \labels[4].label[147] );
tran (\labels[4][155] , \labels[4].label[146] );
tran (\labels[4][154] , \labels[4].label[145] );
tran (\labels[4][153] , \labels[4].label[144] );
tran (\labels[4][152] , \labels[4].label[143] );
tran (\labels[4][151] , \labels[4].label[142] );
tran (\labels[4][150] , \labels[4].label[141] );
tran (\labels[4][149] , \labels[4].label[140] );
tran (\labels[4][148] , \labels[4].label[139] );
tran (\labels[4][147] , \labels[4].label[138] );
tran (\labels[4][146] , \labels[4].label[137] );
tran (\labels[4][145] , \labels[4].label[136] );
tran (\labels[4][144] , \labels[4].label[135] );
tran (\labels[4][143] , \labels[4].label[134] );
tran (\labels[4][142] , \labels[4].label[133] );
tran (\labels[4][141] , \labels[4].label[132] );
tran (\labels[4][140] , \labels[4].label[131] );
tran (\labels[4][139] , \labels[4].label[130] );
tran (\labels[4][138] , \labels[4].label[129] );
tran (\labels[4][137] , \labels[4].label[128] );
tran (\labels[4][136] , \labels[4].label[127] );
tran (\labels[4][135] , \labels[4].label[126] );
tran (\labels[4][134] , \labels[4].label[125] );
tran (\labels[4][133] , \labels[4].label[124] );
tran (\labels[4][132] , \labels[4].label[123] );
tran (\labels[4][131] , \labels[4].label[122] );
tran (\labels[4][130] , \labels[4].label[121] );
tran (\labels[4][129] , \labels[4].label[120] );
tran (\labels[4][128] , \labels[4].label[119] );
tran (\labels[4][127] , \labels[4].label[118] );
tran (\labels[4][126] , \labels[4].label[117] );
tran (\labels[4][125] , \labels[4].label[116] );
tran (\labels[4][124] , \labels[4].label[115] );
tran (\labels[4][123] , \labels[4].label[114] );
tran (\labels[4][122] , \labels[4].label[113] );
tran (\labels[4][121] , \labels[4].label[112] );
tran (\labels[4][120] , \labels[4].label[111] );
tran (\labels[4][119] , \labels[4].label[110] );
tran (\labels[4][118] , \labels[4].label[109] );
tran (\labels[4][117] , \labels[4].label[108] );
tran (\labels[4][116] , \labels[4].label[107] );
tran (\labels[4][115] , \labels[4].label[106] );
tran (\labels[4][114] , \labels[4].label[105] );
tran (\labels[4][113] , \labels[4].label[104] );
tran (\labels[4][112] , \labels[4].label[103] );
tran (\labels[4][111] , \labels[4].label[102] );
tran (\labels[4][110] , \labels[4].label[101] );
tran (\labels[4][109] , \labels[4].label[100] );
tran (\labels[4][108] , \labels[4].label[99] );
tran (\labels[4][107] , \labels[4].label[98] );
tran (\labels[4][106] , \labels[4].label[97] );
tran (\labels[4][105] , \labels[4].label[96] );
tran (\labels[4][104] , \labels[4].label[95] );
tran (\labels[4][103] , \labels[4].label[94] );
tran (\labels[4][102] , \labels[4].label[93] );
tran (\labels[4][101] , \labels[4].label[92] );
tran (\labels[4][100] , \labels[4].label[91] );
tran (\labels[4][99] , \labels[4].label[90] );
tran (\labels[4][98] , \labels[4].label[89] );
tran (\labels[4][97] , \labels[4].label[88] );
tran (\labels[4][96] , \labels[4].label[87] );
tran (\labels[4][95] , \labels[4].label[86] );
tran (\labels[4][94] , \labels[4].label[85] );
tran (\labels[4][93] , \labels[4].label[84] );
tran (\labels[4][92] , \labels[4].label[83] );
tran (\labels[4][91] , \labels[4].label[82] );
tran (\labels[4][90] , \labels[4].label[81] );
tran (\labels[4][89] , \labels[4].label[80] );
tran (\labels[4][88] , \labels[4].label[79] );
tran (\labels[4][87] , \labels[4].label[78] );
tran (\labels[4][86] , \labels[4].label[77] );
tran (\labels[4][85] , \labels[4].label[76] );
tran (\labels[4][84] , \labels[4].label[75] );
tran (\labels[4][83] , \labels[4].label[74] );
tran (\labels[4][82] , \labels[4].label[73] );
tran (\labels[4][81] , \labels[4].label[72] );
tran (\labels[4][80] , \labels[4].label[71] );
tran (\labels[4][79] , \labels[4].label[70] );
tran (\labels[4][78] , \labels[4].label[69] );
tran (\labels[4][77] , \labels[4].label[68] );
tran (\labels[4][76] , \labels[4].label[67] );
tran (\labels[4][75] , \labels[4].label[66] );
tran (\labels[4][74] , \labels[4].label[65] );
tran (\labels[4][73] , \labels[4].label[64] );
tran (\labels[4][72] , \labels[4].label[63] );
tran (\labels[4][71] , \labels[4].label[62] );
tran (\labels[4][70] , \labels[4].label[61] );
tran (\labels[4][69] , \labels[4].label[60] );
tran (\labels[4][68] , \labels[4].label[59] );
tran (\labels[4][67] , \labels[4].label[58] );
tran (\labels[4][66] , \labels[4].label[57] );
tran (\labels[4][65] , \labels[4].label[56] );
tran (\labels[4][64] , \labels[4].label[55] );
tran (\labels[4][63] , \labels[4].label[54] );
tran (\labels[4][62] , \labels[4].label[53] );
tran (\labels[4][61] , \labels[4].label[52] );
tran (\labels[4][60] , \labels[4].label[51] );
tran (\labels[4][59] , \labels[4].label[50] );
tran (\labels[4][58] , \labels[4].label[49] );
tran (\labels[4][57] , \labels[4].label[48] );
tran (\labels[4][56] , \labels[4].label[47] );
tran (\labels[4][55] , \labels[4].label[46] );
tran (\labels[4][54] , \labels[4].label[45] );
tran (\labels[4][53] , \labels[4].label[44] );
tran (\labels[4][52] , \labels[4].label[43] );
tran (\labels[4][51] , \labels[4].label[42] );
tran (\labels[4][50] , \labels[4].label[41] );
tran (\labels[4][49] , \labels[4].label[40] );
tran (\labels[4][48] , \labels[4].label[39] );
tran (\labels[4][47] , \labels[4].label[38] );
tran (\labels[4][46] , \labels[4].label[37] );
tran (\labels[4][45] , \labels[4].label[36] );
tran (\labels[4][44] , \labels[4].label[35] );
tran (\labels[4][43] , \labels[4].label[34] );
tran (\labels[4][42] , \labels[4].label[33] );
tran (\labels[4][41] , \labels[4].label[32] );
tran (\labels[4][40] , \labels[4].label[31] );
tran (\labels[4][39] , \labels[4].label[30] );
tran (\labels[4][38] , \labels[4].label[29] );
tran (\labels[4][37] , \labels[4].label[28] );
tran (\labels[4][36] , \labels[4].label[27] );
tran (\labels[4][35] , \labels[4].label[26] );
tran (\labels[4][34] , \labels[4].label[25] );
tran (\labels[4][33] , \labels[4].label[24] );
tran (\labels[4][32] , \labels[4].label[23] );
tran (\labels[4][31] , \labels[4].label[22] );
tran (\labels[4][30] , \labels[4].label[21] );
tran (\labels[4][29] , \labels[4].label[20] );
tran (\labels[4][28] , \labels[4].label[19] );
tran (\labels[4][27] , \labels[4].label[18] );
tran (\labels[4][26] , \labels[4].label[17] );
tran (\labels[4][25] , \labels[4].label[16] );
tran (\labels[4][24] , \labels[4].label[15] );
tran (\labels[4][23] , \labels[4].label[14] );
tran (\labels[4][22] , \labels[4].label[13] );
tran (\labels[4][21] , \labels[4].label[12] );
tran (\labels[4][20] , \labels[4].label[11] );
tran (\labels[4][19] , \labels[4].label[10] );
tran (\labels[4][18] , \labels[4].label[9] );
tran (\labels[4][17] , \labels[4].label[8] );
tran (\labels[4][16] , \labels[4].label[7] );
tran (\labels[4][15] , \labels[4].label[6] );
tran (\labels[4][14] , \labels[4].label[5] );
tran (\labels[4][13] , \labels[4].label[4] );
tran (\labels[4][12] , \labels[4].label[3] );
tran (\labels[4][11] , \labels[4].label[2] );
tran (\labels[4][10] , \labels[4].label[1] );
tran (\labels[4][9] , \labels[4].label[0] );
tran (\labels[4][8] , \labels[4].delimiter_valid[0] );
tran (\labels[4][7] , \labels[4].delimiter[7] );
tran (\labels[4][6] , \labels[4].delimiter[6] );
tran (\labels[4][5] , \labels[4].delimiter[5] );
tran (\labels[4][4] , \labels[4].delimiter[4] );
tran (\labels[4][3] , \labels[4].delimiter[3] );
tran (\labels[4][2] , \labels[4].delimiter[2] );
tran (\labels[4][1] , \labels[4].delimiter[1] );
tran (\labels[4][0] , \labels[4].delimiter[0] );
tran (\labels[3][271] , \labels[3].guid_size[0] );
tran (\labels[3][270] , \labels[3].label_size[5] );
tran (\labels[3][269] , \labels[3].label_size[4] );
tran (\labels[3][268] , \labels[3].label_size[3] );
tran (\labels[3][267] , \labels[3].label_size[2] );
tran (\labels[3][266] , \labels[3].label_size[1] );
tran (\labels[3][265] , \labels[3].label_size[0] );
tran (\labels[3][264] , \labels[3].label[255] );
tran (\labels[3][263] , \labels[3].label[254] );
tran (\labels[3][262] , \labels[3].label[253] );
tran (\labels[3][261] , \labels[3].label[252] );
tran (\labels[3][260] , \labels[3].label[251] );
tran (\labels[3][259] , \labels[3].label[250] );
tran (\labels[3][258] , \labels[3].label[249] );
tran (\labels[3][257] , \labels[3].label[248] );
tran (\labels[3][256] , \labels[3].label[247] );
tran (\labels[3][255] , \labels[3].label[246] );
tran (\labels[3][254] , \labels[3].label[245] );
tran (\labels[3][253] , \labels[3].label[244] );
tran (\labels[3][252] , \labels[3].label[243] );
tran (\labels[3][251] , \labels[3].label[242] );
tran (\labels[3][250] , \labels[3].label[241] );
tran (\labels[3][249] , \labels[3].label[240] );
tran (\labels[3][248] , \labels[3].label[239] );
tran (\labels[3][247] , \labels[3].label[238] );
tran (\labels[3][246] , \labels[3].label[237] );
tran (\labels[3][245] , \labels[3].label[236] );
tran (\labels[3][244] , \labels[3].label[235] );
tran (\labels[3][243] , \labels[3].label[234] );
tran (\labels[3][242] , \labels[3].label[233] );
tran (\labels[3][241] , \labels[3].label[232] );
tran (\labels[3][240] , \labels[3].label[231] );
tran (\labels[3][239] , \labels[3].label[230] );
tran (\labels[3][238] , \labels[3].label[229] );
tran (\labels[3][237] , \labels[3].label[228] );
tran (\labels[3][236] , \labels[3].label[227] );
tran (\labels[3][235] , \labels[3].label[226] );
tran (\labels[3][234] , \labels[3].label[225] );
tran (\labels[3][233] , \labels[3].label[224] );
tran (\labels[3][232] , \labels[3].label[223] );
tran (\labels[3][231] , \labels[3].label[222] );
tran (\labels[3][230] , \labels[3].label[221] );
tran (\labels[3][229] , \labels[3].label[220] );
tran (\labels[3][228] , \labels[3].label[219] );
tran (\labels[3][227] , \labels[3].label[218] );
tran (\labels[3][226] , \labels[3].label[217] );
tran (\labels[3][225] , \labels[3].label[216] );
tran (\labels[3][224] , \labels[3].label[215] );
tran (\labels[3][223] , \labels[3].label[214] );
tran (\labels[3][222] , \labels[3].label[213] );
tran (\labels[3][221] , \labels[3].label[212] );
tran (\labels[3][220] , \labels[3].label[211] );
tran (\labels[3][219] , \labels[3].label[210] );
tran (\labels[3][218] , \labels[3].label[209] );
tran (\labels[3][217] , \labels[3].label[208] );
tran (\labels[3][216] , \labels[3].label[207] );
tran (\labels[3][215] , \labels[3].label[206] );
tran (\labels[3][214] , \labels[3].label[205] );
tran (\labels[3][213] , \labels[3].label[204] );
tran (\labels[3][212] , \labels[3].label[203] );
tran (\labels[3][211] , \labels[3].label[202] );
tran (\labels[3][210] , \labels[3].label[201] );
tran (\labels[3][209] , \labels[3].label[200] );
tran (\labels[3][208] , \labels[3].label[199] );
tran (\labels[3][207] , \labels[3].label[198] );
tran (\labels[3][206] , \labels[3].label[197] );
tran (\labels[3][205] , \labels[3].label[196] );
tran (\labels[3][204] , \labels[3].label[195] );
tran (\labels[3][203] , \labels[3].label[194] );
tran (\labels[3][202] , \labels[3].label[193] );
tran (\labels[3][201] , \labels[3].label[192] );
tran (\labels[3][200] , \labels[3].label[191] );
tran (\labels[3][199] , \labels[3].label[190] );
tran (\labels[3][198] , \labels[3].label[189] );
tran (\labels[3][197] , \labels[3].label[188] );
tran (\labels[3][196] , \labels[3].label[187] );
tran (\labels[3][195] , \labels[3].label[186] );
tran (\labels[3][194] , \labels[3].label[185] );
tran (\labels[3][193] , \labels[3].label[184] );
tran (\labels[3][192] , \labels[3].label[183] );
tran (\labels[3][191] , \labels[3].label[182] );
tran (\labels[3][190] , \labels[3].label[181] );
tran (\labels[3][189] , \labels[3].label[180] );
tran (\labels[3][188] , \labels[3].label[179] );
tran (\labels[3][187] , \labels[3].label[178] );
tran (\labels[3][186] , \labels[3].label[177] );
tran (\labels[3][185] , \labels[3].label[176] );
tran (\labels[3][184] , \labels[3].label[175] );
tran (\labels[3][183] , \labels[3].label[174] );
tran (\labels[3][182] , \labels[3].label[173] );
tran (\labels[3][181] , \labels[3].label[172] );
tran (\labels[3][180] , \labels[3].label[171] );
tran (\labels[3][179] , \labels[3].label[170] );
tran (\labels[3][178] , \labels[3].label[169] );
tran (\labels[3][177] , \labels[3].label[168] );
tran (\labels[3][176] , \labels[3].label[167] );
tran (\labels[3][175] , \labels[3].label[166] );
tran (\labels[3][174] , \labels[3].label[165] );
tran (\labels[3][173] , \labels[3].label[164] );
tran (\labels[3][172] , \labels[3].label[163] );
tran (\labels[3][171] , \labels[3].label[162] );
tran (\labels[3][170] , \labels[3].label[161] );
tran (\labels[3][169] , \labels[3].label[160] );
tran (\labels[3][168] , \labels[3].label[159] );
tran (\labels[3][167] , \labels[3].label[158] );
tran (\labels[3][166] , \labels[3].label[157] );
tran (\labels[3][165] , \labels[3].label[156] );
tran (\labels[3][164] , \labels[3].label[155] );
tran (\labels[3][163] , \labels[3].label[154] );
tran (\labels[3][162] , \labels[3].label[153] );
tran (\labels[3][161] , \labels[3].label[152] );
tran (\labels[3][160] , \labels[3].label[151] );
tran (\labels[3][159] , \labels[3].label[150] );
tran (\labels[3][158] , \labels[3].label[149] );
tran (\labels[3][157] , \labels[3].label[148] );
tran (\labels[3][156] , \labels[3].label[147] );
tran (\labels[3][155] , \labels[3].label[146] );
tran (\labels[3][154] , \labels[3].label[145] );
tran (\labels[3][153] , \labels[3].label[144] );
tran (\labels[3][152] , \labels[3].label[143] );
tran (\labels[3][151] , \labels[3].label[142] );
tran (\labels[3][150] , \labels[3].label[141] );
tran (\labels[3][149] , \labels[3].label[140] );
tran (\labels[3][148] , \labels[3].label[139] );
tran (\labels[3][147] , \labels[3].label[138] );
tran (\labels[3][146] , \labels[3].label[137] );
tran (\labels[3][145] , \labels[3].label[136] );
tran (\labels[3][144] , \labels[3].label[135] );
tran (\labels[3][143] , \labels[3].label[134] );
tran (\labels[3][142] , \labels[3].label[133] );
tran (\labels[3][141] , \labels[3].label[132] );
tran (\labels[3][140] , \labels[3].label[131] );
tran (\labels[3][139] , \labels[3].label[130] );
tran (\labels[3][138] , \labels[3].label[129] );
tran (\labels[3][137] , \labels[3].label[128] );
tran (\labels[3][136] , \labels[3].label[127] );
tran (\labels[3][135] , \labels[3].label[126] );
tran (\labels[3][134] , \labels[3].label[125] );
tran (\labels[3][133] , \labels[3].label[124] );
tran (\labels[3][132] , \labels[3].label[123] );
tran (\labels[3][131] , \labels[3].label[122] );
tran (\labels[3][130] , \labels[3].label[121] );
tran (\labels[3][129] , \labels[3].label[120] );
tran (\labels[3][128] , \labels[3].label[119] );
tran (\labels[3][127] , \labels[3].label[118] );
tran (\labels[3][126] , \labels[3].label[117] );
tran (\labels[3][125] , \labels[3].label[116] );
tran (\labels[3][124] , \labels[3].label[115] );
tran (\labels[3][123] , \labels[3].label[114] );
tran (\labels[3][122] , \labels[3].label[113] );
tran (\labels[3][121] , \labels[3].label[112] );
tran (\labels[3][120] , \labels[3].label[111] );
tran (\labels[3][119] , \labels[3].label[110] );
tran (\labels[3][118] , \labels[3].label[109] );
tran (\labels[3][117] , \labels[3].label[108] );
tran (\labels[3][116] , \labels[3].label[107] );
tran (\labels[3][115] , \labels[3].label[106] );
tran (\labels[3][114] , \labels[3].label[105] );
tran (\labels[3][113] , \labels[3].label[104] );
tran (\labels[3][112] , \labels[3].label[103] );
tran (\labels[3][111] , \labels[3].label[102] );
tran (\labels[3][110] , \labels[3].label[101] );
tran (\labels[3][109] , \labels[3].label[100] );
tran (\labels[3][108] , \labels[3].label[99] );
tran (\labels[3][107] , \labels[3].label[98] );
tran (\labels[3][106] , \labels[3].label[97] );
tran (\labels[3][105] , \labels[3].label[96] );
tran (\labels[3][104] , \labels[3].label[95] );
tran (\labels[3][103] , \labels[3].label[94] );
tran (\labels[3][102] , \labels[3].label[93] );
tran (\labels[3][101] , \labels[3].label[92] );
tran (\labels[3][100] , \labels[3].label[91] );
tran (\labels[3][99] , \labels[3].label[90] );
tran (\labels[3][98] , \labels[3].label[89] );
tran (\labels[3][97] , \labels[3].label[88] );
tran (\labels[3][96] , \labels[3].label[87] );
tran (\labels[3][95] , \labels[3].label[86] );
tran (\labels[3][94] , \labels[3].label[85] );
tran (\labels[3][93] , \labels[3].label[84] );
tran (\labels[3][92] , \labels[3].label[83] );
tran (\labels[3][91] , \labels[3].label[82] );
tran (\labels[3][90] , \labels[3].label[81] );
tran (\labels[3][89] , \labels[3].label[80] );
tran (\labels[3][88] , \labels[3].label[79] );
tran (\labels[3][87] , \labels[3].label[78] );
tran (\labels[3][86] , \labels[3].label[77] );
tran (\labels[3][85] , \labels[3].label[76] );
tran (\labels[3][84] , \labels[3].label[75] );
tran (\labels[3][83] , \labels[3].label[74] );
tran (\labels[3][82] , \labels[3].label[73] );
tran (\labels[3][81] , \labels[3].label[72] );
tran (\labels[3][80] , \labels[3].label[71] );
tran (\labels[3][79] , \labels[3].label[70] );
tran (\labels[3][78] , \labels[3].label[69] );
tran (\labels[3][77] , \labels[3].label[68] );
tran (\labels[3][76] , \labels[3].label[67] );
tran (\labels[3][75] , \labels[3].label[66] );
tran (\labels[3][74] , \labels[3].label[65] );
tran (\labels[3][73] , \labels[3].label[64] );
tran (\labels[3][72] , \labels[3].label[63] );
tran (\labels[3][71] , \labels[3].label[62] );
tran (\labels[3][70] , \labels[3].label[61] );
tran (\labels[3][69] , \labels[3].label[60] );
tran (\labels[3][68] , \labels[3].label[59] );
tran (\labels[3][67] , \labels[3].label[58] );
tran (\labels[3][66] , \labels[3].label[57] );
tran (\labels[3][65] , \labels[3].label[56] );
tran (\labels[3][64] , \labels[3].label[55] );
tran (\labels[3][63] , \labels[3].label[54] );
tran (\labels[3][62] , \labels[3].label[53] );
tran (\labels[3][61] , \labels[3].label[52] );
tran (\labels[3][60] , \labels[3].label[51] );
tran (\labels[3][59] , \labels[3].label[50] );
tran (\labels[3][58] , \labels[3].label[49] );
tran (\labels[3][57] , \labels[3].label[48] );
tran (\labels[3][56] , \labels[3].label[47] );
tran (\labels[3][55] , \labels[3].label[46] );
tran (\labels[3][54] , \labels[3].label[45] );
tran (\labels[3][53] , \labels[3].label[44] );
tran (\labels[3][52] , \labels[3].label[43] );
tran (\labels[3][51] , \labels[3].label[42] );
tran (\labels[3][50] , \labels[3].label[41] );
tran (\labels[3][49] , \labels[3].label[40] );
tran (\labels[3][48] , \labels[3].label[39] );
tran (\labels[3][47] , \labels[3].label[38] );
tran (\labels[3][46] , \labels[3].label[37] );
tran (\labels[3][45] , \labels[3].label[36] );
tran (\labels[3][44] , \labels[3].label[35] );
tran (\labels[3][43] , \labels[3].label[34] );
tran (\labels[3][42] , \labels[3].label[33] );
tran (\labels[3][41] , \labels[3].label[32] );
tran (\labels[3][40] , \labels[3].label[31] );
tran (\labels[3][39] , \labels[3].label[30] );
tran (\labels[3][38] , \labels[3].label[29] );
tran (\labels[3][37] , \labels[3].label[28] );
tran (\labels[3][36] , \labels[3].label[27] );
tran (\labels[3][35] , \labels[3].label[26] );
tran (\labels[3][34] , \labels[3].label[25] );
tran (\labels[3][33] , \labels[3].label[24] );
tran (\labels[3][32] , \labels[3].label[23] );
tran (\labels[3][31] , \labels[3].label[22] );
tran (\labels[3][30] , \labels[3].label[21] );
tran (\labels[3][29] , \labels[3].label[20] );
tran (\labels[3][28] , \labels[3].label[19] );
tran (\labels[3][27] , \labels[3].label[18] );
tran (\labels[3][26] , \labels[3].label[17] );
tran (\labels[3][25] , \labels[3].label[16] );
tran (\labels[3][24] , \labels[3].label[15] );
tran (\labels[3][23] , \labels[3].label[14] );
tran (\labels[3][22] , \labels[3].label[13] );
tran (\labels[3][21] , \labels[3].label[12] );
tran (\labels[3][20] , \labels[3].label[11] );
tran (\labels[3][19] , \labels[3].label[10] );
tran (\labels[3][18] , \labels[3].label[9] );
tran (\labels[3][17] , \labels[3].label[8] );
tran (\labels[3][16] , \labels[3].label[7] );
tran (\labels[3][15] , \labels[3].label[6] );
tran (\labels[3][14] , \labels[3].label[5] );
tran (\labels[3][13] , \labels[3].label[4] );
tran (\labels[3][12] , \labels[3].label[3] );
tran (\labels[3][11] , \labels[3].label[2] );
tran (\labels[3][10] , \labels[3].label[1] );
tran (\labels[3][9] , \labels[3].label[0] );
tran (\labels[3][8] , \labels[3].delimiter_valid[0] );
tran (\labels[3][7] , \labels[3].delimiter[7] );
tran (\labels[3][6] , \labels[3].delimiter[6] );
tran (\labels[3][5] , \labels[3].delimiter[5] );
tran (\labels[3][4] , \labels[3].delimiter[4] );
tran (\labels[3][3] , \labels[3].delimiter[3] );
tran (\labels[3][2] , \labels[3].delimiter[2] );
tran (\labels[3][1] , \labels[3].delimiter[1] );
tran (\labels[3][0] , \labels[3].delimiter[0] );
tran (\labels[2][271] , \labels[2].guid_size[0] );
tran (\labels[2][270] , \labels[2].label_size[5] );
tran (\labels[2][269] , \labels[2].label_size[4] );
tran (\labels[2][268] , \labels[2].label_size[3] );
tran (\labels[2][267] , \labels[2].label_size[2] );
tran (\labels[2][266] , \labels[2].label_size[1] );
tran (\labels[2][265] , \labels[2].label_size[0] );
tran (\labels[2][264] , \labels[2].label[255] );
tran (\labels[2][263] , \labels[2].label[254] );
tran (\labels[2][262] , \labels[2].label[253] );
tran (\labels[2][261] , \labels[2].label[252] );
tran (\labels[2][260] , \labels[2].label[251] );
tran (\labels[2][259] , \labels[2].label[250] );
tran (\labels[2][258] , \labels[2].label[249] );
tran (\labels[2][257] , \labels[2].label[248] );
tran (\labels[2][256] , \labels[2].label[247] );
tran (\labels[2][255] , \labels[2].label[246] );
tran (\labels[2][254] , \labels[2].label[245] );
tran (\labels[2][253] , \labels[2].label[244] );
tran (\labels[2][252] , \labels[2].label[243] );
tran (\labels[2][251] , \labels[2].label[242] );
tran (\labels[2][250] , \labels[2].label[241] );
tran (\labels[2][249] , \labels[2].label[240] );
tran (\labels[2][248] , \labels[2].label[239] );
tran (\labels[2][247] , \labels[2].label[238] );
tran (\labels[2][246] , \labels[2].label[237] );
tran (\labels[2][245] , \labels[2].label[236] );
tran (\labels[2][244] , \labels[2].label[235] );
tran (\labels[2][243] , \labels[2].label[234] );
tran (\labels[2][242] , \labels[2].label[233] );
tran (\labels[2][241] , \labels[2].label[232] );
tran (\labels[2][240] , \labels[2].label[231] );
tran (\labels[2][239] , \labels[2].label[230] );
tran (\labels[2][238] , \labels[2].label[229] );
tran (\labels[2][237] , \labels[2].label[228] );
tran (\labels[2][236] , \labels[2].label[227] );
tran (\labels[2][235] , \labels[2].label[226] );
tran (\labels[2][234] , \labels[2].label[225] );
tran (\labels[2][233] , \labels[2].label[224] );
tran (\labels[2][232] , \labels[2].label[223] );
tran (\labels[2][231] , \labels[2].label[222] );
tran (\labels[2][230] , \labels[2].label[221] );
tran (\labels[2][229] , \labels[2].label[220] );
tran (\labels[2][228] , \labels[2].label[219] );
tran (\labels[2][227] , \labels[2].label[218] );
tran (\labels[2][226] , \labels[2].label[217] );
tran (\labels[2][225] , \labels[2].label[216] );
tran (\labels[2][224] , \labels[2].label[215] );
tran (\labels[2][223] , \labels[2].label[214] );
tran (\labels[2][222] , \labels[2].label[213] );
tran (\labels[2][221] , \labels[2].label[212] );
tran (\labels[2][220] , \labels[2].label[211] );
tran (\labels[2][219] , \labels[2].label[210] );
tran (\labels[2][218] , \labels[2].label[209] );
tran (\labels[2][217] , \labels[2].label[208] );
tran (\labels[2][216] , \labels[2].label[207] );
tran (\labels[2][215] , \labels[2].label[206] );
tran (\labels[2][214] , \labels[2].label[205] );
tran (\labels[2][213] , \labels[2].label[204] );
tran (\labels[2][212] , \labels[2].label[203] );
tran (\labels[2][211] , \labels[2].label[202] );
tran (\labels[2][210] , \labels[2].label[201] );
tran (\labels[2][209] , \labels[2].label[200] );
tran (\labels[2][208] , \labels[2].label[199] );
tran (\labels[2][207] , \labels[2].label[198] );
tran (\labels[2][206] , \labels[2].label[197] );
tran (\labels[2][205] , \labels[2].label[196] );
tran (\labels[2][204] , \labels[2].label[195] );
tran (\labels[2][203] , \labels[2].label[194] );
tran (\labels[2][202] , \labels[2].label[193] );
tran (\labels[2][201] , \labels[2].label[192] );
tran (\labels[2][200] , \labels[2].label[191] );
tran (\labels[2][199] , \labels[2].label[190] );
tran (\labels[2][198] , \labels[2].label[189] );
tran (\labels[2][197] , \labels[2].label[188] );
tran (\labels[2][196] , \labels[2].label[187] );
tran (\labels[2][195] , \labels[2].label[186] );
tran (\labels[2][194] , \labels[2].label[185] );
tran (\labels[2][193] , \labels[2].label[184] );
tran (\labels[2][192] , \labels[2].label[183] );
tran (\labels[2][191] , \labels[2].label[182] );
tran (\labels[2][190] , \labels[2].label[181] );
tran (\labels[2][189] , \labels[2].label[180] );
tran (\labels[2][188] , \labels[2].label[179] );
tran (\labels[2][187] , \labels[2].label[178] );
tran (\labels[2][186] , \labels[2].label[177] );
tran (\labels[2][185] , \labels[2].label[176] );
tran (\labels[2][184] , \labels[2].label[175] );
tran (\labels[2][183] , \labels[2].label[174] );
tran (\labels[2][182] , \labels[2].label[173] );
tran (\labels[2][181] , \labels[2].label[172] );
tran (\labels[2][180] , \labels[2].label[171] );
tran (\labels[2][179] , \labels[2].label[170] );
tran (\labels[2][178] , \labels[2].label[169] );
tran (\labels[2][177] , \labels[2].label[168] );
tran (\labels[2][176] , \labels[2].label[167] );
tran (\labels[2][175] , \labels[2].label[166] );
tran (\labels[2][174] , \labels[2].label[165] );
tran (\labels[2][173] , \labels[2].label[164] );
tran (\labels[2][172] , \labels[2].label[163] );
tran (\labels[2][171] , \labels[2].label[162] );
tran (\labels[2][170] , \labels[2].label[161] );
tran (\labels[2][169] , \labels[2].label[160] );
tran (\labels[2][168] , \labels[2].label[159] );
tran (\labels[2][167] , \labels[2].label[158] );
tran (\labels[2][166] , \labels[2].label[157] );
tran (\labels[2][165] , \labels[2].label[156] );
tran (\labels[2][164] , \labels[2].label[155] );
tran (\labels[2][163] , \labels[2].label[154] );
tran (\labels[2][162] , \labels[2].label[153] );
tran (\labels[2][161] , \labels[2].label[152] );
tran (\labels[2][160] , \labels[2].label[151] );
tran (\labels[2][159] , \labels[2].label[150] );
tran (\labels[2][158] , \labels[2].label[149] );
tran (\labels[2][157] , \labels[2].label[148] );
tran (\labels[2][156] , \labels[2].label[147] );
tran (\labels[2][155] , \labels[2].label[146] );
tran (\labels[2][154] , \labels[2].label[145] );
tran (\labels[2][153] , \labels[2].label[144] );
tran (\labels[2][152] , \labels[2].label[143] );
tran (\labels[2][151] , \labels[2].label[142] );
tran (\labels[2][150] , \labels[2].label[141] );
tran (\labels[2][149] , \labels[2].label[140] );
tran (\labels[2][148] , \labels[2].label[139] );
tran (\labels[2][147] , \labels[2].label[138] );
tran (\labels[2][146] , \labels[2].label[137] );
tran (\labels[2][145] , \labels[2].label[136] );
tran (\labels[2][144] , \labels[2].label[135] );
tran (\labels[2][143] , \labels[2].label[134] );
tran (\labels[2][142] , \labels[2].label[133] );
tran (\labels[2][141] , \labels[2].label[132] );
tran (\labels[2][140] , \labels[2].label[131] );
tran (\labels[2][139] , \labels[2].label[130] );
tran (\labels[2][138] , \labels[2].label[129] );
tran (\labels[2][137] , \labels[2].label[128] );
tran (\labels[2][136] , \labels[2].label[127] );
tran (\labels[2][135] , \labels[2].label[126] );
tran (\labels[2][134] , \labels[2].label[125] );
tran (\labels[2][133] , \labels[2].label[124] );
tran (\labels[2][132] , \labels[2].label[123] );
tran (\labels[2][131] , \labels[2].label[122] );
tran (\labels[2][130] , \labels[2].label[121] );
tran (\labels[2][129] , \labels[2].label[120] );
tran (\labels[2][128] , \labels[2].label[119] );
tran (\labels[2][127] , \labels[2].label[118] );
tran (\labels[2][126] , \labels[2].label[117] );
tran (\labels[2][125] , \labels[2].label[116] );
tran (\labels[2][124] , \labels[2].label[115] );
tran (\labels[2][123] , \labels[2].label[114] );
tran (\labels[2][122] , \labels[2].label[113] );
tran (\labels[2][121] , \labels[2].label[112] );
tran (\labels[2][120] , \labels[2].label[111] );
tran (\labels[2][119] , \labels[2].label[110] );
tran (\labels[2][118] , \labels[2].label[109] );
tran (\labels[2][117] , \labels[2].label[108] );
tran (\labels[2][116] , \labels[2].label[107] );
tran (\labels[2][115] , \labels[2].label[106] );
tran (\labels[2][114] , \labels[2].label[105] );
tran (\labels[2][113] , \labels[2].label[104] );
tran (\labels[2][112] , \labels[2].label[103] );
tran (\labels[2][111] , \labels[2].label[102] );
tran (\labels[2][110] , \labels[2].label[101] );
tran (\labels[2][109] , \labels[2].label[100] );
tran (\labels[2][108] , \labels[2].label[99] );
tran (\labels[2][107] , \labels[2].label[98] );
tran (\labels[2][106] , \labels[2].label[97] );
tran (\labels[2][105] , \labels[2].label[96] );
tran (\labels[2][104] , \labels[2].label[95] );
tran (\labels[2][103] , \labels[2].label[94] );
tran (\labels[2][102] , \labels[2].label[93] );
tran (\labels[2][101] , \labels[2].label[92] );
tran (\labels[2][100] , \labels[2].label[91] );
tran (\labels[2][99] , \labels[2].label[90] );
tran (\labels[2][98] , \labels[2].label[89] );
tran (\labels[2][97] , \labels[2].label[88] );
tran (\labels[2][96] , \labels[2].label[87] );
tran (\labels[2][95] , \labels[2].label[86] );
tran (\labels[2][94] , \labels[2].label[85] );
tran (\labels[2][93] , \labels[2].label[84] );
tran (\labels[2][92] , \labels[2].label[83] );
tran (\labels[2][91] , \labels[2].label[82] );
tran (\labels[2][90] , \labels[2].label[81] );
tran (\labels[2][89] , \labels[2].label[80] );
tran (\labels[2][88] , \labels[2].label[79] );
tran (\labels[2][87] , \labels[2].label[78] );
tran (\labels[2][86] , \labels[2].label[77] );
tran (\labels[2][85] , \labels[2].label[76] );
tran (\labels[2][84] , \labels[2].label[75] );
tran (\labels[2][83] , \labels[2].label[74] );
tran (\labels[2][82] , \labels[2].label[73] );
tran (\labels[2][81] , \labels[2].label[72] );
tran (\labels[2][80] , \labels[2].label[71] );
tran (\labels[2][79] , \labels[2].label[70] );
tran (\labels[2][78] , \labels[2].label[69] );
tran (\labels[2][77] , \labels[2].label[68] );
tran (\labels[2][76] , \labels[2].label[67] );
tran (\labels[2][75] , \labels[2].label[66] );
tran (\labels[2][74] , \labels[2].label[65] );
tran (\labels[2][73] , \labels[2].label[64] );
tran (\labels[2][72] , \labels[2].label[63] );
tran (\labels[2][71] , \labels[2].label[62] );
tran (\labels[2][70] , \labels[2].label[61] );
tran (\labels[2][69] , \labels[2].label[60] );
tran (\labels[2][68] , \labels[2].label[59] );
tran (\labels[2][67] , \labels[2].label[58] );
tran (\labels[2][66] , \labels[2].label[57] );
tran (\labels[2][65] , \labels[2].label[56] );
tran (\labels[2][64] , \labels[2].label[55] );
tran (\labels[2][63] , \labels[2].label[54] );
tran (\labels[2][62] , \labels[2].label[53] );
tran (\labels[2][61] , \labels[2].label[52] );
tran (\labels[2][60] , \labels[2].label[51] );
tran (\labels[2][59] , \labels[2].label[50] );
tran (\labels[2][58] , \labels[2].label[49] );
tran (\labels[2][57] , \labels[2].label[48] );
tran (\labels[2][56] , \labels[2].label[47] );
tran (\labels[2][55] , \labels[2].label[46] );
tran (\labels[2][54] , \labels[2].label[45] );
tran (\labels[2][53] , \labels[2].label[44] );
tran (\labels[2][52] , \labels[2].label[43] );
tran (\labels[2][51] , \labels[2].label[42] );
tran (\labels[2][50] , \labels[2].label[41] );
tran (\labels[2][49] , \labels[2].label[40] );
tran (\labels[2][48] , \labels[2].label[39] );
tran (\labels[2][47] , \labels[2].label[38] );
tran (\labels[2][46] , \labels[2].label[37] );
tran (\labels[2][45] , \labels[2].label[36] );
tran (\labels[2][44] , \labels[2].label[35] );
tran (\labels[2][43] , \labels[2].label[34] );
tran (\labels[2][42] , \labels[2].label[33] );
tran (\labels[2][41] , \labels[2].label[32] );
tran (\labels[2][40] , \labels[2].label[31] );
tran (\labels[2][39] , \labels[2].label[30] );
tran (\labels[2][38] , \labels[2].label[29] );
tran (\labels[2][37] , \labels[2].label[28] );
tran (\labels[2][36] , \labels[2].label[27] );
tran (\labels[2][35] , \labels[2].label[26] );
tran (\labels[2][34] , \labels[2].label[25] );
tran (\labels[2][33] , \labels[2].label[24] );
tran (\labels[2][32] , \labels[2].label[23] );
tran (\labels[2][31] , \labels[2].label[22] );
tran (\labels[2][30] , \labels[2].label[21] );
tran (\labels[2][29] , \labels[2].label[20] );
tran (\labels[2][28] , \labels[2].label[19] );
tran (\labels[2][27] , \labels[2].label[18] );
tran (\labels[2][26] , \labels[2].label[17] );
tran (\labels[2][25] , \labels[2].label[16] );
tran (\labels[2][24] , \labels[2].label[15] );
tran (\labels[2][23] , \labels[2].label[14] );
tran (\labels[2][22] , \labels[2].label[13] );
tran (\labels[2][21] , \labels[2].label[12] );
tran (\labels[2][20] , \labels[2].label[11] );
tran (\labels[2][19] , \labels[2].label[10] );
tran (\labels[2][18] , \labels[2].label[9] );
tran (\labels[2][17] , \labels[2].label[8] );
tran (\labels[2][16] , \labels[2].label[7] );
tran (\labels[2][15] , \labels[2].label[6] );
tran (\labels[2][14] , \labels[2].label[5] );
tran (\labels[2][13] , \labels[2].label[4] );
tran (\labels[2][12] , \labels[2].label[3] );
tran (\labels[2][11] , \labels[2].label[2] );
tran (\labels[2][10] , \labels[2].label[1] );
tran (\labels[2][9] , \labels[2].label[0] );
tran (\labels[2][8] , \labels[2].delimiter_valid[0] );
tran (\labels[2][7] , \labels[2].delimiter[7] );
tran (\labels[2][6] , \labels[2].delimiter[6] );
tran (\labels[2][5] , \labels[2].delimiter[5] );
tran (\labels[2][4] , \labels[2].delimiter[4] );
tran (\labels[2][3] , \labels[2].delimiter[3] );
tran (\labels[2][2] , \labels[2].delimiter[2] );
tran (\labels[2][1] , \labels[2].delimiter[1] );
tran (\labels[2][0] , \labels[2].delimiter[0] );
tran (\labels[1][271] , \labels[1].guid_size[0] );
tran (\labels[1][270] , \labels[1].label_size[5] );
tran (\labels[1][269] , \labels[1].label_size[4] );
tran (\labels[1][268] , \labels[1].label_size[3] );
tran (\labels[1][267] , \labels[1].label_size[2] );
tran (\labels[1][266] , \labels[1].label_size[1] );
tran (\labels[1][265] , \labels[1].label_size[0] );
tran (\labels[1][264] , \labels[1].label[255] );
tran (\labels[1][263] , \labels[1].label[254] );
tran (\labels[1][262] , \labels[1].label[253] );
tran (\labels[1][261] , \labels[1].label[252] );
tran (\labels[1][260] , \labels[1].label[251] );
tran (\labels[1][259] , \labels[1].label[250] );
tran (\labels[1][258] , \labels[1].label[249] );
tran (\labels[1][257] , \labels[1].label[248] );
tran (\labels[1][256] , \labels[1].label[247] );
tran (\labels[1][255] , \labels[1].label[246] );
tran (\labels[1][254] , \labels[1].label[245] );
tran (\labels[1][253] , \labels[1].label[244] );
tran (\labels[1][252] , \labels[1].label[243] );
tran (\labels[1][251] , \labels[1].label[242] );
tran (\labels[1][250] , \labels[1].label[241] );
tran (\labels[1][249] , \labels[1].label[240] );
tran (\labels[1][248] , \labels[1].label[239] );
tran (\labels[1][247] , \labels[1].label[238] );
tran (\labels[1][246] , \labels[1].label[237] );
tran (\labels[1][245] , \labels[1].label[236] );
tran (\labels[1][244] , \labels[1].label[235] );
tran (\labels[1][243] , \labels[1].label[234] );
tran (\labels[1][242] , \labels[1].label[233] );
tran (\labels[1][241] , \labels[1].label[232] );
tran (\labels[1][240] , \labels[1].label[231] );
tran (\labels[1][239] , \labels[1].label[230] );
tran (\labels[1][238] , \labels[1].label[229] );
tran (\labels[1][237] , \labels[1].label[228] );
tran (\labels[1][236] , \labels[1].label[227] );
tran (\labels[1][235] , \labels[1].label[226] );
tran (\labels[1][234] , \labels[1].label[225] );
tran (\labels[1][233] , \labels[1].label[224] );
tran (\labels[1][232] , \labels[1].label[223] );
tran (\labels[1][231] , \labels[1].label[222] );
tran (\labels[1][230] , \labels[1].label[221] );
tran (\labels[1][229] , \labels[1].label[220] );
tran (\labels[1][228] , \labels[1].label[219] );
tran (\labels[1][227] , \labels[1].label[218] );
tran (\labels[1][226] , \labels[1].label[217] );
tran (\labels[1][225] , \labels[1].label[216] );
tran (\labels[1][224] , \labels[1].label[215] );
tran (\labels[1][223] , \labels[1].label[214] );
tran (\labels[1][222] , \labels[1].label[213] );
tran (\labels[1][221] , \labels[1].label[212] );
tran (\labels[1][220] , \labels[1].label[211] );
tran (\labels[1][219] , \labels[1].label[210] );
tran (\labels[1][218] , \labels[1].label[209] );
tran (\labels[1][217] , \labels[1].label[208] );
tran (\labels[1][216] , \labels[1].label[207] );
tran (\labels[1][215] , \labels[1].label[206] );
tran (\labels[1][214] , \labels[1].label[205] );
tran (\labels[1][213] , \labels[1].label[204] );
tran (\labels[1][212] , \labels[1].label[203] );
tran (\labels[1][211] , \labels[1].label[202] );
tran (\labels[1][210] , \labels[1].label[201] );
tran (\labels[1][209] , \labels[1].label[200] );
tran (\labels[1][208] , \labels[1].label[199] );
tran (\labels[1][207] , \labels[1].label[198] );
tran (\labels[1][206] , \labels[1].label[197] );
tran (\labels[1][205] , \labels[1].label[196] );
tran (\labels[1][204] , \labels[1].label[195] );
tran (\labels[1][203] , \labels[1].label[194] );
tran (\labels[1][202] , \labels[1].label[193] );
tran (\labels[1][201] , \labels[1].label[192] );
tran (\labels[1][200] , \labels[1].label[191] );
tran (\labels[1][199] , \labels[1].label[190] );
tran (\labels[1][198] , \labels[1].label[189] );
tran (\labels[1][197] , \labels[1].label[188] );
tran (\labels[1][196] , \labels[1].label[187] );
tran (\labels[1][195] , \labels[1].label[186] );
tran (\labels[1][194] , \labels[1].label[185] );
tran (\labels[1][193] , \labels[1].label[184] );
tran (\labels[1][192] , \labels[1].label[183] );
tran (\labels[1][191] , \labels[1].label[182] );
tran (\labels[1][190] , \labels[1].label[181] );
tran (\labels[1][189] , \labels[1].label[180] );
tran (\labels[1][188] , \labels[1].label[179] );
tran (\labels[1][187] , \labels[1].label[178] );
tran (\labels[1][186] , \labels[1].label[177] );
tran (\labels[1][185] , \labels[1].label[176] );
tran (\labels[1][184] , \labels[1].label[175] );
tran (\labels[1][183] , \labels[1].label[174] );
tran (\labels[1][182] , \labels[1].label[173] );
tran (\labels[1][181] , \labels[1].label[172] );
tran (\labels[1][180] , \labels[1].label[171] );
tran (\labels[1][179] , \labels[1].label[170] );
tran (\labels[1][178] , \labels[1].label[169] );
tran (\labels[1][177] , \labels[1].label[168] );
tran (\labels[1][176] , \labels[1].label[167] );
tran (\labels[1][175] , \labels[1].label[166] );
tran (\labels[1][174] , \labels[1].label[165] );
tran (\labels[1][173] , \labels[1].label[164] );
tran (\labels[1][172] , \labels[1].label[163] );
tran (\labels[1][171] , \labels[1].label[162] );
tran (\labels[1][170] , \labels[1].label[161] );
tran (\labels[1][169] , \labels[1].label[160] );
tran (\labels[1][168] , \labels[1].label[159] );
tran (\labels[1][167] , \labels[1].label[158] );
tran (\labels[1][166] , \labels[1].label[157] );
tran (\labels[1][165] , \labels[1].label[156] );
tran (\labels[1][164] , \labels[1].label[155] );
tran (\labels[1][163] , \labels[1].label[154] );
tran (\labels[1][162] , \labels[1].label[153] );
tran (\labels[1][161] , \labels[1].label[152] );
tran (\labels[1][160] , \labels[1].label[151] );
tran (\labels[1][159] , \labels[1].label[150] );
tran (\labels[1][158] , \labels[1].label[149] );
tran (\labels[1][157] , \labels[1].label[148] );
tran (\labels[1][156] , \labels[1].label[147] );
tran (\labels[1][155] , \labels[1].label[146] );
tran (\labels[1][154] , \labels[1].label[145] );
tran (\labels[1][153] , \labels[1].label[144] );
tran (\labels[1][152] , \labels[1].label[143] );
tran (\labels[1][151] , \labels[1].label[142] );
tran (\labels[1][150] , \labels[1].label[141] );
tran (\labels[1][149] , \labels[1].label[140] );
tran (\labels[1][148] , \labels[1].label[139] );
tran (\labels[1][147] , \labels[1].label[138] );
tran (\labels[1][146] , \labels[1].label[137] );
tran (\labels[1][145] , \labels[1].label[136] );
tran (\labels[1][144] , \labels[1].label[135] );
tran (\labels[1][143] , \labels[1].label[134] );
tran (\labels[1][142] , \labels[1].label[133] );
tran (\labels[1][141] , \labels[1].label[132] );
tran (\labels[1][140] , \labels[1].label[131] );
tran (\labels[1][139] , \labels[1].label[130] );
tran (\labels[1][138] , \labels[1].label[129] );
tran (\labels[1][137] , \labels[1].label[128] );
tran (\labels[1][136] , \labels[1].label[127] );
tran (\labels[1][135] , \labels[1].label[126] );
tran (\labels[1][134] , \labels[1].label[125] );
tran (\labels[1][133] , \labels[1].label[124] );
tran (\labels[1][132] , \labels[1].label[123] );
tran (\labels[1][131] , \labels[1].label[122] );
tran (\labels[1][130] , \labels[1].label[121] );
tran (\labels[1][129] , \labels[1].label[120] );
tran (\labels[1][128] , \labels[1].label[119] );
tran (\labels[1][127] , \labels[1].label[118] );
tran (\labels[1][126] , \labels[1].label[117] );
tran (\labels[1][125] , \labels[1].label[116] );
tran (\labels[1][124] , \labels[1].label[115] );
tran (\labels[1][123] , \labels[1].label[114] );
tran (\labels[1][122] , \labels[1].label[113] );
tran (\labels[1][121] , \labels[1].label[112] );
tran (\labels[1][120] , \labels[1].label[111] );
tran (\labels[1][119] , \labels[1].label[110] );
tran (\labels[1][118] , \labels[1].label[109] );
tran (\labels[1][117] , \labels[1].label[108] );
tran (\labels[1][116] , \labels[1].label[107] );
tran (\labels[1][115] , \labels[1].label[106] );
tran (\labels[1][114] , \labels[1].label[105] );
tran (\labels[1][113] , \labels[1].label[104] );
tran (\labels[1][112] , \labels[1].label[103] );
tran (\labels[1][111] , \labels[1].label[102] );
tran (\labels[1][110] , \labels[1].label[101] );
tran (\labels[1][109] , \labels[1].label[100] );
tran (\labels[1][108] , \labels[1].label[99] );
tran (\labels[1][107] , \labels[1].label[98] );
tran (\labels[1][106] , \labels[1].label[97] );
tran (\labels[1][105] , \labels[1].label[96] );
tran (\labels[1][104] , \labels[1].label[95] );
tran (\labels[1][103] , \labels[1].label[94] );
tran (\labels[1][102] , \labels[1].label[93] );
tran (\labels[1][101] , \labels[1].label[92] );
tran (\labels[1][100] , \labels[1].label[91] );
tran (\labels[1][99] , \labels[1].label[90] );
tran (\labels[1][98] , \labels[1].label[89] );
tran (\labels[1][97] , \labels[1].label[88] );
tran (\labels[1][96] , \labels[1].label[87] );
tran (\labels[1][95] , \labels[1].label[86] );
tran (\labels[1][94] , \labels[1].label[85] );
tran (\labels[1][93] , \labels[1].label[84] );
tran (\labels[1][92] , \labels[1].label[83] );
tran (\labels[1][91] , \labels[1].label[82] );
tran (\labels[1][90] , \labels[1].label[81] );
tran (\labels[1][89] , \labels[1].label[80] );
tran (\labels[1][88] , \labels[1].label[79] );
tran (\labels[1][87] , \labels[1].label[78] );
tran (\labels[1][86] , \labels[1].label[77] );
tran (\labels[1][85] , \labels[1].label[76] );
tran (\labels[1][84] , \labels[1].label[75] );
tran (\labels[1][83] , \labels[1].label[74] );
tran (\labels[1][82] , \labels[1].label[73] );
tran (\labels[1][81] , \labels[1].label[72] );
tran (\labels[1][80] , \labels[1].label[71] );
tran (\labels[1][79] , \labels[1].label[70] );
tran (\labels[1][78] , \labels[1].label[69] );
tran (\labels[1][77] , \labels[1].label[68] );
tran (\labels[1][76] , \labels[1].label[67] );
tran (\labels[1][75] , \labels[1].label[66] );
tran (\labels[1][74] , \labels[1].label[65] );
tran (\labels[1][73] , \labels[1].label[64] );
tran (\labels[1][72] , \labels[1].label[63] );
tran (\labels[1][71] , \labels[1].label[62] );
tran (\labels[1][70] , \labels[1].label[61] );
tran (\labels[1][69] , \labels[1].label[60] );
tran (\labels[1][68] , \labels[1].label[59] );
tran (\labels[1][67] , \labels[1].label[58] );
tran (\labels[1][66] , \labels[1].label[57] );
tran (\labels[1][65] , \labels[1].label[56] );
tran (\labels[1][64] , \labels[1].label[55] );
tran (\labels[1][63] , \labels[1].label[54] );
tran (\labels[1][62] , \labels[1].label[53] );
tran (\labels[1][61] , \labels[1].label[52] );
tran (\labels[1][60] , \labels[1].label[51] );
tran (\labels[1][59] , \labels[1].label[50] );
tran (\labels[1][58] , \labels[1].label[49] );
tran (\labels[1][57] , \labels[1].label[48] );
tran (\labels[1][56] , \labels[1].label[47] );
tran (\labels[1][55] , \labels[1].label[46] );
tran (\labels[1][54] , \labels[1].label[45] );
tran (\labels[1][53] , \labels[1].label[44] );
tran (\labels[1][52] , \labels[1].label[43] );
tran (\labels[1][51] , \labels[1].label[42] );
tran (\labels[1][50] , \labels[1].label[41] );
tran (\labels[1][49] , \labels[1].label[40] );
tran (\labels[1][48] , \labels[1].label[39] );
tran (\labels[1][47] , \labels[1].label[38] );
tran (\labels[1][46] , \labels[1].label[37] );
tran (\labels[1][45] , \labels[1].label[36] );
tran (\labels[1][44] , \labels[1].label[35] );
tran (\labels[1][43] , \labels[1].label[34] );
tran (\labels[1][42] , \labels[1].label[33] );
tran (\labels[1][41] , \labels[1].label[32] );
tran (\labels[1][40] , \labels[1].label[31] );
tran (\labels[1][39] , \labels[1].label[30] );
tran (\labels[1][38] , \labels[1].label[29] );
tran (\labels[1][37] , \labels[1].label[28] );
tran (\labels[1][36] , \labels[1].label[27] );
tran (\labels[1][35] , \labels[1].label[26] );
tran (\labels[1][34] , \labels[1].label[25] );
tran (\labels[1][33] , \labels[1].label[24] );
tran (\labels[1][32] , \labels[1].label[23] );
tran (\labels[1][31] , \labels[1].label[22] );
tran (\labels[1][30] , \labels[1].label[21] );
tran (\labels[1][29] , \labels[1].label[20] );
tran (\labels[1][28] , \labels[1].label[19] );
tran (\labels[1][27] , \labels[1].label[18] );
tran (\labels[1][26] , \labels[1].label[17] );
tran (\labels[1][25] , \labels[1].label[16] );
tran (\labels[1][24] , \labels[1].label[15] );
tran (\labels[1][23] , \labels[1].label[14] );
tran (\labels[1][22] , \labels[1].label[13] );
tran (\labels[1][21] , \labels[1].label[12] );
tran (\labels[1][20] , \labels[1].label[11] );
tran (\labels[1][19] , \labels[1].label[10] );
tran (\labels[1][18] , \labels[1].label[9] );
tran (\labels[1][17] , \labels[1].label[8] );
tran (\labels[1][16] , \labels[1].label[7] );
tran (\labels[1][15] , \labels[1].label[6] );
tran (\labels[1][14] , \labels[1].label[5] );
tran (\labels[1][13] , \labels[1].label[4] );
tran (\labels[1][12] , \labels[1].label[3] );
tran (\labels[1][11] , \labels[1].label[2] );
tran (\labels[1][10] , \labels[1].label[1] );
tran (\labels[1][9] , \labels[1].label[0] );
tran (\labels[1][8] , \labels[1].delimiter_valid[0] );
tran (\labels[1][7] , \labels[1].delimiter[7] );
tran (\labels[1][6] , \labels[1].delimiter[6] );
tran (\labels[1][5] , \labels[1].delimiter[5] );
tran (\labels[1][4] , \labels[1].delimiter[4] );
tran (\labels[1][3] , \labels[1].delimiter[3] );
tran (\labels[1][2] , \labels[1].delimiter[2] );
tran (\labels[1][1] , \labels[1].delimiter[1] );
tran (\labels[1][0] , \labels[1].delimiter[0] );
tran (\labels[0][271] , \labels[0].guid_size[0] );
tran (\labels[0][270] , \labels[0].label_size[5] );
tran (\labels[0][269] , \labels[0].label_size[4] );
tran (\labels[0][268] , \labels[0].label_size[3] );
tran (\labels[0][267] , \labels[0].label_size[2] );
tran (\labels[0][266] , \labels[0].label_size[1] );
tran (\labels[0][265] , \labels[0].label_size[0] );
tran (\labels[0][264] , \labels[0].label[255] );
tran (\labels[0][263] , \labels[0].label[254] );
tran (\labels[0][262] , \labels[0].label[253] );
tran (\labels[0][261] , \labels[0].label[252] );
tran (\labels[0][260] , \labels[0].label[251] );
tran (\labels[0][259] , \labels[0].label[250] );
tran (\labels[0][258] , \labels[0].label[249] );
tran (\labels[0][257] , \labels[0].label[248] );
tran (\labels[0][256] , \labels[0].label[247] );
tran (\labels[0][255] , \labels[0].label[246] );
tran (\labels[0][254] , \labels[0].label[245] );
tran (\labels[0][253] , \labels[0].label[244] );
tran (\labels[0][252] , \labels[0].label[243] );
tran (\labels[0][251] , \labels[0].label[242] );
tran (\labels[0][250] , \labels[0].label[241] );
tran (\labels[0][249] , \labels[0].label[240] );
tran (\labels[0][248] , \labels[0].label[239] );
tran (\labels[0][247] , \labels[0].label[238] );
tran (\labels[0][246] , \labels[0].label[237] );
tran (\labels[0][245] , \labels[0].label[236] );
tran (\labels[0][244] , \labels[0].label[235] );
tran (\labels[0][243] , \labels[0].label[234] );
tran (\labels[0][242] , \labels[0].label[233] );
tran (\labels[0][241] , \labels[0].label[232] );
tran (\labels[0][240] , \labels[0].label[231] );
tran (\labels[0][239] , \labels[0].label[230] );
tran (\labels[0][238] , \labels[0].label[229] );
tran (\labels[0][237] , \labels[0].label[228] );
tran (\labels[0][236] , \labels[0].label[227] );
tran (\labels[0][235] , \labels[0].label[226] );
tran (\labels[0][234] , \labels[0].label[225] );
tran (\labels[0][233] , \labels[0].label[224] );
tran (\labels[0][232] , \labels[0].label[223] );
tran (\labels[0][231] , \labels[0].label[222] );
tran (\labels[0][230] , \labels[0].label[221] );
tran (\labels[0][229] , \labels[0].label[220] );
tran (\labels[0][228] , \labels[0].label[219] );
tran (\labels[0][227] , \labels[0].label[218] );
tran (\labels[0][226] , \labels[0].label[217] );
tran (\labels[0][225] , \labels[0].label[216] );
tran (\labels[0][224] , \labels[0].label[215] );
tran (\labels[0][223] , \labels[0].label[214] );
tran (\labels[0][222] , \labels[0].label[213] );
tran (\labels[0][221] , \labels[0].label[212] );
tran (\labels[0][220] , \labels[0].label[211] );
tran (\labels[0][219] , \labels[0].label[210] );
tran (\labels[0][218] , \labels[0].label[209] );
tran (\labels[0][217] , \labels[0].label[208] );
tran (\labels[0][216] , \labels[0].label[207] );
tran (\labels[0][215] , \labels[0].label[206] );
tran (\labels[0][214] , \labels[0].label[205] );
tran (\labels[0][213] , \labels[0].label[204] );
tran (\labels[0][212] , \labels[0].label[203] );
tran (\labels[0][211] , \labels[0].label[202] );
tran (\labels[0][210] , \labels[0].label[201] );
tran (\labels[0][209] , \labels[0].label[200] );
tran (\labels[0][208] , \labels[0].label[199] );
tran (\labels[0][207] , \labels[0].label[198] );
tran (\labels[0][206] , \labels[0].label[197] );
tran (\labels[0][205] , \labels[0].label[196] );
tran (\labels[0][204] , \labels[0].label[195] );
tran (\labels[0][203] , \labels[0].label[194] );
tran (\labels[0][202] , \labels[0].label[193] );
tran (\labels[0][201] , \labels[0].label[192] );
tran (\labels[0][200] , \labels[0].label[191] );
tran (\labels[0][199] , \labels[0].label[190] );
tran (\labels[0][198] , \labels[0].label[189] );
tran (\labels[0][197] , \labels[0].label[188] );
tran (\labels[0][196] , \labels[0].label[187] );
tran (\labels[0][195] , \labels[0].label[186] );
tran (\labels[0][194] , \labels[0].label[185] );
tran (\labels[0][193] , \labels[0].label[184] );
tran (\labels[0][192] , \labels[0].label[183] );
tran (\labels[0][191] , \labels[0].label[182] );
tran (\labels[0][190] , \labels[0].label[181] );
tran (\labels[0][189] , \labels[0].label[180] );
tran (\labels[0][188] , \labels[0].label[179] );
tran (\labels[0][187] , \labels[0].label[178] );
tran (\labels[0][186] , \labels[0].label[177] );
tran (\labels[0][185] , \labels[0].label[176] );
tran (\labels[0][184] , \labels[0].label[175] );
tran (\labels[0][183] , \labels[0].label[174] );
tran (\labels[0][182] , \labels[0].label[173] );
tran (\labels[0][181] , \labels[0].label[172] );
tran (\labels[0][180] , \labels[0].label[171] );
tran (\labels[0][179] , \labels[0].label[170] );
tran (\labels[0][178] , \labels[0].label[169] );
tran (\labels[0][177] , \labels[0].label[168] );
tran (\labels[0][176] , \labels[0].label[167] );
tran (\labels[0][175] , \labels[0].label[166] );
tran (\labels[0][174] , \labels[0].label[165] );
tran (\labels[0][173] , \labels[0].label[164] );
tran (\labels[0][172] , \labels[0].label[163] );
tran (\labels[0][171] , \labels[0].label[162] );
tran (\labels[0][170] , \labels[0].label[161] );
tran (\labels[0][169] , \labels[0].label[160] );
tran (\labels[0][168] , \labels[0].label[159] );
tran (\labels[0][167] , \labels[0].label[158] );
tran (\labels[0][166] , \labels[0].label[157] );
tran (\labels[0][165] , \labels[0].label[156] );
tran (\labels[0][164] , \labels[0].label[155] );
tran (\labels[0][163] , \labels[0].label[154] );
tran (\labels[0][162] , \labels[0].label[153] );
tran (\labels[0][161] , \labels[0].label[152] );
tran (\labels[0][160] , \labels[0].label[151] );
tran (\labels[0][159] , \labels[0].label[150] );
tran (\labels[0][158] , \labels[0].label[149] );
tran (\labels[0][157] , \labels[0].label[148] );
tran (\labels[0][156] , \labels[0].label[147] );
tran (\labels[0][155] , \labels[0].label[146] );
tran (\labels[0][154] , \labels[0].label[145] );
tran (\labels[0][153] , \labels[0].label[144] );
tran (\labels[0][152] , \labels[0].label[143] );
tran (\labels[0][151] , \labels[0].label[142] );
tran (\labels[0][150] , \labels[0].label[141] );
tran (\labels[0][149] , \labels[0].label[140] );
tran (\labels[0][148] , \labels[0].label[139] );
tran (\labels[0][147] , \labels[0].label[138] );
tran (\labels[0][146] , \labels[0].label[137] );
tran (\labels[0][145] , \labels[0].label[136] );
tran (\labels[0][144] , \labels[0].label[135] );
tran (\labels[0][143] , \labels[0].label[134] );
tran (\labels[0][142] , \labels[0].label[133] );
tran (\labels[0][141] , \labels[0].label[132] );
tran (\labels[0][140] , \labels[0].label[131] );
tran (\labels[0][139] , \labels[0].label[130] );
tran (\labels[0][138] , \labels[0].label[129] );
tran (\labels[0][137] , \labels[0].label[128] );
tran (\labels[0][136] , \labels[0].label[127] );
tran (\labels[0][135] , \labels[0].label[126] );
tran (\labels[0][134] , \labels[0].label[125] );
tran (\labels[0][133] , \labels[0].label[124] );
tran (\labels[0][132] , \labels[0].label[123] );
tran (\labels[0][131] , \labels[0].label[122] );
tran (\labels[0][130] , \labels[0].label[121] );
tran (\labels[0][129] , \labels[0].label[120] );
tran (\labels[0][128] , \labels[0].label[119] );
tran (\labels[0][127] , \labels[0].label[118] );
tran (\labels[0][126] , \labels[0].label[117] );
tran (\labels[0][125] , \labels[0].label[116] );
tran (\labels[0][124] , \labels[0].label[115] );
tran (\labels[0][123] , \labels[0].label[114] );
tran (\labels[0][122] , \labels[0].label[113] );
tran (\labels[0][121] , \labels[0].label[112] );
tran (\labels[0][120] , \labels[0].label[111] );
tran (\labels[0][119] , \labels[0].label[110] );
tran (\labels[0][118] , \labels[0].label[109] );
tran (\labels[0][117] , \labels[0].label[108] );
tran (\labels[0][116] , \labels[0].label[107] );
tran (\labels[0][115] , \labels[0].label[106] );
tran (\labels[0][114] , \labels[0].label[105] );
tran (\labels[0][113] , \labels[0].label[104] );
tran (\labels[0][112] , \labels[0].label[103] );
tran (\labels[0][111] , \labels[0].label[102] );
tran (\labels[0][110] , \labels[0].label[101] );
tran (\labels[0][109] , \labels[0].label[100] );
tran (\labels[0][108] , \labels[0].label[99] );
tran (\labels[0][107] , \labels[0].label[98] );
tran (\labels[0][106] , \labels[0].label[97] );
tran (\labels[0][105] , \labels[0].label[96] );
tran (\labels[0][104] , \labels[0].label[95] );
tran (\labels[0][103] , \labels[0].label[94] );
tran (\labels[0][102] , \labels[0].label[93] );
tran (\labels[0][101] , \labels[0].label[92] );
tran (\labels[0][100] , \labels[0].label[91] );
tran (\labels[0][99] , \labels[0].label[90] );
tran (\labels[0][98] , \labels[0].label[89] );
tran (\labels[0][97] , \labels[0].label[88] );
tran (\labels[0][96] , \labels[0].label[87] );
tran (\labels[0][95] , \labels[0].label[86] );
tran (\labels[0][94] , \labels[0].label[85] );
tran (\labels[0][93] , \labels[0].label[84] );
tran (\labels[0][92] , \labels[0].label[83] );
tran (\labels[0][91] , \labels[0].label[82] );
tran (\labels[0][90] , \labels[0].label[81] );
tran (\labels[0][89] , \labels[0].label[80] );
tran (\labels[0][88] , \labels[0].label[79] );
tran (\labels[0][87] , \labels[0].label[78] );
tran (\labels[0][86] , \labels[0].label[77] );
tran (\labels[0][85] , \labels[0].label[76] );
tran (\labels[0][84] , \labels[0].label[75] );
tran (\labels[0][83] , \labels[0].label[74] );
tran (\labels[0][82] , \labels[0].label[73] );
tran (\labels[0][81] , \labels[0].label[72] );
tran (\labels[0][80] , \labels[0].label[71] );
tran (\labels[0][79] , \labels[0].label[70] );
tran (\labels[0][78] , \labels[0].label[69] );
tran (\labels[0][77] , \labels[0].label[68] );
tran (\labels[0][76] , \labels[0].label[67] );
tran (\labels[0][75] , \labels[0].label[66] );
tran (\labels[0][74] , \labels[0].label[65] );
tran (\labels[0][73] , \labels[0].label[64] );
tran (\labels[0][72] , \labels[0].label[63] );
tran (\labels[0][71] , \labels[0].label[62] );
tran (\labels[0][70] , \labels[0].label[61] );
tran (\labels[0][69] , \labels[0].label[60] );
tran (\labels[0][68] , \labels[0].label[59] );
tran (\labels[0][67] , \labels[0].label[58] );
tran (\labels[0][66] , \labels[0].label[57] );
tran (\labels[0][65] , \labels[0].label[56] );
tran (\labels[0][64] , \labels[0].label[55] );
tran (\labels[0][63] , \labels[0].label[54] );
tran (\labels[0][62] , \labels[0].label[53] );
tran (\labels[0][61] , \labels[0].label[52] );
tran (\labels[0][60] , \labels[0].label[51] );
tran (\labels[0][59] , \labels[0].label[50] );
tran (\labels[0][58] , \labels[0].label[49] );
tran (\labels[0][57] , \labels[0].label[48] );
tran (\labels[0][56] , \labels[0].label[47] );
tran (\labels[0][55] , \labels[0].label[46] );
tran (\labels[0][54] , \labels[0].label[45] );
tran (\labels[0][53] , \labels[0].label[44] );
tran (\labels[0][52] , \labels[0].label[43] );
tran (\labels[0][51] , \labels[0].label[42] );
tran (\labels[0][50] , \labels[0].label[41] );
tran (\labels[0][49] , \labels[0].label[40] );
tran (\labels[0][48] , \labels[0].label[39] );
tran (\labels[0][47] , \labels[0].label[38] );
tran (\labels[0][46] , \labels[0].label[37] );
tran (\labels[0][45] , \labels[0].label[36] );
tran (\labels[0][44] , \labels[0].label[35] );
tran (\labels[0][43] , \labels[0].label[34] );
tran (\labels[0][42] , \labels[0].label[33] );
tran (\labels[0][41] , \labels[0].label[32] );
tran (\labels[0][40] , \labels[0].label[31] );
tran (\labels[0][39] , \labels[0].label[30] );
tran (\labels[0][38] , \labels[0].label[29] );
tran (\labels[0][37] , \labels[0].label[28] );
tran (\labels[0][36] , \labels[0].label[27] );
tran (\labels[0][35] , \labels[0].label[26] );
tran (\labels[0][34] , \labels[0].label[25] );
tran (\labels[0][33] , \labels[0].label[24] );
tran (\labels[0][32] , \labels[0].label[23] );
tran (\labels[0][31] , \labels[0].label[22] );
tran (\labels[0][30] , \labels[0].label[21] );
tran (\labels[0][29] , \labels[0].label[20] );
tran (\labels[0][28] , \labels[0].label[19] );
tran (\labels[0][27] , \labels[0].label[18] );
tran (\labels[0][26] , \labels[0].label[17] );
tran (\labels[0][25] , \labels[0].label[16] );
tran (\labels[0][24] , \labels[0].label[15] );
tran (\labels[0][23] , \labels[0].label[14] );
tran (\labels[0][22] , \labels[0].label[13] );
tran (\labels[0][21] , \labels[0].label[12] );
tran (\labels[0][20] , \labels[0].label[11] );
tran (\labels[0][19] , \labels[0].label[10] );
tran (\labels[0][18] , \labels[0].label[9] );
tran (\labels[0][17] , \labels[0].label[8] );
tran (\labels[0][16] , \labels[0].label[7] );
tran (\labels[0][15] , \labels[0].label[6] );
tran (\labels[0][14] , \labels[0].label[5] );
tran (\labels[0][13] , \labels[0].label[4] );
tran (\labels[0][12] , \labels[0].label[3] );
tran (\labels[0][11] , \labels[0].label[2] );
tran (\labels[0][10] , \labels[0].label[1] );
tran (\labels[0][9] , \labels[0].label[0] );
tran (\labels[0][8] , \labels[0].delimiter_valid[0] );
tran (\labels[0][7] , \labels[0].delimiter[7] );
tran (\labels[0][6] , \labels[0].delimiter[6] );
tran (\labels[0][5] , \labels[0].delimiter[5] );
tran (\labels[0][4] , \labels[0].delimiter[4] );
tran (\labels[0][3] , \labels[0].delimiter[3] );
tran (\labels[0][2] , \labels[0].delimiter[2] );
tran (\labels[0][1] , \labels[0].delimiter[1] );
tran (\labels[0][0] , \labels[0].delimiter[0] );
tran (tready_override[8], \tready_override.r.part0 [8]);
tran (tready_override[8], \tready_override.f.txc_tready_override );
tran (tready_override[7], \tready_override.r.part0 [7]);
tran (tready_override[7], \tready_override.f.engine_7_tready_override );
tran (tready_override[6], \tready_override.r.part0 [6]);
tran (tready_override[6], \tready_override.f.engine_6_tready_override );
tran (tready_override[5], \tready_override.r.part0 [5]);
tran (tready_override[5], \tready_override.f.engine_5_tready_override );
tran (tready_override[4], \tready_override.r.part0 [4]);
tran (tready_override[4], \tready_override.f.engine_4_tready_override );
tran (tready_override[3], \tready_override.r.part0 [3]);
tran (tready_override[3], \tready_override.f.engine_3_tready_override );
tran (tready_override[2], \tready_override.r.part0 [2]);
tran (tready_override[2], \tready_override.f.engine_2_tready_override );
tran (tready_override[1], \tready_override.r.part0 [1]);
tran (tready_override[1], \tready_override.f.engine_1_tready_override );
tran (tready_override[0], \tready_override.r.part0 [0]);
tran (tready_override[0], \tready_override.f.engine_0_tready_override );
tran (cceip_encrypt_kop_fifo_override[6], \cceip_encrypt_kop_fifo_override.r.part0 [6]);
tran (cceip_encrypt_kop_fifo_override[6], \cceip_encrypt_kop_fifo_override.f.gcm_status_data_fifo );
tran (cceip_encrypt_kop_fifo_override[5], \cceip_encrypt_kop_fifo_override.r.part0 [5]);
tran (cceip_encrypt_kop_fifo_override[5], \cceip_encrypt_kop_fifo_override.f.tlv_sb_data_fifo );
tran (cceip_encrypt_kop_fifo_override[4], \cceip_encrypt_kop_fifo_override.r.part0 [4]);
tran (cceip_encrypt_kop_fifo_override[4], \cceip_encrypt_kop_fifo_override.f.kdf_cmd_fifo );
tran (cceip_encrypt_kop_fifo_override[3], \cceip_encrypt_kop_fifo_override.r.part0 [3]);
tran (cceip_encrypt_kop_fifo_override[3], \cceip_encrypt_kop_fifo_override.f.kdfstream_cmd_fifo );
tran (cceip_encrypt_kop_fifo_override[2], \cceip_encrypt_kop_fifo_override.r.part0 [2]);
tran (cceip_encrypt_kop_fifo_override[2], \cceip_encrypt_kop_fifo_override.f.keyfilter_cmd_fifo );
tran (cceip_encrypt_kop_fifo_override[1], \cceip_encrypt_kop_fifo_override.r.part0 [1]);
tran (cceip_encrypt_kop_fifo_override[1], \cceip_encrypt_kop_fifo_override.f.gcm_tag_data_fifo );
tran (cceip_encrypt_kop_fifo_override[0], \cceip_encrypt_kop_fifo_override.r.part0 [0]);
tran (cceip_encrypt_kop_fifo_override[0], \cceip_encrypt_kop_fifo_override.f.gcm_cmd_fifo );
tran (cceip_validate_kop_fifo_override[6], \cceip_validate_kop_fifo_override.r.part0 [6]);
tran (cceip_validate_kop_fifo_override[6], \cceip_validate_kop_fifo_override.f.gcm_status_data_fifo );
tran (cceip_validate_kop_fifo_override[5], \cceip_validate_kop_fifo_override.r.part0 [5]);
tran (cceip_validate_kop_fifo_override[5], \cceip_validate_kop_fifo_override.f.tlv_sb_data_fifo );
tran (cceip_validate_kop_fifo_override[4], \cceip_validate_kop_fifo_override.r.part0 [4]);
tran (cceip_validate_kop_fifo_override[4], \cceip_validate_kop_fifo_override.f.kdf_cmd_fifo );
tran (cceip_validate_kop_fifo_override[3], \cceip_validate_kop_fifo_override.r.part0 [3]);
tran (cceip_validate_kop_fifo_override[3], \cceip_validate_kop_fifo_override.f.kdfstream_cmd_fifo );
tran (cceip_validate_kop_fifo_override[2], \cceip_validate_kop_fifo_override.r.part0 [2]);
tran (cceip_validate_kop_fifo_override[2], \cceip_validate_kop_fifo_override.f.keyfilter_cmd_fifo );
tran (cceip_validate_kop_fifo_override[1], \cceip_validate_kop_fifo_override.r.part0 [1]);
tran (cceip_validate_kop_fifo_override[1], \cceip_validate_kop_fifo_override.f.gcm_tag_data_fifo );
tran (cceip_validate_kop_fifo_override[0], \cceip_validate_kop_fifo_override.r.part0 [0]);
tran (cceip_validate_kop_fifo_override[0], \cceip_validate_kop_fifo_override.f.gcm_cmd_fifo );
tran (cddip_decrypt_kop_fifo_override[6], \cddip_decrypt_kop_fifo_override.r.part0 [6]);
tran (cddip_decrypt_kop_fifo_override[6], \cddip_decrypt_kop_fifo_override.f.gcm_status_data_fifo );
tran (cddip_decrypt_kop_fifo_override[5], \cddip_decrypt_kop_fifo_override.r.part0 [5]);
tran (cddip_decrypt_kop_fifo_override[5], \cddip_decrypt_kop_fifo_override.f.tlv_sb_data_fifo );
tran (cddip_decrypt_kop_fifo_override[4], \cddip_decrypt_kop_fifo_override.r.part0 [4]);
tran (cddip_decrypt_kop_fifo_override[4], \cddip_decrypt_kop_fifo_override.f.kdf_cmd_fifo );
tran (cddip_decrypt_kop_fifo_override[3], \cddip_decrypt_kop_fifo_override.r.part0 [3]);
tran (cddip_decrypt_kop_fifo_override[3], \cddip_decrypt_kop_fifo_override.f.kdfstream_cmd_fifo );
tran (cddip_decrypt_kop_fifo_override[2], \cddip_decrypt_kop_fifo_override.r.part0 [2]);
tran (cddip_decrypt_kop_fifo_override[2], \cddip_decrypt_kop_fifo_override.f.keyfilter_cmd_fifo );
tran (cddip_decrypt_kop_fifo_override[1], \cddip_decrypt_kop_fifo_override.r.part0 [1]);
tran (cddip_decrypt_kop_fifo_override[1], \cddip_decrypt_kop_fifo_override.f.gcm_tag_data_fifo );
tran (cddip_decrypt_kop_fifo_override[0], \cddip_decrypt_kop_fifo_override.r.part0 [0]);
tran (cddip_decrypt_kop_fifo_override[0], \cddip_decrypt_kop_fifo_override.f.gcm_cmd_fifo );
tran (sa_global_ctrl[31], \sa_global_ctrl.r.part0 [31]);
tran (sa_global_ctrl[31], \sa_global_ctrl.f.spare [29]);
tran (sa_global_ctrl[30], \sa_global_ctrl.r.part0 [30]);
tran (sa_global_ctrl[30], \sa_global_ctrl.f.spare [28]);
tran (sa_global_ctrl[29], \sa_global_ctrl.r.part0 [29]);
tran (sa_global_ctrl[29], \sa_global_ctrl.f.spare [27]);
tran (sa_global_ctrl[28], \sa_global_ctrl.r.part0 [28]);
tran (sa_global_ctrl[28], \sa_global_ctrl.f.spare [26]);
tran (sa_global_ctrl[27], \sa_global_ctrl.r.part0 [27]);
tran (sa_global_ctrl[27], \sa_global_ctrl.f.spare [25]);
tran (sa_global_ctrl[26], \sa_global_ctrl.r.part0 [26]);
tran (sa_global_ctrl[26], \sa_global_ctrl.f.spare [24]);
tran (sa_global_ctrl[25], \sa_global_ctrl.r.part0 [25]);
tran (sa_global_ctrl[25], \sa_global_ctrl.f.spare [23]);
tran (sa_global_ctrl[24], \sa_global_ctrl.r.part0 [24]);
tran (sa_global_ctrl[24], \sa_global_ctrl.f.spare [22]);
tran (sa_global_ctrl[23], \sa_global_ctrl.r.part0 [23]);
tran (sa_global_ctrl[23], \sa_global_ctrl.f.spare [21]);
tran (sa_global_ctrl[22], \sa_global_ctrl.r.part0 [22]);
tran (sa_global_ctrl[22], \sa_global_ctrl.f.spare [20]);
tran (sa_global_ctrl[21], \sa_global_ctrl.r.part0 [21]);
tran (sa_global_ctrl[21], \sa_global_ctrl.f.spare [19]);
tran (sa_global_ctrl[20], \sa_global_ctrl.r.part0 [20]);
tran (sa_global_ctrl[20], \sa_global_ctrl.f.spare [18]);
tran (sa_global_ctrl[19], \sa_global_ctrl.r.part0 [19]);
tran (sa_global_ctrl[19], \sa_global_ctrl.f.spare [17]);
tran (sa_global_ctrl[18], \sa_global_ctrl.r.part0 [18]);
tran (sa_global_ctrl[18], \sa_global_ctrl.f.spare [16]);
tran (sa_global_ctrl[17], \sa_global_ctrl.r.part0 [17]);
tran (sa_global_ctrl[17], \sa_global_ctrl.f.spare [15]);
tran (sa_global_ctrl[16], \sa_global_ctrl.r.part0 [16]);
tran (sa_global_ctrl[16], \sa_global_ctrl.f.spare [14]);
tran (sa_global_ctrl[15], \sa_global_ctrl.r.part0 [15]);
tran (sa_global_ctrl[15], \sa_global_ctrl.f.spare [13]);
tran (sa_global_ctrl[14], \sa_global_ctrl.r.part0 [14]);
tran (sa_global_ctrl[14], \sa_global_ctrl.f.spare [12]);
tran (sa_global_ctrl[13], \sa_global_ctrl.r.part0 [13]);
tran (sa_global_ctrl[13], \sa_global_ctrl.f.spare [11]);
tran (sa_global_ctrl[12], \sa_global_ctrl.r.part0 [12]);
tran (sa_global_ctrl[12], \sa_global_ctrl.f.spare [10]);
tran (sa_global_ctrl[11], \sa_global_ctrl.r.part0 [11]);
tran (sa_global_ctrl[11], \sa_global_ctrl.f.spare [9]);
tran (sa_global_ctrl[10], \sa_global_ctrl.r.part0 [10]);
tran (sa_global_ctrl[10], \sa_global_ctrl.f.spare [8]);
tran (sa_global_ctrl[9], \sa_global_ctrl.r.part0 [9]);
tran (sa_global_ctrl[9], \sa_global_ctrl.f.spare [7]);
tran (sa_global_ctrl[8], \sa_global_ctrl.r.part0 [8]);
tran (sa_global_ctrl[8], \sa_global_ctrl.f.spare [6]);
tran (sa_global_ctrl[7], \sa_global_ctrl.r.part0 [7]);
tran (sa_global_ctrl[7], \sa_global_ctrl.f.spare [5]);
tran (sa_global_ctrl[6], \sa_global_ctrl.r.part0 [6]);
tran (sa_global_ctrl[6], \sa_global_ctrl.f.spare [4]);
tran (sa_global_ctrl[5], \sa_global_ctrl.r.part0 [5]);
tran (sa_global_ctrl[5], \sa_global_ctrl.f.spare [3]);
tran (sa_global_ctrl[4], \sa_global_ctrl.r.part0 [4]);
tran (sa_global_ctrl[4], \sa_global_ctrl.f.spare [2]);
tran (sa_global_ctrl[3], \sa_global_ctrl.r.part0 [3]);
tran (sa_global_ctrl[3], \sa_global_ctrl.f.spare [1]);
tran (sa_global_ctrl[2], \sa_global_ctrl.r.part0 [2]);
tran (sa_global_ctrl[2], \sa_global_ctrl.f.spare [0]);
tran (sa_global_ctrl[1], \sa_global_ctrl.r.part0 [1]);
tran (sa_global_ctrl[1], \sa_global_ctrl.f.sa_snap );
tran (sa_global_ctrl[0], \sa_global_ctrl.r.part0 [0]);
tran (sa_global_ctrl[0], \sa_global_ctrl.f.sa_clear_live );
tran (kme_cceip1_ob_in[0], \kme_cceip1_ob_in.tready );
tran (kme_cceip2_ob_in[0], \kme_cceip2_ob_in.tready );
tran (kme_cceip3_ob_in[0], \kme_cceip3_ob_in.tready );
tran (kme_cddip0_ob_in[0], \kme_cddip0_ob_in.tready );
tran (kme_cddip1_ob_in[0], \kme_cddip1_ob_in.tready );
tran (kme_cddip2_ob_in[0], \kme_cddip2_ob_in.tready );
tran (kme_cddip3_ob_in[0], \kme_cddip3_ob_in.tready );
tran (rbus_ring_i[1], \rbus_ring_i.ack );
tran (rbus_ring_i[0], \rbus_ring_i.err_ack );
tran (rbus_ring_i[33], \rbus_ring_i.rd_data [31]);
tran (rbus_ring_i[32], \rbus_ring_i.rd_data [30]);
tran (rbus_ring_i[31], \rbus_ring_i.rd_data [29]);
tran (rbus_ring_i[30], \rbus_ring_i.rd_data [28]);
tran (rbus_ring_i[29], \rbus_ring_i.rd_data [27]);
tran (rbus_ring_i[28], \rbus_ring_i.rd_data [26]);
tran (rbus_ring_i[27], \rbus_ring_i.rd_data [25]);
tran (rbus_ring_i[26], \rbus_ring_i.rd_data [24]);
tran (rbus_ring_i[25], \rbus_ring_i.rd_data [23]);
tran (rbus_ring_i[24], \rbus_ring_i.rd_data [22]);
tran (rbus_ring_i[23], \rbus_ring_i.rd_data [21]);
tran (rbus_ring_i[22], \rbus_ring_i.rd_data [20]);
tran (rbus_ring_i[21], \rbus_ring_i.rd_data [19]);
tran (rbus_ring_i[20], \rbus_ring_i.rd_data [18]);
tran (rbus_ring_i[19], \rbus_ring_i.rd_data [17]);
tran (rbus_ring_i[18], \rbus_ring_i.rd_data [16]);
tran (rbus_ring_i[17], \rbus_ring_i.rd_data [15]);
tran (rbus_ring_i[16], \rbus_ring_i.rd_data [14]);
tran (rbus_ring_i[15], \rbus_ring_i.rd_data [13]);
tran (rbus_ring_i[14], \rbus_ring_i.rd_data [12]);
tran (rbus_ring_i[13], \rbus_ring_i.rd_data [11]);
tran (rbus_ring_i[12], \rbus_ring_i.rd_data [10]);
tran (rbus_ring_i[11], \rbus_ring_i.rd_data [9]);
tran (rbus_ring_i[10], \rbus_ring_i.rd_data [8]);
tran (rbus_ring_i[9], \rbus_ring_i.rd_data [7]);
tran (rbus_ring_i[8], \rbus_ring_i.rd_data [6]);
tran (rbus_ring_i[7], \rbus_ring_i.rd_data [5]);
tran (rbus_ring_i[6], \rbus_ring_i.rd_data [4]);
tran (rbus_ring_i[5], \rbus_ring_i.rd_data [3]);
tran (rbus_ring_i[4], \rbus_ring_i.rd_data [2]);
tran (rbus_ring_i[3], \rbus_ring_i.rd_data [1]);
tran (rbus_ring_i[2], \rbus_ring_i.rd_data [0]);
tran (\sa_snapshot[31][63] , \sa_snapshot[31].r.part1[31] );
tran (\sa_snapshot[31][63] , \sa_snapshot[31].f.unused[13] );
tran (\sa_snapshot[31][62] , \sa_snapshot[31].r.part1[30] );
tran (\sa_snapshot[31][62] , \sa_snapshot[31].f.unused[12] );
tran (\sa_snapshot[31][61] , \sa_snapshot[31].r.part1[29] );
tran (\sa_snapshot[31][61] , \sa_snapshot[31].f.unused[11] );
tran (\sa_snapshot[31][60] , \sa_snapshot[31].r.part1[28] );
tran (\sa_snapshot[31][60] , \sa_snapshot[31].f.unused[10] );
tran (\sa_snapshot[31][59] , \sa_snapshot[31].r.part1[27] );
tran (\sa_snapshot[31][59] , \sa_snapshot[31].f.unused[9] );
tran (\sa_snapshot[31][58] , \sa_snapshot[31].r.part1[26] );
tran (\sa_snapshot[31][58] , \sa_snapshot[31].f.unused[8] );
tran (\sa_snapshot[31][57] , \sa_snapshot[31].r.part1[25] );
tran (\sa_snapshot[31][57] , \sa_snapshot[31].f.unused[7] );
tran (\sa_snapshot[31][56] , \sa_snapshot[31].r.part1[24] );
tran (\sa_snapshot[31][56] , \sa_snapshot[31].f.unused[6] );
tran (\sa_snapshot[31][55] , \sa_snapshot[31].r.part1[23] );
tran (\sa_snapshot[31][55] , \sa_snapshot[31].f.unused[5] );
tran (\sa_snapshot[31][54] , \sa_snapshot[31].r.part1[22] );
tran (\sa_snapshot[31][54] , \sa_snapshot[31].f.unused[4] );
tran (\sa_snapshot[31][53] , \sa_snapshot[31].r.part1[21] );
tran (\sa_snapshot[31][53] , \sa_snapshot[31].f.unused[3] );
tran (\sa_snapshot[31][52] , \sa_snapshot[31].r.part1[20] );
tran (\sa_snapshot[31][52] , \sa_snapshot[31].f.unused[2] );
tran (\sa_snapshot[31][51] , \sa_snapshot[31].r.part1[19] );
tran (\sa_snapshot[31][51] , \sa_snapshot[31].f.unused[1] );
tran (\sa_snapshot[31][50] , \sa_snapshot[31].r.part1[18] );
tran (\sa_snapshot[31][50] , \sa_snapshot[31].f.unused[0] );
tran (\sa_snapshot[31][49] , \sa_snapshot[31].r.part1[17] );
tran (\sa_snapshot[31][49] , \sa_snapshot[31].f.upper[17] );
tran (\sa_snapshot[31][48] , \sa_snapshot[31].r.part1[16] );
tran (\sa_snapshot[31][48] , \sa_snapshot[31].f.upper[16] );
tran (\sa_snapshot[31][47] , \sa_snapshot[31].r.part1[15] );
tran (\sa_snapshot[31][47] , \sa_snapshot[31].f.upper[15] );
tran (\sa_snapshot[31][46] , \sa_snapshot[31].r.part1[14] );
tran (\sa_snapshot[31][46] , \sa_snapshot[31].f.upper[14] );
tran (\sa_snapshot[31][45] , \sa_snapshot[31].r.part1[13] );
tran (\sa_snapshot[31][45] , \sa_snapshot[31].f.upper[13] );
tran (\sa_snapshot[31][44] , \sa_snapshot[31].r.part1[12] );
tran (\sa_snapshot[31][44] , \sa_snapshot[31].f.upper[12] );
tran (\sa_snapshot[31][43] , \sa_snapshot[31].r.part1[11] );
tran (\sa_snapshot[31][43] , \sa_snapshot[31].f.upper[11] );
tran (\sa_snapshot[31][42] , \sa_snapshot[31].r.part1[10] );
tran (\sa_snapshot[31][42] , \sa_snapshot[31].f.upper[10] );
tran (\sa_snapshot[31][41] , \sa_snapshot[31].r.part1[9] );
tran (\sa_snapshot[31][41] , \sa_snapshot[31].f.upper[9] );
tran (\sa_snapshot[31][40] , \sa_snapshot[31].r.part1[8] );
tran (\sa_snapshot[31][40] , \sa_snapshot[31].f.upper[8] );
tran (\sa_snapshot[31][39] , \sa_snapshot[31].r.part1[7] );
tran (\sa_snapshot[31][39] , \sa_snapshot[31].f.upper[7] );
tran (\sa_snapshot[31][38] , \sa_snapshot[31].r.part1[6] );
tran (\sa_snapshot[31][38] , \sa_snapshot[31].f.upper[6] );
tran (\sa_snapshot[31][37] , \sa_snapshot[31].r.part1[5] );
tran (\sa_snapshot[31][37] , \sa_snapshot[31].f.upper[5] );
tran (\sa_snapshot[31][36] , \sa_snapshot[31].r.part1[4] );
tran (\sa_snapshot[31][36] , \sa_snapshot[31].f.upper[4] );
tran (\sa_snapshot[31][35] , \sa_snapshot[31].r.part1[3] );
tran (\sa_snapshot[31][35] , \sa_snapshot[31].f.upper[3] );
tran (\sa_snapshot[31][34] , \sa_snapshot[31].r.part1[2] );
tran (\sa_snapshot[31][34] , \sa_snapshot[31].f.upper[2] );
tran (\sa_snapshot[31][33] , \sa_snapshot[31].r.part1[1] );
tran (\sa_snapshot[31][33] , \sa_snapshot[31].f.upper[1] );
tran (\sa_snapshot[31][32] , \sa_snapshot[31].r.part1[0] );
tran (\sa_snapshot[31][32] , \sa_snapshot[31].f.upper[0] );
tran (\sa_snapshot[31][31] , \sa_snapshot[31].r.part0[31] );
tran (\sa_snapshot[31][31] , \sa_snapshot[31].f.lower[31] );
tran (\sa_snapshot[31][30] , \sa_snapshot[31].r.part0[30] );
tran (\sa_snapshot[31][30] , \sa_snapshot[31].f.lower[30] );
tran (\sa_snapshot[31][29] , \sa_snapshot[31].r.part0[29] );
tran (\sa_snapshot[31][29] , \sa_snapshot[31].f.lower[29] );
tran (\sa_snapshot[31][28] , \sa_snapshot[31].r.part0[28] );
tran (\sa_snapshot[31][28] , \sa_snapshot[31].f.lower[28] );
tran (\sa_snapshot[31][27] , \sa_snapshot[31].r.part0[27] );
tran (\sa_snapshot[31][27] , \sa_snapshot[31].f.lower[27] );
tran (\sa_snapshot[31][26] , \sa_snapshot[31].r.part0[26] );
tran (\sa_snapshot[31][26] , \sa_snapshot[31].f.lower[26] );
tran (\sa_snapshot[31][25] , \sa_snapshot[31].r.part0[25] );
tran (\sa_snapshot[31][25] , \sa_snapshot[31].f.lower[25] );
tran (\sa_snapshot[31][24] , \sa_snapshot[31].r.part0[24] );
tran (\sa_snapshot[31][24] , \sa_snapshot[31].f.lower[24] );
tran (\sa_snapshot[31][23] , \sa_snapshot[31].r.part0[23] );
tran (\sa_snapshot[31][23] , \sa_snapshot[31].f.lower[23] );
tran (\sa_snapshot[31][22] , \sa_snapshot[31].r.part0[22] );
tran (\sa_snapshot[31][22] , \sa_snapshot[31].f.lower[22] );
tran (\sa_snapshot[31][21] , \sa_snapshot[31].r.part0[21] );
tran (\sa_snapshot[31][21] , \sa_snapshot[31].f.lower[21] );
tran (\sa_snapshot[31][20] , \sa_snapshot[31].r.part0[20] );
tran (\sa_snapshot[31][20] , \sa_snapshot[31].f.lower[20] );
tran (\sa_snapshot[31][19] , \sa_snapshot[31].r.part0[19] );
tran (\sa_snapshot[31][19] , \sa_snapshot[31].f.lower[19] );
tran (\sa_snapshot[31][18] , \sa_snapshot[31].r.part0[18] );
tran (\sa_snapshot[31][18] , \sa_snapshot[31].f.lower[18] );
tran (\sa_snapshot[31][17] , \sa_snapshot[31].r.part0[17] );
tran (\sa_snapshot[31][17] , \sa_snapshot[31].f.lower[17] );
tran (\sa_snapshot[31][16] , \sa_snapshot[31].r.part0[16] );
tran (\sa_snapshot[31][16] , \sa_snapshot[31].f.lower[16] );
tran (\sa_snapshot[31][15] , \sa_snapshot[31].r.part0[15] );
tran (\sa_snapshot[31][15] , \sa_snapshot[31].f.lower[15] );
tran (\sa_snapshot[31][14] , \sa_snapshot[31].r.part0[14] );
tran (\sa_snapshot[31][14] , \sa_snapshot[31].f.lower[14] );
tran (\sa_snapshot[31][13] , \sa_snapshot[31].r.part0[13] );
tran (\sa_snapshot[31][13] , \sa_snapshot[31].f.lower[13] );
tran (\sa_snapshot[31][12] , \sa_snapshot[31].r.part0[12] );
tran (\sa_snapshot[31][12] , \sa_snapshot[31].f.lower[12] );
tran (\sa_snapshot[31][11] , \sa_snapshot[31].r.part0[11] );
tran (\sa_snapshot[31][11] , \sa_snapshot[31].f.lower[11] );
tran (\sa_snapshot[31][10] , \sa_snapshot[31].r.part0[10] );
tran (\sa_snapshot[31][10] , \sa_snapshot[31].f.lower[10] );
tran (\sa_snapshot[31][9] , \sa_snapshot[31].r.part0[9] );
tran (\sa_snapshot[31][9] , \sa_snapshot[31].f.lower[9] );
tran (\sa_snapshot[31][8] , \sa_snapshot[31].r.part0[8] );
tran (\sa_snapshot[31][8] , \sa_snapshot[31].f.lower[8] );
tran (\sa_snapshot[31][7] , \sa_snapshot[31].r.part0[7] );
tran (\sa_snapshot[31][7] , \sa_snapshot[31].f.lower[7] );
tran (\sa_snapshot[31][6] , \sa_snapshot[31].r.part0[6] );
tran (\sa_snapshot[31][6] , \sa_snapshot[31].f.lower[6] );
tran (\sa_snapshot[31][5] , \sa_snapshot[31].r.part0[5] );
tran (\sa_snapshot[31][5] , \sa_snapshot[31].f.lower[5] );
tran (\sa_snapshot[31][4] , \sa_snapshot[31].r.part0[4] );
tran (\sa_snapshot[31][4] , \sa_snapshot[31].f.lower[4] );
tran (\sa_snapshot[31][3] , \sa_snapshot[31].r.part0[3] );
tran (\sa_snapshot[31][3] , \sa_snapshot[31].f.lower[3] );
tran (\sa_snapshot[31][2] , \sa_snapshot[31].r.part0[2] );
tran (\sa_snapshot[31][2] , \sa_snapshot[31].f.lower[2] );
tran (\sa_snapshot[31][1] , \sa_snapshot[31].r.part0[1] );
tran (\sa_snapshot[31][1] , \sa_snapshot[31].f.lower[1] );
tran (\sa_snapshot[31][0] , \sa_snapshot[31].r.part0[0] );
tran (\sa_snapshot[31][0] , \sa_snapshot[31].f.lower[0] );
tran (\sa_snapshot[30][63] , \sa_snapshot[30].r.part1[31] );
tran (\sa_snapshot[30][63] , \sa_snapshot[30].f.unused[13] );
tran (\sa_snapshot[30][62] , \sa_snapshot[30].r.part1[30] );
tran (\sa_snapshot[30][62] , \sa_snapshot[30].f.unused[12] );
tran (\sa_snapshot[30][61] , \sa_snapshot[30].r.part1[29] );
tran (\sa_snapshot[30][61] , \sa_snapshot[30].f.unused[11] );
tran (\sa_snapshot[30][60] , \sa_snapshot[30].r.part1[28] );
tran (\sa_snapshot[30][60] , \sa_snapshot[30].f.unused[10] );
tran (\sa_snapshot[30][59] , \sa_snapshot[30].r.part1[27] );
tran (\sa_snapshot[30][59] , \sa_snapshot[30].f.unused[9] );
tran (\sa_snapshot[30][58] , \sa_snapshot[30].r.part1[26] );
tran (\sa_snapshot[30][58] , \sa_snapshot[30].f.unused[8] );
tran (\sa_snapshot[30][57] , \sa_snapshot[30].r.part1[25] );
tran (\sa_snapshot[30][57] , \sa_snapshot[30].f.unused[7] );
tran (\sa_snapshot[30][56] , \sa_snapshot[30].r.part1[24] );
tran (\sa_snapshot[30][56] , \sa_snapshot[30].f.unused[6] );
tran (\sa_snapshot[30][55] , \sa_snapshot[30].r.part1[23] );
tran (\sa_snapshot[30][55] , \sa_snapshot[30].f.unused[5] );
tran (\sa_snapshot[30][54] , \sa_snapshot[30].r.part1[22] );
tran (\sa_snapshot[30][54] , \sa_snapshot[30].f.unused[4] );
tran (\sa_snapshot[30][53] , \sa_snapshot[30].r.part1[21] );
tran (\sa_snapshot[30][53] , \sa_snapshot[30].f.unused[3] );
tran (\sa_snapshot[30][52] , \sa_snapshot[30].r.part1[20] );
tran (\sa_snapshot[30][52] , \sa_snapshot[30].f.unused[2] );
tran (\sa_snapshot[30][51] , \sa_snapshot[30].r.part1[19] );
tran (\sa_snapshot[30][51] , \sa_snapshot[30].f.unused[1] );
tran (\sa_snapshot[30][50] , \sa_snapshot[30].r.part1[18] );
tran (\sa_snapshot[30][50] , \sa_snapshot[30].f.unused[0] );
tran (\sa_snapshot[30][49] , \sa_snapshot[30].r.part1[17] );
tran (\sa_snapshot[30][49] , \sa_snapshot[30].f.upper[17] );
tran (\sa_snapshot[30][48] , \sa_snapshot[30].r.part1[16] );
tran (\sa_snapshot[30][48] , \sa_snapshot[30].f.upper[16] );
tran (\sa_snapshot[30][47] , \sa_snapshot[30].r.part1[15] );
tran (\sa_snapshot[30][47] , \sa_snapshot[30].f.upper[15] );
tran (\sa_snapshot[30][46] , \sa_snapshot[30].r.part1[14] );
tran (\sa_snapshot[30][46] , \sa_snapshot[30].f.upper[14] );
tran (\sa_snapshot[30][45] , \sa_snapshot[30].r.part1[13] );
tran (\sa_snapshot[30][45] , \sa_snapshot[30].f.upper[13] );
tran (\sa_snapshot[30][44] , \sa_snapshot[30].r.part1[12] );
tran (\sa_snapshot[30][44] , \sa_snapshot[30].f.upper[12] );
tran (\sa_snapshot[30][43] , \sa_snapshot[30].r.part1[11] );
tran (\sa_snapshot[30][43] , \sa_snapshot[30].f.upper[11] );
tran (\sa_snapshot[30][42] , \sa_snapshot[30].r.part1[10] );
tran (\sa_snapshot[30][42] , \sa_snapshot[30].f.upper[10] );
tran (\sa_snapshot[30][41] , \sa_snapshot[30].r.part1[9] );
tran (\sa_snapshot[30][41] , \sa_snapshot[30].f.upper[9] );
tran (\sa_snapshot[30][40] , \sa_snapshot[30].r.part1[8] );
tran (\sa_snapshot[30][40] , \sa_snapshot[30].f.upper[8] );
tran (\sa_snapshot[30][39] , \sa_snapshot[30].r.part1[7] );
tran (\sa_snapshot[30][39] , \sa_snapshot[30].f.upper[7] );
tran (\sa_snapshot[30][38] , \sa_snapshot[30].r.part1[6] );
tran (\sa_snapshot[30][38] , \sa_snapshot[30].f.upper[6] );
tran (\sa_snapshot[30][37] , \sa_snapshot[30].r.part1[5] );
tran (\sa_snapshot[30][37] , \sa_snapshot[30].f.upper[5] );
tran (\sa_snapshot[30][36] , \sa_snapshot[30].r.part1[4] );
tran (\sa_snapshot[30][36] , \sa_snapshot[30].f.upper[4] );
tran (\sa_snapshot[30][35] , \sa_snapshot[30].r.part1[3] );
tran (\sa_snapshot[30][35] , \sa_snapshot[30].f.upper[3] );
tran (\sa_snapshot[30][34] , \sa_snapshot[30].r.part1[2] );
tran (\sa_snapshot[30][34] , \sa_snapshot[30].f.upper[2] );
tran (\sa_snapshot[30][33] , \sa_snapshot[30].r.part1[1] );
tran (\sa_snapshot[30][33] , \sa_snapshot[30].f.upper[1] );
tran (\sa_snapshot[30][32] , \sa_snapshot[30].r.part1[0] );
tran (\sa_snapshot[30][32] , \sa_snapshot[30].f.upper[0] );
tran (\sa_snapshot[30][31] , \sa_snapshot[30].r.part0[31] );
tran (\sa_snapshot[30][31] , \sa_snapshot[30].f.lower[31] );
tran (\sa_snapshot[30][30] , \sa_snapshot[30].r.part0[30] );
tran (\sa_snapshot[30][30] , \sa_snapshot[30].f.lower[30] );
tran (\sa_snapshot[30][29] , \sa_snapshot[30].r.part0[29] );
tran (\sa_snapshot[30][29] , \sa_snapshot[30].f.lower[29] );
tran (\sa_snapshot[30][28] , \sa_snapshot[30].r.part0[28] );
tran (\sa_snapshot[30][28] , \sa_snapshot[30].f.lower[28] );
tran (\sa_snapshot[30][27] , \sa_snapshot[30].r.part0[27] );
tran (\sa_snapshot[30][27] , \sa_snapshot[30].f.lower[27] );
tran (\sa_snapshot[30][26] , \sa_snapshot[30].r.part0[26] );
tran (\sa_snapshot[30][26] , \sa_snapshot[30].f.lower[26] );
tran (\sa_snapshot[30][25] , \sa_snapshot[30].r.part0[25] );
tran (\sa_snapshot[30][25] , \sa_snapshot[30].f.lower[25] );
tran (\sa_snapshot[30][24] , \sa_snapshot[30].r.part0[24] );
tran (\sa_snapshot[30][24] , \sa_snapshot[30].f.lower[24] );
tran (\sa_snapshot[30][23] , \sa_snapshot[30].r.part0[23] );
tran (\sa_snapshot[30][23] , \sa_snapshot[30].f.lower[23] );
tran (\sa_snapshot[30][22] , \sa_snapshot[30].r.part0[22] );
tran (\sa_snapshot[30][22] , \sa_snapshot[30].f.lower[22] );
tran (\sa_snapshot[30][21] , \sa_snapshot[30].r.part0[21] );
tran (\sa_snapshot[30][21] , \sa_snapshot[30].f.lower[21] );
tran (\sa_snapshot[30][20] , \sa_snapshot[30].r.part0[20] );
tran (\sa_snapshot[30][20] , \sa_snapshot[30].f.lower[20] );
tran (\sa_snapshot[30][19] , \sa_snapshot[30].r.part0[19] );
tran (\sa_snapshot[30][19] , \sa_snapshot[30].f.lower[19] );
tran (\sa_snapshot[30][18] , \sa_snapshot[30].r.part0[18] );
tran (\sa_snapshot[30][18] , \sa_snapshot[30].f.lower[18] );
tran (\sa_snapshot[30][17] , \sa_snapshot[30].r.part0[17] );
tran (\sa_snapshot[30][17] , \sa_snapshot[30].f.lower[17] );
tran (\sa_snapshot[30][16] , \sa_snapshot[30].r.part0[16] );
tran (\sa_snapshot[30][16] , \sa_snapshot[30].f.lower[16] );
tran (\sa_snapshot[30][15] , \sa_snapshot[30].r.part0[15] );
tran (\sa_snapshot[30][15] , \sa_snapshot[30].f.lower[15] );
tran (\sa_snapshot[30][14] , \sa_snapshot[30].r.part0[14] );
tran (\sa_snapshot[30][14] , \sa_snapshot[30].f.lower[14] );
tran (\sa_snapshot[30][13] , \sa_snapshot[30].r.part0[13] );
tran (\sa_snapshot[30][13] , \sa_snapshot[30].f.lower[13] );
tran (\sa_snapshot[30][12] , \sa_snapshot[30].r.part0[12] );
tran (\sa_snapshot[30][12] , \sa_snapshot[30].f.lower[12] );
tran (\sa_snapshot[30][11] , \sa_snapshot[30].r.part0[11] );
tran (\sa_snapshot[30][11] , \sa_snapshot[30].f.lower[11] );
tran (\sa_snapshot[30][10] , \sa_snapshot[30].r.part0[10] );
tran (\sa_snapshot[30][10] , \sa_snapshot[30].f.lower[10] );
tran (\sa_snapshot[30][9] , \sa_snapshot[30].r.part0[9] );
tran (\sa_snapshot[30][9] , \sa_snapshot[30].f.lower[9] );
tran (\sa_snapshot[30][8] , \sa_snapshot[30].r.part0[8] );
tran (\sa_snapshot[30][8] , \sa_snapshot[30].f.lower[8] );
tran (\sa_snapshot[30][7] , \sa_snapshot[30].r.part0[7] );
tran (\sa_snapshot[30][7] , \sa_snapshot[30].f.lower[7] );
tran (\sa_snapshot[30][6] , \sa_snapshot[30].r.part0[6] );
tran (\sa_snapshot[30][6] , \sa_snapshot[30].f.lower[6] );
tran (\sa_snapshot[30][5] , \sa_snapshot[30].r.part0[5] );
tran (\sa_snapshot[30][5] , \sa_snapshot[30].f.lower[5] );
tran (\sa_snapshot[30][4] , \sa_snapshot[30].r.part0[4] );
tran (\sa_snapshot[30][4] , \sa_snapshot[30].f.lower[4] );
tran (\sa_snapshot[30][3] , \sa_snapshot[30].r.part0[3] );
tran (\sa_snapshot[30][3] , \sa_snapshot[30].f.lower[3] );
tran (\sa_snapshot[30][2] , \sa_snapshot[30].r.part0[2] );
tran (\sa_snapshot[30][2] , \sa_snapshot[30].f.lower[2] );
tran (\sa_snapshot[30][1] , \sa_snapshot[30].r.part0[1] );
tran (\sa_snapshot[30][1] , \sa_snapshot[30].f.lower[1] );
tran (\sa_snapshot[30][0] , \sa_snapshot[30].r.part0[0] );
tran (\sa_snapshot[30][0] , \sa_snapshot[30].f.lower[0] );
tran (\sa_snapshot[29][63] , \sa_snapshot[29].r.part1[31] );
tran (\sa_snapshot[29][63] , \sa_snapshot[29].f.unused[13] );
tran (\sa_snapshot[29][62] , \sa_snapshot[29].r.part1[30] );
tran (\sa_snapshot[29][62] , \sa_snapshot[29].f.unused[12] );
tran (\sa_snapshot[29][61] , \sa_snapshot[29].r.part1[29] );
tran (\sa_snapshot[29][61] , \sa_snapshot[29].f.unused[11] );
tran (\sa_snapshot[29][60] , \sa_snapshot[29].r.part1[28] );
tran (\sa_snapshot[29][60] , \sa_snapshot[29].f.unused[10] );
tran (\sa_snapshot[29][59] , \sa_snapshot[29].r.part1[27] );
tran (\sa_snapshot[29][59] , \sa_snapshot[29].f.unused[9] );
tran (\sa_snapshot[29][58] , \sa_snapshot[29].r.part1[26] );
tran (\sa_snapshot[29][58] , \sa_snapshot[29].f.unused[8] );
tran (\sa_snapshot[29][57] , \sa_snapshot[29].r.part1[25] );
tran (\sa_snapshot[29][57] , \sa_snapshot[29].f.unused[7] );
tran (\sa_snapshot[29][56] , \sa_snapshot[29].r.part1[24] );
tran (\sa_snapshot[29][56] , \sa_snapshot[29].f.unused[6] );
tran (\sa_snapshot[29][55] , \sa_snapshot[29].r.part1[23] );
tran (\sa_snapshot[29][55] , \sa_snapshot[29].f.unused[5] );
tran (\sa_snapshot[29][54] , \sa_snapshot[29].r.part1[22] );
tran (\sa_snapshot[29][54] , \sa_snapshot[29].f.unused[4] );
tran (\sa_snapshot[29][53] , \sa_snapshot[29].r.part1[21] );
tran (\sa_snapshot[29][53] , \sa_snapshot[29].f.unused[3] );
tran (\sa_snapshot[29][52] , \sa_snapshot[29].r.part1[20] );
tran (\sa_snapshot[29][52] , \sa_snapshot[29].f.unused[2] );
tran (\sa_snapshot[29][51] , \sa_snapshot[29].r.part1[19] );
tran (\sa_snapshot[29][51] , \sa_snapshot[29].f.unused[1] );
tran (\sa_snapshot[29][50] , \sa_snapshot[29].r.part1[18] );
tran (\sa_snapshot[29][50] , \sa_snapshot[29].f.unused[0] );
tran (\sa_snapshot[29][49] , \sa_snapshot[29].r.part1[17] );
tran (\sa_snapshot[29][49] , \sa_snapshot[29].f.upper[17] );
tran (\sa_snapshot[29][48] , \sa_snapshot[29].r.part1[16] );
tran (\sa_snapshot[29][48] , \sa_snapshot[29].f.upper[16] );
tran (\sa_snapshot[29][47] , \sa_snapshot[29].r.part1[15] );
tran (\sa_snapshot[29][47] , \sa_snapshot[29].f.upper[15] );
tran (\sa_snapshot[29][46] , \sa_snapshot[29].r.part1[14] );
tran (\sa_snapshot[29][46] , \sa_snapshot[29].f.upper[14] );
tran (\sa_snapshot[29][45] , \sa_snapshot[29].r.part1[13] );
tran (\sa_snapshot[29][45] , \sa_snapshot[29].f.upper[13] );
tran (\sa_snapshot[29][44] , \sa_snapshot[29].r.part1[12] );
tran (\sa_snapshot[29][44] , \sa_snapshot[29].f.upper[12] );
tran (\sa_snapshot[29][43] , \sa_snapshot[29].r.part1[11] );
tran (\sa_snapshot[29][43] , \sa_snapshot[29].f.upper[11] );
tran (\sa_snapshot[29][42] , \sa_snapshot[29].r.part1[10] );
tran (\sa_snapshot[29][42] , \sa_snapshot[29].f.upper[10] );
tran (\sa_snapshot[29][41] , \sa_snapshot[29].r.part1[9] );
tran (\sa_snapshot[29][41] , \sa_snapshot[29].f.upper[9] );
tran (\sa_snapshot[29][40] , \sa_snapshot[29].r.part1[8] );
tran (\sa_snapshot[29][40] , \sa_snapshot[29].f.upper[8] );
tran (\sa_snapshot[29][39] , \sa_snapshot[29].r.part1[7] );
tran (\sa_snapshot[29][39] , \sa_snapshot[29].f.upper[7] );
tran (\sa_snapshot[29][38] , \sa_snapshot[29].r.part1[6] );
tran (\sa_snapshot[29][38] , \sa_snapshot[29].f.upper[6] );
tran (\sa_snapshot[29][37] , \sa_snapshot[29].r.part1[5] );
tran (\sa_snapshot[29][37] , \sa_snapshot[29].f.upper[5] );
tran (\sa_snapshot[29][36] , \sa_snapshot[29].r.part1[4] );
tran (\sa_snapshot[29][36] , \sa_snapshot[29].f.upper[4] );
tran (\sa_snapshot[29][35] , \sa_snapshot[29].r.part1[3] );
tran (\sa_snapshot[29][35] , \sa_snapshot[29].f.upper[3] );
tran (\sa_snapshot[29][34] , \sa_snapshot[29].r.part1[2] );
tran (\sa_snapshot[29][34] , \sa_snapshot[29].f.upper[2] );
tran (\sa_snapshot[29][33] , \sa_snapshot[29].r.part1[1] );
tran (\sa_snapshot[29][33] , \sa_snapshot[29].f.upper[1] );
tran (\sa_snapshot[29][32] , \sa_snapshot[29].r.part1[0] );
tran (\sa_snapshot[29][32] , \sa_snapshot[29].f.upper[0] );
tran (\sa_snapshot[29][31] , \sa_snapshot[29].r.part0[31] );
tran (\sa_snapshot[29][31] , \sa_snapshot[29].f.lower[31] );
tran (\sa_snapshot[29][30] , \sa_snapshot[29].r.part0[30] );
tran (\sa_snapshot[29][30] , \sa_snapshot[29].f.lower[30] );
tran (\sa_snapshot[29][29] , \sa_snapshot[29].r.part0[29] );
tran (\sa_snapshot[29][29] , \sa_snapshot[29].f.lower[29] );
tran (\sa_snapshot[29][28] , \sa_snapshot[29].r.part0[28] );
tran (\sa_snapshot[29][28] , \sa_snapshot[29].f.lower[28] );
tran (\sa_snapshot[29][27] , \sa_snapshot[29].r.part0[27] );
tran (\sa_snapshot[29][27] , \sa_snapshot[29].f.lower[27] );
tran (\sa_snapshot[29][26] , \sa_snapshot[29].r.part0[26] );
tran (\sa_snapshot[29][26] , \sa_snapshot[29].f.lower[26] );
tran (\sa_snapshot[29][25] , \sa_snapshot[29].r.part0[25] );
tran (\sa_snapshot[29][25] , \sa_snapshot[29].f.lower[25] );
tran (\sa_snapshot[29][24] , \sa_snapshot[29].r.part0[24] );
tran (\sa_snapshot[29][24] , \sa_snapshot[29].f.lower[24] );
tran (\sa_snapshot[29][23] , \sa_snapshot[29].r.part0[23] );
tran (\sa_snapshot[29][23] , \sa_snapshot[29].f.lower[23] );
tran (\sa_snapshot[29][22] , \sa_snapshot[29].r.part0[22] );
tran (\sa_snapshot[29][22] , \sa_snapshot[29].f.lower[22] );
tran (\sa_snapshot[29][21] , \sa_snapshot[29].r.part0[21] );
tran (\sa_snapshot[29][21] , \sa_snapshot[29].f.lower[21] );
tran (\sa_snapshot[29][20] , \sa_snapshot[29].r.part0[20] );
tran (\sa_snapshot[29][20] , \sa_snapshot[29].f.lower[20] );
tran (\sa_snapshot[29][19] , \sa_snapshot[29].r.part0[19] );
tran (\sa_snapshot[29][19] , \sa_snapshot[29].f.lower[19] );
tran (\sa_snapshot[29][18] , \sa_snapshot[29].r.part0[18] );
tran (\sa_snapshot[29][18] , \sa_snapshot[29].f.lower[18] );
tran (\sa_snapshot[29][17] , \sa_snapshot[29].r.part0[17] );
tran (\sa_snapshot[29][17] , \sa_snapshot[29].f.lower[17] );
tran (\sa_snapshot[29][16] , \sa_snapshot[29].r.part0[16] );
tran (\sa_snapshot[29][16] , \sa_snapshot[29].f.lower[16] );
tran (\sa_snapshot[29][15] , \sa_snapshot[29].r.part0[15] );
tran (\sa_snapshot[29][15] , \sa_snapshot[29].f.lower[15] );
tran (\sa_snapshot[29][14] , \sa_snapshot[29].r.part0[14] );
tran (\sa_snapshot[29][14] , \sa_snapshot[29].f.lower[14] );
tran (\sa_snapshot[29][13] , \sa_snapshot[29].r.part0[13] );
tran (\sa_snapshot[29][13] , \sa_snapshot[29].f.lower[13] );
tran (\sa_snapshot[29][12] , \sa_snapshot[29].r.part0[12] );
tran (\sa_snapshot[29][12] , \sa_snapshot[29].f.lower[12] );
tran (\sa_snapshot[29][11] , \sa_snapshot[29].r.part0[11] );
tran (\sa_snapshot[29][11] , \sa_snapshot[29].f.lower[11] );
tran (\sa_snapshot[29][10] , \sa_snapshot[29].r.part0[10] );
tran (\sa_snapshot[29][10] , \sa_snapshot[29].f.lower[10] );
tran (\sa_snapshot[29][9] , \sa_snapshot[29].r.part0[9] );
tran (\sa_snapshot[29][9] , \sa_snapshot[29].f.lower[9] );
tran (\sa_snapshot[29][8] , \sa_snapshot[29].r.part0[8] );
tran (\sa_snapshot[29][8] , \sa_snapshot[29].f.lower[8] );
tran (\sa_snapshot[29][7] , \sa_snapshot[29].r.part0[7] );
tran (\sa_snapshot[29][7] , \sa_snapshot[29].f.lower[7] );
tran (\sa_snapshot[29][6] , \sa_snapshot[29].r.part0[6] );
tran (\sa_snapshot[29][6] , \sa_snapshot[29].f.lower[6] );
tran (\sa_snapshot[29][5] , \sa_snapshot[29].r.part0[5] );
tran (\sa_snapshot[29][5] , \sa_snapshot[29].f.lower[5] );
tran (\sa_snapshot[29][4] , \sa_snapshot[29].r.part0[4] );
tran (\sa_snapshot[29][4] , \sa_snapshot[29].f.lower[4] );
tran (\sa_snapshot[29][3] , \sa_snapshot[29].r.part0[3] );
tran (\sa_snapshot[29][3] , \sa_snapshot[29].f.lower[3] );
tran (\sa_snapshot[29][2] , \sa_snapshot[29].r.part0[2] );
tran (\sa_snapshot[29][2] , \sa_snapshot[29].f.lower[2] );
tran (\sa_snapshot[29][1] , \sa_snapshot[29].r.part0[1] );
tran (\sa_snapshot[29][1] , \sa_snapshot[29].f.lower[1] );
tran (\sa_snapshot[29][0] , \sa_snapshot[29].r.part0[0] );
tran (\sa_snapshot[29][0] , \sa_snapshot[29].f.lower[0] );
tran (\sa_snapshot[28][63] , \sa_snapshot[28].r.part1[31] );
tran (\sa_snapshot[28][63] , \sa_snapshot[28].f.unused[13] );
tran (\sa_snapshot[28][62] , \sa_snapshot[28].r.part1[30] );
tran (\sa_snapshot[28][62] , \sa_snapshot[28].f.unused[12] );
tran (\sa_snapshot[28][61] , \sa_snapshot[28].r.part1[29] );
tran (\sa_snapshot[28][61] , \sa_snapshot[28].f.unused[11] );
tran (\sa_snapshot[28][60] , \sa_snapshot[28].r.part1[28] );
tran (\sa_snapshot[28][60] , \sa_snapshot[28].f.unused[10] );
tran (\sa_snapshot[28][59] , \sa_snapshot[28].r.part1[27] );
tran (\sa_snapshot[28][59] , \sa_snapshot[28].f.unused[9] );
tran (\sa_snapshot[28][58] , \sa_snapshot[28].r.part1[26] );
tran (\sa_snapshot[28][58] , \sa_snapshot[28].f.unused[8] );
tran (\sa_snapshot[28][57] , \sa_snapshot[28].r.part1[25] );
tran (\sa_snapshot[28][57] , \sa_snapshot[28].f.unused[7] );
tran (\sa_snapshot[28][56] , \sa_snapshot[28].r.part1[24] );
tran (\sa_snapshot[28][56] , \sa_snapshot[28].f.unused[6] );
tran (\sa_snapshot[28][55] , \sa_snapshot[28].r.part1[23] );
tran (\sa_snapshot[28][55] , \sa_snapshot[28].f.unused[5] );
tran (\sa_snapshot[28][54] , \sa_snapshot[28].r.part1[22] );
tran (\sa_snapshot[28][54] , \sa_snapshot[28].f.unused[4] );
tran (\sa_snapshot[28][53] , \sa_snapshot[28].r.part1[21] );
tran (\sa_snapshot[28][53] , \sa_snapshot[28].f.unused[3] );
tran (\sa_snapshot[28][52] , \sa_snapshot[28].r.part1[20] );
tran (\sa_snapshot[28][52] , \sa_snapshot[28].f.unused[2] );
tran (\sa_snapshot[28][51] , \sa_snapshot[28].r.part1[19] );
tran (\sa_snapshot[28][51] , \sa_snapshot[28].f.unused[1] );
tran (\sa_snapshot[28][50] , \sa_snapshot[28].r.part1[18] );
tran (\sa_snapshot[28][50] , \sa_snapshot[28].f.unused[0] );
tran (\sa_snapshot[28][49] , \sa_snapshot[28].r.part1[17] );
tran (\sa_snapshot[28][49] , \sa_snapshot[28].f.upper[17] );
tran (\sa_snapshot[28][48] , \sa_snapshot[28].r.part1[16] );
tran (\sa_snapshot[28][48] , \sa_snapshot[28].f.upper[16] );
tran (\sa_snapshot[28][47] , \sa_snapshot[28].r.part1[15] );
tran (\sa_snapshot[28][47] , \sa_snapshot[28].f.upper[15] );
tran (\sa_snapshot[28][46] , \sa_snapshot[28].r.part1[14] );
tran (\sa_snapshot[28][46] , \sa_snapshot[28].f.upper[14] );
tran (\sa_snapshot[28][45] , \sa_snapshot[28].r.part1[13] );
tran (\sa_snapshot[28][45] , \sa_snapshot[28].f.upper[13] );
tran (\sa_snapshot[28][44] , \sa_snapshot[28].r.part1[12] );
tran (\sa_snapshot[28][44] , \sa_snapshot[28].f.upper[12] );
tran (\sa_snapshot[28][43] , \sa_snapshot[28].r.part1[11] );
tran (\sa_snapshot[28][43] , \sa_snapshot[28].f.upper[11] );
tran (\sa_snapshot[28][42] , \sa_snapshot[28].r.part1[10] );
tran (\sa_snapshot[28][42] , \sa_snapshot[28].f.upper[10] );
tran (\sa_snapshot[28][41] , \sa_snapshot[28].r.part1[9] );
tran (\sa_snapshot[28][41] , \sa_snapshot[28].f.upper[9] );
tran (\sa_snapshot[28][40] , \sa_snapshot[28].r.part1[8] );
tran (\sa_snapshot[28][40] , \sa_snapshot[28].f.upper[8] );
tran (\sa_snapshot[28][39] , \sa_snapshot[28].r.part1[7] );
tran (\sa_snapshot[28][39] , \sa_snapshot[28].f.upper[7] );
tran (\sa_snapshot[28][38] , \sa_snapshot[28].r.part1[6] );
tran (\sa_snapshot[28][38] , \sa_snapshot[28].f.upper[6] );
tran (\sa_snapshot[28][37] , \sa_snapshot[28].r.part1[5] );
tran (\sa_snapshot[28][37] , \sa_snapshot[28].f.upper[5] );
tran (\sa_snapshot[28][36] , \sa_snapshot[28].r.part1[4] );
tran (\sa_snapshot[28][36] , \sa_snapshot[28].f.upper[4] );
tran (\sa_snapshot[28][35] , \sa_snapshot[28].r.part1[3] );
tran (\sa_snapshot[28][35] , \sa_snapshot[28].f.upper[3] );
tran (\sa_snapshot[28][34] , \sa_snapshot[28].r.part1[2] );
tran (\sa_snapshot[28][34] , \sa_snapshot[28].f.upper[2] );
tran (\sa_snapshot[28][33] , \sa_snapshot[28].r.part1[1] );
tran (\sa_snapshot[28][33] , \sa_snapshot[28].f.upper[1] );
tran (\sa_snapshot[28][32] , \sa_snapshot[28].r.part1[0] );
tran (\sa_snapshot[28][32] , \sa_snapshot[28].f.upper[0] );
tran (\sa_snapshot[28][31] , \sa_snapshot[28].r.part0[31] );
tran (\sa_snapshot[28][31] , \sa_snapshot[28].f.lower[31] );
tran (\sa_snapshot[28][30] , \sa_snapshot[28].r.part0[30] );
tran (\sa_snapshot[28][30] , \sa_snapshot[28].f.lower[30] );
tran (\sa_snapshot[28][29] , \sa_snapshot[28].r.part0[29] );
tran (\sa_snapshot[28][29] , \sa_snapshot[28].f.lower[29] );
tran (\sa_snapshot[28][28] , \sa_snapshot[28].r.part0[28] );
tran (\sa_snapshot[28][28] , \sa_snapshot[28].f.lower[28] );
tran (\sa_snapshot[28][27] , \sa_snapshot[28].r.part0[27] );
tran (\sa_snapshot[28][27] , \sa_snapshot[28].f.lower[27] );
tran (\sa_snapshot[28][26] , \sa_snapshot[28].r.part0[26] );
tran (\sa_snapshot[28][26] , \sa_snapshot[28].f.lower[26] );
tran (\sa_snapshot[28][25] , \sa_snapshot[28].r.part0[25] );
tran (\sa_snapshot[28][25] , \sa_snapshot[28].f.lower[25] );
tran (\sa_snapshot[28][24] , \sa_snapshot[28].r.part0[24] );
tran (\sa_snapshot[28][24] , \sa_snapshot[28].f.lower[24] );
tran (\sa_snapshot[28][23] , \sa_snapshot[28].r.part0[23] );
tran (\sa_snapshot[28][23] , \sa_snapshot[28].f.lower[23] );
tran (\sa_snapshot[28][22] , \sa_snapshot[28].r.part0[22] );
tran (\sa_snapshot[28][22] , \sa_snapshot[28].f.lower[22] );
tran (\sa_snapshot[28][21] , \sa_snapshot[28].r.part0[21] );
tran (\sa_snapshot[28][21] , \sa_snapshot[28].f.lower[21] );
tran (\sa_snapshot[28][20] , \sa_snapshot[28].r.part0[20] );
tran (\sa_snapshot[28][20] , \sa_snapshot[28].f.lower[20] );
tran (\sa_snapshot[28][19] , \sa_snapshot[28].r.part0[19] );
tran (\sa_snapshot[28][19] , \sa_snapshot[28].f.lower[19] );
tran (\sa_snapshot[28][18] , \sa_snapshot[28].r.part0[18] );
tran (\sa_snapshot[28][18] , \sa_snapshot[28].f.lower[18] );
tran (\sa_snapshot[28][17] , \sa_snapshot[28].r.part0[17] );
tran (\sa_snapshot[28][17] , \sa_snapshot[28].f.lower[17] );
tran (\sa_snapshot[28][16] , \sa_snapshot[28].r.part0[16] );
tran (\sa_snapshot[28][16] , \sa_snapshot[28].f.lower[16] );
tran (\sa_snapshot[28][15] , \sa_snapshot[28].r.part0[15] );
tran (\sa_snapshot[28][15] , \sa_snapshot[28].f.lower[15] );
tran (\sa_snapshot[28][14] , \sa_snapshot[28].r.part0[14] );
tran (\sa_snapshot[28][14] , \sa_snapshot[28].f.lower[14] );
tran (\sa_snapshot[28][13] , \sa_snapshot[28].r.part0[13] );
tran (\sa_snapshot[28][13] , \sa_snapshot[28].f.lower[13] );
tran (\sa_snapshot[28][12] , \sa_snapshot[28].r.part0[12] );
tran (\sa_snapshot[28][12] , \sa_snapshot[28].f.lower[12] );
tran (\sa_snapshot[28][11] , \sa_snapshot[28].r.part0[11] );
tran (\sa_snapshot[28][11] , \sa_snapshot[28].f.lower[11] );
tran (\sa_snapshot[28][10] , \sa_snapshot[28].r.part0[10] );
tran (\sa_snapshot[28][10] , \sa_snapshot[28].f.lower[10] );
tran (\sa_snapshot[28][9] , \sa_snapshot[28].r.part0[9] );
tran (\sa_snapshot[28][9] , \sa_snapshot[28].f.lower[9] );
tran (\sa_snapshot[28][8] , \sa_snapshot[28].r.part0[8] );
tran (\sa_snapshot[28][8] , \sa_snapshot[28].f.lower[8] );
tran (\sa_snapshot[28][7] , \sa_snapshot[28].r.part0[7] );
tran (\sa_snapshot[28][7] , \sa_snapshot[28].f.lower[7] );
tran (\sa_snapshot[28][6] , \sa_snapshot[28].r.part0[6] );
tran (\sa_snapshot[28][6] , \sa_snapshot[28].f.lower[6] );
tran (\sa_snapshot[28][5] , \sa_snapshot[28].r.part0[5] );
tran (\sa_snapshot[28][5] , \sa_snapshot[28].f.lower[5] );
tran (\sa_snapshot[28][4] , \sa_snapshot[28].r.part0[4] );
tran (\sa_snapshot[28][4] , \sa_snapshot[28].f.lower[4] );
tran (\sa_snapshot[28][3] , \sa_snapshot[28].r.part0[3] );
tran (\sa_snapshot[28][3] , \sa_snapshot[28].f.lower[3] );
tran (\sa_snapshot[28][2] , \sa_snapshot[28].r.part0[2] );
tran (\sa_snapshot[28][2] , \sa_snapshot[28].f.lower[2] );
tran (\sa_snapshot[28][1] , \sa_snapshot[28].r.part0[1] );
tran (\sa_snapshot[28][1] , \sa_snapshot[28].f.lower[1] );
tran (\sa_snapshot[28][0] , \sa_snapshot[28].r.part0[0] );
tran (\sa_snapshot[28][0] , \sa_snapshot[28].f.lower[0] );
tran (\sa_snapshot[27][63] , \sa_snapshot[27].r.part1[31] );
tran (\sa_snapshot[27][63] , \sa_snapshot[27].f.unused[13] );
tran (\sa_snapshot[27][62] , \sa_snapshot[27].r.part1[30] );
tran (\sa_snapshot[27][62] , \sa_snapshot[27].f.unused[12] );
tran (\sa_snapshot[27][61] , \sa_snapshot[27].r.part1[29] );
tran (\sa_snapshot[27][61] , \sa_snapshot[27].f.unused[11] );
tran (\sa_snapshot[27][60] , \sa_snapshot[27].r.part1[28] );
tran (\sa_snapshot[27][60] , \sa_snapshot[27].f.unused[10] );
tran (\sa_snapshot[27][59] , \sa_snapshot[27].r.part1[27] );
tran (\sa_snapshot[27][59] , \sa_snapshot[27].f.unused[9] );
tran (\sa_snapshot[27][58] , \sa_snapshot[27].r.part1[26] );
tran (\sa_snapshot[27][58] , \sa_snapshot[27].f.unused[8] );
tran (\sa_snapshot[27][57] , \sa_snapshot[27].r.part1[25] );
tran (\sa_snapshot[27][57] , \sa_snapshot[27].f.unused[7] );
tran (\sa_snapshot[27][56] , \sa_snapshot[27].r.part1[24] );
tran (\sa_snapshot[27][56] , \sa_snapshot[27].f.unused[6] );
tran (\sa_snapshot[27][55] , \sa_snapshot[27].r.part1[23] );
tran (\sa_snapshot[27][55] , \sa_snapshot[27].f.unused[5] );
tran (\sa_snapshot[27][54] , \sa_snapshot[27].r.part1[22] );
tran (\sa_snapshot[27][54] , \sa_snapshot[27].f.unused[4] );
tran (\sa_snapshot[27][53] , \sa_snapshot[27].r.part1[21] );
tran (\sa_snapshot[27][53] , \sa_snapshot[27].f.unused[3] );
tran (\sa_snapshot[27][52] , \sa_snapshot[27].r.part1[20] );
tran (\sa_snapshot[27][52] , \sa_snapshot[27].f.unused[2] );
tran (\sa_snapshot[27][51] , \sa_snapshot[27].r.part1[19] );
tran (\sa_snapshot[27][51] , \sa_snapshot[27].f.unused[1] );
tran (\sa_snapshot[27][50] , \sa_snapshot[27].r.part1[18] );
tran (\sa_snapshot[27][50] , \sa_snapshot[27].f.unused[0] );
tran (\sa_snapshot[27][49] , \sa_snapshot[27].r.part1[17] );
tran (\sa_snapshot[27][49] , \sa_snapshot[27].f.upper[17] );
tran (\sa_snapshot[27][48] , \sa_snapshot[27].r.part1[16] );
tran (\sa_snapshot[27][48] , \sa_snapshot[27].f.upper[16] );
tran (\sa_snapshot[27][47] , \sa_snapshot[27].r.part1[15] );
tran (\sa_snapshot[27][47] , \sa_snapshot[27].f.upper[15] );
tran (\sa_snapshot[27][46] , \sa_snapshot[27].r.part1[14] );
tran (\sa_snapshot[27][46] , \sa_snapshot[27].f.upper[14] );
tran (\sa_snapshot[27][45] , \sa_snapshot[27].r.part1[13] );
tran (\sa_snapshot[27][45] , \sa_snapshot[27].f.upper[13] );
tran (\sa_snapshot[27][44] , \sa_snapshot[27].r.part1[12] );
tran (\sa_snapshot[27][44] , \sa_snapshot[27].f.upper[12] );
tran (\sa_snapshot[27][43] , \sa_snapshot[27].r.part1[11] );
tran (\sa_snapshot[27][43] , \sa_snapshot[27].f.upper[11] );
tran (\sa_snapshot[27][42] , \sa_snapshot[27].r.part1[10] );
tran (\sa_snapshot[27][42] , \sa_snapshot[27].f.upper[10] );
tran (\sa_snapshot[27][41] , \sa_snapshot[27].r.part1[9] );
tran (\sa_snapshot[27][41] , \sa_snapshot[27].f.upper[9] );
tran (\sa_snapshot[27][40] , \sa_snapshot[27].r.part1[8] );
tran (\sa_snapshot[27][40] , \sa_snapshot[27].f.upper[8] );
tran (\sa_snapshot[27][39] , \sa_snapshot[27].r.part1[7] );
tran (\sa_snapshot[27][39] , \sa_snapshot[27].f.upper[7] );
tran (\sa_snapshot[27][38] , \sa_snapshot[27].r.part1[6] );
tran (\sa_snapshot[27][38] , \sa_snapshot[27].f.upper[6] );
tran (\sa_snapshot[27][37] , \sa_snapshot[27].r.part1[5] );
tran (\sa_snapshot[27][37] , \sa_snapshot[27].f.upper[5] );
tran (\sa_snapshot[27][36] , \sa_snapshot[27].r.part1[4] );
tran (\sa_snapshot[27][36] , \sa_snapshot[27].f.upper[4] );
tran (\sa_snapshot[27][35] , \sa_snapshot[27].r.part1[3] );
tran (\sa_snapshot[27][35] , \sa_snapshot[27].f.upper[3] );
tran (\sa_snapshot[27][34] , \sa_snapshot[27].r.part1[2] );
tran (\sa_snapshot[27][34] , \sa_snapshot[27].f.upper[2] );
tran (\sa_snapshot[27][33] , \sa_snapshot[27].r.part1[1] );
tran (\sa_snapshot[27][33] , \sa_snapshot[27].f.upper[1] );
tran (\sa_snapshot[27][32] , \sa_snapshot[27].r.part1[0] );
tran (\sa_snapshot[27][32] , \sa_snapshot[27].f.upper[0] );
tran (\sa_snapshot[27][31] , \sa_snapshot[27].r.part0[31] );
tran (\sa_snapshot[27][31] , \sa_snapshot[27].f.lower[31] );
tran (\sa_snapshot[27][30] , \sa_snapshot[27].r.part0[30] );
tran (\sa_snapshot[27][30] , \sa_snapshot[27].f.lower[30] );
tran (\sa_snapshot[27][29] , \sa_snapshot[27].r.part0[29] );
tran (\sa_snapshot[27][29] , \sa_snapshot[27].f.lower[29] );
tran (\sa_snapshot[27][28] , \sa_snapshot[27].r.part0[28] );
tran (\sa_snapshot[27][28] , \sa_snapshot[27].f.lower[28] );
tran (\sa_snapshot[27][27] , \sa_snapshot[27].r.part0[27] );
tran (\sa_snapshot[27][27] , \sa_snapshot[27].f.lower[27] );
tran (\sa_snapshot[27][26] , \sa_snapshot[27].r.part0[26] );
tran (\sa_snapshot[27][26] , \sa_snapshot[27].f.lower[26] );
tran (\sa_snapshot[27][25] , \sa_snapshot[27].r.part0[25] );
tran (\sa_snapshot[27][25] , \sa_snapshot[27].f.lower[25] );
tran (\sa_snapshot[27][24] , \sa_snapshot[27].r.part0[24] );
tran (\sa_snapshot[27][24] , \sa_snapshot[27].f.lower[24] );
tran (\sa_snapshot[27][23] , \sa_snapshot[27].r.part0[23] );
tran (\sa_snapshot[27][23] , \sa_snapshot[27].f.lower[23] );
tran (\sa_snapshot[27][22] , \sa_snapshot[27].r.part0[22] );
tran (\sa_snapshot[27][22] , \sa_snapshot[27].f.lower[22] );
tran (\sa_snapshot[27][21] , \sa_snapshot[27].r.part0[21] );
tran (\sa_snapshot[27][21] , \sa_snapshot[27].f.lower[21] );
tran (\sa_snapshot[27][20] , \sa_snapshot[27].r.part0[20] );
tran (\sa_snapshot[27][20] , \sa_snapshot[27].f.lower[20] );
tran (\sa_snapshot[27][19] , \sa_snapshot[27].r.part0[19] );
tran (\sa_snapshot[27][19] , \sa_snapshot[27].f.lower[19] );
tran (\sa_snapshot[27][18] , \sa_snapshot[27].r.part0[18] );
tran (\sa_snapshot[27][18] , \sa_snapshot[27].f.lower[18] );
tran (\sa_snapshot[27][17] , \sa_snapshot[27].r.part0[17] );
tran (\sa_snapshot[27][17] , \sa_snapshot[27].f.lower[17] );
tran (\sa_snapshot[27][16] , \sa_snapshot[27].r.part0[16] );
tran (\sa_snapshot[27][16] , \sa_snapshot[27].f.lower[16] );
tran (\sa_snapshot[27][15] , \sa_snapshot[27].r.part0[15] );
tran (\sa_snapshot[27][15] , \sa_snapshot[27].f.lower[15] );
tran (\sa_snapshot[27][14] , \sa_snapshot[27].r.part0[14] );
tran (\sa_snapshot[27][14] , \sa_snapshot[27].f.lower[14] );
tran (\sa_snapshot[27][13] , \sa_snapshot[27].r.part0[13] );
tran (\sa_snapshot[27][13] , \sa_snapshot[27].f.lower[13] );
tran (\sa_snapshot[27][12] , \sa_snapshot[27].r.part0[12] );
tran (\sa_snapshot[27][12] , \sa_snapshot[27].f.lower[12] );
tran (\sa_snapshot[27][11] , \sa_snapshot[27].r.part0[11] );
tran (\sa_snapshot[27][11] , \sa_snapshot[27].f.lower[11] );
tran (\sa_snapshot[27][10] , \sa_snapshot[27].r.part0[10] );
tran (\sa_snapshot[27][10] , \sa_snapshot[27].f.lower[10] );
tran (\sa_snapshot[27][9] , \sa_snapshot[27].r.part0[9] );
tran (\sa_snapshot[27][9] , \sa_snapshot[27].f.lower[9] );
tran (\sa_snapshot[27][8] , \sa_snapshot[27].r.part0[8] );
tran (\sa_snapshot[27][8] , \sa_snapshot[27].f.lower[8] );
tran (\sa_snapshot[27][7] , \sa_snapshot[27].r.part0[7] );
tran (\sa_snapshot[27][7] , \sa_snapshot[27].f.lower[7] );
tran (\sa_snapshot[27][6] , \sa_snapshot[27].r.part0[6] );
tran (\sa_snapshot[27][6] , \sa_snapshot[27].f.lower[6] );
tran (\sa_snapshot[27][5] , \sa_snapshot[27].r.part0[5] );
tran (\sa_snapshot[27][5] , \sa_snapshot[27].f.lower[5] );
tran (\sa_snapshot[27][4] , \sa_snapshot[27].r.part0[4] );
tran (\sa_snapshot[27][4] , \sa_snapshot[27].f.lower[4] );
tran (\sa_snapshot[27][3] , \sa_snapshot[27].r.part0[3] );
tran (\sa_snapshot[27][3] , \sa_snapshot[27].f.lower[3] );
tran (\sa_snapshot[27][2] , \sa_snapshot[27].r.part0[2] );
tran (\sa_snapshot[27][2] , \sa_snapshot[27].f.lower[2] );
tran (\sa_snapshot[27][1] , \sa_snapshot[27].r.part0[1] );
tran (\sa_snapshot[27][1] , \sa_snapshot[27].f.lower[1] );
tran (\sa_snapshot[27][0] , \sa_snapshot[27].r.part0[0] );
tran (\sa_snapshot[27][0] , \sa_snapshot[27].f.lower[0] );
tran (\sa_snapshot[26][63] , \sa_snapshot[26].r.part1[31] );
tran (\sa_snapshot[26][63] , \sa_snapshot[26].f.unused[13] );
tran (\sa_snapshot[26][62] , \sa_snapshot[26].r.part1[30] );
tran (\sa_snapshot[26][62] , \sa_snapshot[26].f.unused[12] );
tran (\sa_snapshot[26][61] , \sa_snapshot[26].r.part1[29] );
tran (\sa_snapshot[26][61] , \sa_snapshot[26].f.unused[11] );
tran (\sa_snapshot[26][60] , \sa_snapshot[26].r.part1[28] );
tran (\sa_snapshot[26][60] , \sa_snapshot[26].f.unused[10] );
tran (\sa_snapshot[26][59] , \sa_snapshot[26].r.part1[27] );
tran (\sa_snapshot[26][59] , \sa_snapshot[26].f.unused[9] );
tran (\sa_snapshot[26][58] , \sa_snapshot[26].r.part1[26] );
tran (\sa_snapshot[26][58] , \sa_snapshot[26].f.unused[8] );
tran (\sa_snapshot[26][57] , \sa_snapshot[26].r.part1[25] );
tran (\sa_snapshot[26][57] , \sa_snapshot[26].f.unused[7] );
tran (\sa_snapshot[26][56] , \sa_snapshot[26].r.part1[24] );
tran (\sa_snapshot[26][56] , \sa_snapshot[26].f.unused[6] );
tran (\sa_snapshot[26][55] , \sa_snapshot[26].r.part1[23] );
tran (\sa_snapshot[26][55] , \sa_snapshot[26].f.unused[5] );
tran (\sa_snapshot[26][54] , \sa_snapshot[26].r.part1[22] );
tran (\sa_snapshot[26][54] , \sa_snapshot[26].f.unused[4] );
tran (\sa_snapshot[26][53] , \sa_snapshot[26].r.part1[21] );
tran (\sa_snapshot[26][53] , \sa_snapshot[26].f.unused[3] );
tran (\sa_snapshot[26][52] , \sa_snapshot[26].r.part1[20] );
tran (\sa_snapshot[26][52] , \sa_snapshot[26].f.unused[2] );
tran (\sa_snapshot[26][51] , \sa_snapshot[26].r.part1[19] );
tran (\sa_snapshot[26][51] , \sa_snapshot[26].f.unused[1] );
tran (\sa_snapshot[26][50] , \sa_snapshot[26].r.part1[18] );
tran (\sa_snapshot[26][50] , \sa_snapshot[26].f.unused[0] );
tran (\sa_snapshot[26][49] , \sa_snapshot[26].r.part1[17] );
tran (\sa_snapshot[26][49] , \sa_snapshot[26].f.upper[17] );
tran (\sa_snapshot[26][48] , \sa_snapshot[26].r.part1[16] );
tran (\sa_snapshot[26][48] , \sa_snapshot[26].f.upper[16] );
tran (\sa_snapshot[26][47] , \sa_snapshot[26].r.part1[15] );
tran (\sa_snapshot[26][47] , \sa_snapshot[26].f.upper[15] );
tran (\sa_snapshot[26][46] , \sa_snapshot[26].r.part1[14] );
tran (\sa_snapshot[26][46] , \sa_snapshot[26].f.upper[14] );
tran (\sa_snapshot[26][45] , \sa_snapshot[26].r.part1[13] );
tran (\sa_snapshot[26][45] , \sa_snapshot[26].f.upper[13] );
tran (\sa_snapshot[26][44] , \sa_snapshot[26].r.part1[12] );
tran (\sa_snapshot[26][44] , \sa_snapshot[26].f.upper[12] );
tran (\sa_snapshot[26][43] , \sa_snapshot[26].r.part1[11] );
tran (\sa_snapshot[26][43] , \sa_snapshot[26].f.upper[11] );
tran (\sa_snapshot[26][42] , \sa_snapshot[26].r.part1[10] );
tran (\sa_snapshot[26][42] , \sa_snapshot[26].f.upper[10] );
tran (\sa_snapshot[26][41] , \sa_snapshot[26].r.part1[9] );
tran (\sa_snapshot[26][41] , \sa_snapshot[26].f.upper[9] );
tran (\sa_snapshot[26][40] , \sa_snapshot[26].r.part1[8] );
tran (\sa_snapshot[26][40] , \sa_snapshot[26].f.upper[8] );
tran (\sa_snapshot[26][39] , \sa_snapshot[26].r.part1[7] );
tran (\sa_snapshot[26][39] , \sa_snapshot[26].f.upper[7] );
tran (\sa_snapshot[26][38] , \sa_snapshot[26].r.part1[6] );
tran (\sa_snapshot[26][38] , \sa_snapshot[26].f.upper[6] );
tran (\sa_snapshot[26][37] , \sa_snapshot[26].r.part1[5] );
tran (\sa_snapshot[26][37] , \sa_snapshot[26].f.upper[5] );
tran (\sa_snapshot[26][36] , \sa_snapshot[26].r.part1[4] );
tran (\sa_snapshot[26][36] , \sa_snapshot[26].f.upper[4] );
tran (\sa_snapshot[26][35] , \sa_snapshot[26].r.part1[3] );
tran (\sa_snapshot[26][35] , \sa_snapshot[26].f.upper[3] );
tran (\sa_snapshot[26][34] , \sa_snapshot[26].r.part1[2] );
tran (\sa_snapshot[26][34] , \sa_snapshot[26].f.upper[2] );
tran (\sa_snapshot[26][33] , \sa_snapshot[26].r.part1[1] );
tran (\sa_snapshot[26][33] , \sa_snapshot[26].f.upper[1] );
tran (\sa_snapshot[26][32] , \sa_snapshot[26].r.part1[0] );
tran (\sa_snapshot[26][32] , \sa_snapshot[26].f.upper[0] );
tran (\sa_snapshot[26][31] , \sa_snapshot[26].r.part0[31] );
tran (\sa_snapshot[26][31] , \sa_snapshot[26].f.lower[31] );
tran (\sa_snapshot[26][30] , \sa_snapshot[26].r.part0[30] );
tran (\sa_snapshot[26][30] , \sa_snapshot[26].f.lower[30] );
tran (\sa_snapshot[26][29] , \sa_snapshot[26].r.part0[29] );
tran (\sa_snapshot[26][29] , \sa_snapshot[26].f.lower[29] );
tran (\sa_snapshot[26][28] , \sa_snapshot[26].r.part0[28] );
tran (\sa_snapshot[26][28] , \sa_snapshot[26].f.lower[28] );
tran (\sa_snapshot[26][27] , \sa_snapshot[26].r.part0[27] );
tran (\sa_snapshot[26][27] , \sa_snapshot[26].f.lower[27] );
tran (\sa_snapshot[26][26] , \sa_snapshot[26].r.part0[26] );
tran (\sa_snapshot[26][26] , \sa_snapshot[26].f.lower[26] );
tran (\sa_snapshot[26][25] , \sa_snapshot[26].r.part0[25] );
tran (\sa_snapshot[26][25] , \sa_snapshot[26].f.lower[25] );
tran (\sa_snapshot[26][24] , \sa_snapshot[26].r.part0[24] );
tran (\sa_snapshot[26][24] , \sa_snapshot[26].f.lower[24] );
tran (\sa_snapshot[26][23] , \sa_snapshot[26].r.part0[23] );
tran (\sa_snapshot[26][23] , \sa_snapshot[26].f.lower[23] );
tran (\sa_snapshot[26][22] , \sa_snapshot[26].r.part0[22] );
tran (\sa_snapshot[26][22] , \sa_snapshot[26].f.lower[22] );
tran (\sa_snapshot[26][21] , \sa_snapshot[26].r.part0[21] );
tran (\sa_snapshot[26][21] , \sa_snapshot[26].f.lower[21] );
tran (\sa_snapshot[26][20] , \sa_snapshot[26].r.part0[20] );
tran (\sa_snapshot[26][20] , \sa_snapshot[26].f.lower[20] );
tran (\sa_snapshot[26][19] , \sa_snapshot[26].r.part0[19] );
tran (\sa_snapshot[26][19] , \sa_snapshot[26].f.lower[19] );
tran (\sa_snapshot[26][18] , \sa_snapshot[26].r.part0[18] );
tran (\sa_snapshot[26][18] , \sa_snapshot[26].f.lower[18] );
tran (\sa_snapshot[26][17] , \sa_snapshot[26].r.part0[17] );
tran (\sa_snapshot[26][17] , \sa_snapshot[26].f.lower[17] );
tran (\sa_snapshot[26][16] , \sa_snapshot[26].r.part0[16] );
tran (\sa_snapshot[26][16] , \sa_snapshot[26].f.lower[16] );
tran (\sa_snapshot[26][15] , \sa_snapshot[26].r.part0[15] );
tran (\sa_snapshot[26][15] , \sa_snapshot[26].f.lower[15] );
tran (\sa_snapshot[26][14] , \sa_snapshot[26].r.part0[14] );
tran (\sa_snapshot[26][14] , \sa_snapshot[26].f.lower[14] );
tran (\sa_snapshot[26][13] , \sa_snapshot[26].r.part0[13] );
tran (\sa_snapshot[26][13] , \sa_snapshot[26].f.lower[13] );
tran (\sa_snapshot[26][12] , \sa_snapshot[26].r.part0[12] );
tran (\sa_snapshot[26][12] , \sa_snapshot[26].f.lower[12] );
tran (\sa_snapshot[26][11] , \sa_snapshot[26].r.part0[11] );
tran (\sa_snapshot[26][11] , \sa_snapshot[26].f.lower[11] );
tran (\sa_snapshot[26][10] , \sa_snapshot[26].r.part0[10] );
tran (\sa_snapshot[26][10] , \sa_snapshot[26].f.lower[10] );
tran (\sa_snapshot[26][9] , \sa_snapshot[26].r.part0[9] );
tran (\sa_snapshot[26][9] , \sa_snapshot[26].f.lower[9] );
tran (\sa_snapshot[26][8] , \sa_snapshot[26].r.part0[8] );
tran (\sa_snapshot[26][8] , \sa_snapshot[26].f.lower[8] );
tran (\sa_snapshot[26][7] , \sa_snapshot[26].r.part0[7] );
tran (\sa_snapshot[26][7] , \sa_snapshot[26].f.lower[7] );
tran (\sa_snapshot[26][6] , \sa_snapshot[26].r.part0[6] );
tran (\sa_snapshot[26][6] , \sa_snapshot[26].f.lower[6] );
tran (\sa_snapshot[26][5] , \sa_snapshot[26].r.part0[5] );
tran (\sa_snapshot[26][5] , \sa_snapshot[26].f.lower[5] );
tran (\sa_snapshot[26][4] , \sa_snapshot[26].r.part0[4] );
tran (\sa_snapshot[26][4] , \sa_snapshot[26].f.lower[4] );
tran (\sa_snapshot[26][3] , \sa_snapshot[26].r.part0[3] );
tran (\sa_snapshot[26][3] , \sa_snapshot[26].f.lower[3] );
tran (\sa_snapshot[26][2] , \sa_snapshot[26].r.part0[2] );
tran (\sa_snapshot[26][2] , \sa_snapshot[26].f.lower[2] );
tran (\sa_snapshot[26][1] , \sa_snapshot[26].r.part0[1] );
tran (\sa_snapshot[26][1] , \sa_snapshot[26].f.lower[1] );
tran (\sa_snapshot[26][0] , \sa_snapshot[26].r.part0[0] );
tran (\sa_snapshot[26][0] , \sa_snapshot[26].f.lower[0] );
tran (\sa_snapshot[25][63] , \sa_snapshot[25].r.part1[31] );
tran (\sa_snapshot[25][63] , \sa_snapshot[25].f.unused[13] );
tran (\sa_snapshot[25][62] , \sa_snapshot[25].r.part1[30] );
tran (\sa_snapshot[25][62] , \sa_snapshot[25].f.unused[12] );
tran (\sa_snapshot[25][61] , \sa_snapshot[25].r.part1[29] );
tran (\sa_snapshot[25][61] , \sa_snapshot[25].f.unused[11] );
tran (\sa_snapshot[25][60] , \sa_snapshot[25].r.part1[28] );
tran (\sa_snapshot[25][60] , \sa_snapshot[25].f.unused[10] );
tran (\sa_snapshot[25][59] , \sa_snapshot[25].r.part1[27] );
tran (\sa_snapshot[25][59] , \sa_snapshot[25].f.unused[9] );
tran (\sa_snapshot[25][58] , \sa_snapshot[25].r.part1[26] );
tran (\sa_snapshot[25][58] , \sa_snapshot[25].f.unused[8] );
tran (\sa_snapshot[25][57] , \sa_snapshot[25].r.part1[25] );
tran (\sa_snapshot[25][57] , \sa_snapshot[25].f.unused[7] );
tran (\sa_snapshot[25][56] , \sa_snapshot[25].r.part1[24] );
tran (\sa_snapshot[25][56] , \sa_snapshot[25].f.unused[6] );
tran (\sa_snapshot[25][55] , \sa_snapshot[25].r.part1[23] );
tran (\sa_snapshot[25][55] , \sa_snapshot[25].f.unused[5] );
tran (\sa_snapshot[25][54] , \sa_snapshot[25].r.part1[22] );
tran (\sa_snapshot[25][54] , \sa_snapshot[25].f.unused[4] );
tran (\sa_snapshot[25][53] , \sa_snapshot[25].r.part1[21] );
tran (\sa_snapshot[25][53] , \sa_snapshot[25].f.unused[3] );
tran (\sa_snapshot[25][52] , \sa_snapshot[25].r.part1[20] );
tran (\sa_snapshot[25][52] , \sa_snapshot[25].f.unused[2] );
tran (\sa_snapshot[25][51] , \sa_snapshot[25].r.part1[19] );
tran (\sa_snapshot[25][51] , \sa_snapshot[25].f.unused[1] );
tran (\sa_snapshot[25][50] , \sa_snapshot[25].r.part1[18] );
tran (\sa_snapshot[25][50] , \sa_snapshot[25].f.unused[0] );
tran (\sa_snapshot[25][49] , \sa_snapshot[25].r.part1[17] );
tran (\sa_snapshot[25][49] , \sa_snapshot[25].f.upper[17] );
tran (\sa_snapshot[25][48] , \sa_snapshot[25].r.part1[16] );
tran (\sa_snapshot[25][48] , \sa_snapshot[25].f.upper[16] );
tran (\sa_snapshot[25][47] , \sa_snapshot[25].r.part1[15] );
tran (\sa_snapshot[25][47] , \sa_snapshot[25].f.upper[15] );
tran (\sa_snapshot[25][46] , \sa_snapshot[25].r.part1[14] );
tran (\sa_snapshot[25][46] , \sa_snapshot[25].f.upper[14] );
tran (\sa_snapshot[25][45] , \sa_snapshot[25].r.part1[13] );
tran (\sa_snapshot[25][45] , \sa_snapshot[25].f.upper[13] );
tran (\sa_snapshot[25][44] , \sa_snapshot[25].r.part1[12] );
tran (\sa_snapshot[25][44] , \sa_snapshot[25].f.upper[12] );
tran (\sa_snapshot[25][43] , \sa_snapshot[25].r.part1[11] );
tran (\sa_snapshot[25][43] , \sa_snapshot[25].f.upper[11] );
tran (\sa_snapshot[25][42] , \sa_snapshot[25].r.part1[10] );
tran (\sa_snapshot[25][42] , \sa_snapshot[25].f.upper[10] );
tran (\sa_snapshot[25][41] , \sa_snapshot[25].r.part1[9] );
tran (\sa_snapshot[25][41] , \sa_snapshot[25].f.upper[9] );
tran (\sa_snapshot[25][40] , \sa_snapshot[25].r.part1[8] );
tran (\sa_snapshot[25][40] , \sa_snapshot[25].f.upper[8] );
tran (\sa_snapshot[25][39] , \sa_snapshot[25].r.part1[7] );
tran (\sa_snapshot[25][39] , \sa_snapshot[25].f.upper[7] );
tran (\sa_snapshot[25][38] , \sa_snapshot[25].r.part1[6] );
tran (\sa_snapshot[25][38] , \sa_snapshot[25].f.upper[6] );
tran (\sa_snapshot[25][37] , \sa_snapshot[25].r.part1[5] );
tran (\sa_snapshot[25][37] , \sa_snapshot[25].f.upper[5] );
tran (\sa_snapshot[25][36] , \sa_snapshot[25].r.part1[4] );
tran (\sa_snapshot[25][36] , \sa_snapshot[25].f.upper[4] );
tran (\sa_snapshot[25][35] , \sa_snapshot[25].r.part1[3] );
tran (\sa_snapshot[25][35] , \sa_snapshot[25].f.upper[3] );
tran (\sa_snapshot[25][34] , \sa_snapshot[25].r.part1[2] );
tran (\sa_snapshot[25][34] , \sa_snapshot[25].f.upper[2] );
tran (\sa_snapshot[25][33] , \sa_snapshot[25].r.part1[1] );
tran (\sa_snapshot[25][33] , \sa_snapshot[25].f.upper[1] );
tran (\sa_snapshot[25][32] , \sa_snapshot[25].r.part1[0] );
tran (\sa_snapshot[25][32] , \sa_snapshot[25].f.upper[0] );
tran (\sa_snapshot[25][31] , \sa_snapshot[25].r.part0[31] );
tran (\sa_snapshot[25][31] , \sa_snapshot[25].f.lower[31] );
tran (\sa_snapshot[25][30] , \sa_snapshot[25].r.part0[30] );
tran (\sa_snapshot[25][30] , \sa_snapshot[25].f.lower[30] );
tran (\sa_snapshot[25][29] , \sa_snapshot[25].r.part0[29] );
tran (\sa_snapshot[25][29] , \sa_snapshot[25].f.lower[29] );
tran (\sa_snapshot[25][28] , \sa_snapshot[25].r.part0[28] );
tran (\sa_snapshot[25][28] , \sa_snapshot[25].f.lower[28] );
tran (\sa_snapshot[25][27] , \sa_snapshot[25].r.part0[27] );
tran (\sa_snapshot[25][27] , \sa_snapshot[25].f.lower[27] );
tran (\sa_snapshot[25][26] , \sa_snapshot[25].r.part0[26] );
tran (\sa_snapshot[25][26] , \sa_snapshot[25].f.lower[26] );
tran (\sa_snapshot[25][25] , \sa_snapshot[25].r.part0[25] );
tran (\sa_snapshot[25][25] , \sa_snapshot[25].f.lower[25] );
tran (\sa_snapshot[25][24] , \sa_snapshot[25].r.part0[24] );
tran (\sa_snapshot[25][24] , \sa_snapshot[25].f.lower[24] );
tran (\sa_snapshot[25][23] , \sa_snapshot[25].r.part0[23] );
tran (\sa_snapshot[25][23] , \sa_snapshot[25].f.lower[23] );
tran (\sa_snapshot[25][22] , \sa_snapshot[25].r.part0[22] );
tran (\sa_snapshot[25][22] , \sa_snapshot[25].f.lower[22] );
tran (\sa_snapshot[25][21] , \sa_snapshot[25].r.part0[21] );
tran (\sa_snapshot[25][21] , \sa_snapshot[25].f.lower[21] );
tran (\sa_snapshot[25][20] , \sa_snapshot[25].r.part0[20] );
tran (\sa_snapshot[25][20] , \sa_snapshot[25].f.lower[20] );
tran (\sa_snapshot[25][19] , \sa_snapshot[25].r.part0[19] );
tran (\sa_snapshot[25][19] , \sa_snapshot[25].f.lower[19] );
tran (\sa_snapshot[25][18] , \sa_snapshot[25].r.part0[18] );
tran (\sa_snapshot[25][18] , \sa_snapshot[25].f.lower[18] );
tran (\sa_snapshot[25][17] , \sa_snapshot[25].r.part0[17] );
tran (\sa_snapshot[25][17] , \sa_snapshot[25].f.lower[17] );
tran (\sa_snapshot[25][16] , \sa_snapshot[25].r.part0[16] );
tran (\sa_snapshot[25][16] , \sa_snapshot[25].f.lower[16] );
tran (\sa_snapshot[25][15] , \sa_snapshot[25].r.part0[15] );
tran (\sa_snapshot[25][15] , \sa_snapshot[25].f.lower[15] );
tran (\sa_snapshot[25][14] , \sa_snapshot[25].r.part0[14] );
tran (\sa_snapshot[25][14] , \sa_snapshot[25].f.lower[14] );
tran (\sa_snapshot[25][13] , \sa_snapshot[25].r.part0[13] );
tran (\sa_snapshot[25][13] , \sa_snapshot[25].f.lower[13] );
tran (\sa_snapshot[25][12] , \sa_snapshot[25].r.part0[12] );
tran (\sa_snapshot[25][12] , \sa_snapshot[25].f.lower[12] );
tran (\sa_snapshot[25][11] , \sa_snapshot[25].r.part0[11] );
tran (\sa_snapshot[25][11] , \sa_snapshot[25].f.lower[11] );
tran (\sa_snapshot[25][10] , \sa_snapshot[25].r.part0[10] );
tran (\sa_snapshot[25][10] , \sa_snapshot[25].f.lower[10] );
tran (\sa_snapshot[25][9] , \sa_snapshot[25].r.part0[9] );
tran (\sa_snapshot[25][9] , \sa_snapshot[25].f.lower[9] );
tran (\sa_snapshot[25][8] , \sa_snapshot[25].r.part0[8] );
tran (\sa_snapshot[25][8] , \sa_snapshot[25].f.lower[8] );
tran (\sa_snapshot[25][7] , \sa_snapshot[25].r.part0[7] );
tran (\sa_snapshot[25][7] , \sa_snapshot[25].f.lower[7] );
tran (\sa_snapshot[25][6] , \sa_snapshot[25].r.part0[6] );
tran (\sa_snapshot[25][6] , \sa_snapshot[25].f.lower[6] );
tran (\sa_snapshot[25][5] , \sa_snapshot[25].r.part0[5] );
tran (\sa_snapshot[25][5] , \sa_snapshot[25].f.lower[5] );
tran (\sa_snapshot[25][4] , \sa_snapshot[25].r.part0[4] );
tran (\sa_snapshot[25][4] , \sa_snapshot[25].f.lower[4] );
tran (\sa_snapshot[25][3] , \sa_snapshot[25].r.part0[3] );
tran (\sa_snapshot[25][3] , \sa_snapshot[25].f.lower[3] );
tran (\sa_snapshot[25][2] , \sa_snapshot[25].r.part0[2] );
tran (\sa_snapshot[25][2] , \sa_snapshot[25].f.lower[2] );
tran (\sa_snapshot[25][1] , \sa_snapshot[25].r.part0[1] );
tran (\sa_snapshot[25][1] , \sa_snapshot[25].f.lower[1] );
tran (\sa_snapshot[25][0] , \sa_snapshot[25].r.part0[0] );
tran (\sa_snapshot[25][0] , \sa_snapshot[25].f.lower[0] );
tran (\sa_snapshot[24][63] , \sa_snapshot[24].r.part1[31] );
tran (\sa_snapshot[24][63] , \sa_snapshot[24].f.unused[13] );
tran (\sa_snapshot[24][62] , \sa_snapshot[24].r.part1[30] );
tran (\sa_snapshot[24][62] , \sa_snapshot[24].f.unused[12] );
tran (\sa_snapshot[24][61] , \sa_snapshot[24].r.part1[29] );
tran (\sa_snapshot[24][61] , \sa_snapshot[24].f.unused[11] );
tran (\sa_snapshot[24][60] , \sa_snapshot[24].r.part1[28] );
tran (\sa_snapshot[24][60] , \sa_snapshot[24].f.unused[10] );
tran (\sa_snapshot[24][59] , \sa_snapshot[24].r.part1[27] );
tran (\sa_snapshot[24][59] , \sa_snapshot[24].f.unused[9] );
tran (\sa_snapshot[24][58] , \sa_snapshot[24].r.part1[26] );
tran (\sa_snapshot[24][58] , \sa_snapshot[24].f.unused[8] );
tran (\sa_snapshot[24][57] , \sa_snapshot[24].r.part1[25] );
tran (\sa_snapshot[24][57] , \sa_snapshot[24].f.unused[7] );
tran (\sa_snapshot[24][56] , \sa_snapshot[24].r.part1[24] );
tran (\sa_snapshot[24][56] , \sa_snapshot[24].f.unused[6] );
tran (\sa_snapshot[24][55] , \sa_snapshot[24].r.part1[23] );
tran (\sa_snapshot[24][55] , \sa_snapshot[24].f.unused[5] );
tran (\sa_snapshot[24][54] , \sa_snapshot[24].r.part1[22] );
tran (\sa_snapshot[24][54] , \sa_snapshot[24].f.unused[4] );
tran (\sa_snapshot[24][53] , \sa_snapshot[24].r.part1[21] );
tran (\sa_snapshot[24][53] , \sa_snapshot[24].f.unused[3] );
tran (\sa_snapshot[24][52] , \sa_snapshot[24].r.part1[20] );
tran (\sa_snapshot[24][52] , \sa_snapshot[24].f.unused[2] );
tran (\sa_snapshot[24][51] , \sa_snapshot[24].r.part1[19] );
tran (\sa_snapshot[24][51] , \sa_snapshot[24].f.unused[1] );
tran (\sa_snapshot[24][50] , \sa_snapshot[24].r.part1[18] );
tran (\sa_snapshot[24][50] , \sa_snapshot[24].f.unused[0] );
tran (\sa_snapshot[24][49] , \sa_snapshot[24].r.part1[17] );
tran (\sa_snapshot[24][49] , \sa_snapshot[24].f.upper[17] );
tran (\sa_snapshot[24][48] , \sa_snapshot[24].r.part1[16] );
tran (\sa_snapshot[24][48] , \sa_snapshot[24].f.upper[16] );
tran (\sa_snapshot[24][47] , \sa_snapshot[24].r.part1[15] );
tran (\sa_snapshot[24][47] , \sa_snapshot[24].f.upper[15] );
tran (\sa_snapshot[24][46] , \sa_snapshot[24].r.part1[14] );
tran (\sa_snapshot[24][46] , \sa_snapshot[24].f.upper[14] );
tran (\sa_snapshot[24][45] , \sa_snapshot[24].r.part1[13] );
tran (\sa_snapshot[24][45] , \sa_snapshot[24].f.upper[13] );
tran (\sa_snapshot[24][44] , \sa_snapshot[24].r.part1[12] );
tran (\sa_snapshot[24][44] , \sa_snapshot[24].f.upper[12] );
tran (\sa_snapshot[24][43] , \sa_snapshot[24].r.part1[11] );
tran (\sa_snapshot[24][43] , \sa_snapshot[24].f.upper[11] );
tran (\sa_snapshot[24][42] , \sa_snapshot[24].r.part1[10] );
tran (\sa_snapshot[24][42] , \sa_snapshot[24].f.upper[10] );
tran (\sa_snapshot[24][41] , \sa_snapshot[24].r.part1[9] );
tran (\sa_snapshot[24][41] , \sa_snapshot[24].f.upper[9] );
tran (\sa_snapshot[24][40] , \sa_snapshot[24].r.part1[8] );
tran (\sa_snapshot[24][40] , \sa_snapshot[24].f.upper[8] );
tran (\sa_snapshot[24][39] , \sa_snapshot[24].r.part1[7] );
tran (\sa_snapshot[24][39] , \sa_snapshot[24].f.upper[7] );
tran (\sa_snapshot[24][38] , \sa_snapshot[24].r.part1[6] );
tran (\sa_snapshot[24][38] , \sa_snapshot[24].f.upper[6] );
tran (\sa_snapshot[24][37] , \sa_snapshot[24].r.part1[5] );
tran (\sa_snapshot[24][37] , \sa_snapshot[24].f.upper[5] );
tran (\sa_snapshot[24][36] , \sa_snapshot[24].r.part1[4] );
tran (\sa_snapshot[24][36] , \sa_snapshot[24].f.upper[4] );
tran (\sa_snapshot[24][35] , \sa_snapshot[24].r.part1[3] );
tran (\sa_snapshot[24][35] , \sa_snapshot[24].f.upper[3] );
tran (\sa_snapshot[24][34] , \sa_snapshot[24].r.part1[2] );
tran (\sa_snapshot[24][34] , \sa_snapshot[24].f.upper[2] );
tran (\sa_snapshot[24][33] , \sa_snapshot[24].r.part1[1] );
tran (\sa_snapshot[24][33] , \sa_snapshot[24].f.upper[1] );
tran (\sa_snapshot[24][32] , \sa_snapshot[24].r.part1[0] );
tran (\sa_snapshot[24][32] , \sa_snapshot[24].f.upper[0] );
tran (\sa_snapshot[24][31] , \sa_snapshot[24].r.part0[31] );
tran (\sa_snapshot[24][31] , \sa_snapshot[24].f.lower[31] );
tran (\sa_snapshot[24][30] , \sa_snapshot[24].r.part0[30] );
tran (\sa_snapshot[24][30] , \sa_snapshot[24].f.lower[30] );
tran (\sa_snapshot[24][29] , \sa_snapshot[24].r.part0[29] );
tran (\sa_snapshot[24][29] , \sa_snapshot[24].f.lower[29] );
tran (\sa_snapshot[24][28] , \sa_snapshot[24].r.part0[28] );
tran (\sa_snapshot[24][28] , \sa_snapshot[24].f.lower[28] );
tran (\sa_snapshot[24][27] , \sa_snapshot[24].r.part0[27] );
tran (\sa_snapshot[24][27] , \sa_snapshot[24].f.lower[27] );
tran (\sa_snapshot[24][26] , \sa_snapshot[24].r.part0[26] );
tran (\sa_snapshot[24][26] , \sa_snapshot[24].f.lower[26] );
tran (\sa_snapshot[24][25] , \sa_snapshot[24].r.part0[25] );
tran (\sa_snapshot[24][25] , \sa_snapshot[24].f.lower[25] );
tran (\sa_snapshot[24][24] , \sa_snapshot[24].r.part0[24] );
tran (\sa_snapshot[24][24] , \sa_snapshot[24].f.lower[24] );
tran (\sa_snapshot[24][23] , \sa_snapshot[24].r.part0[23] );
tran (\sa_snapshot[24][23] , \sa_snapshot[24].f.lower[23] );
tran (\sa_snapshot[24][22] , \sa_snapshot[24].r.part0[22] );
tran (\sa_snapshot[24][22] , \sa_snapshot[24].f.lower[22] );
tran (\sa_snapshot[24][21] , \sa_snapshot[24].r.part0[21] );
tran (\sa_snapshot[24][21] , \sa_snapshot[24].f.lower[21] );
tran (\sa_snapshot[24][20] , \sa_snapshot[24].r.part0[20] );
tran (\sa_snapshot[24][20] , \sa_snapshot[24].f.lower[20] );
tran (\sa_snapshot[24][19] , \sa_snapshot[24].r.part0[19] );
tran (\sa_snapshot[24][19] , \sa_snapshot[24].f.lower[19] );
tran (\sa_snapshot[24][18] , \sa_snapshot[24].r.part0[18] );
tran (\sa_snapshot[24][18] , \sa_snapshot[24].f.lower[18] );
tran (\sa_snapshot[24][17] , \sa_snapshot[24].r.part0[17] );
tran (\sa_snapshot[24][17] , \sa_snapshot[24].f.lower[17] );
tran (\sa_snapshot[24][16] , \sa_snapshot[24].r.part0[16] );
tran (\sa_snapshot[24][16] , \sa_snapshot[24].f.lower[16] );
tran (\sa_snapshot[24][15] , \sa_snapshot[24].r.part0[15] );
tran (\sa_snapshot[24][15] , \sa_snapshot[24].f.lower[15] );
tran (\sa_snapshot[24][14] , \sa_snapshot[24].r.part0[14] );
tran (\sa_snapshot[24][14] , \sa_snapshot[24].f.lower[14] );
tran (\sa_snapshot[24][13] , \sa_snapshot[24].r.part0[13] );
tran (\sa_snapshot[24][13] , \sa_snapshot[24].f.lower[13] );
tran (\sa_snapshot[24][12] , \sa_snapshot[24].r.part0[12] );
tran (\sa_snapshot[24][12] , \sa_snapshot[24].f.lower[12] );
tran (\sa_snapshot[24][11] , \sa_snapshot[24].r.part0[11] );
tran (\sa_snapshot[24][11] , \sa_snapshot[24].f.lower[11] );
tran (\sa_snapshot[24][10] , \sa_snapshot[24].r.part0[10] );
tran (\sa_snapshot[24][10] , \sa_snapshot[24].f.lower[10] );
tran (\sa_snapshot[24][9] , \sa_snapshot[24].r.part0[9] );
tran (\sa_snapshot[24][9] , \sa_snapshot[24].f.lower[9] );
tran (\sa_snapshot[24][8] , \sa_snapshot[24].r.part0[8] );
tran (\sa_snapshot[24][8] , \sa_snapshot[24].f.lower[8] );
tran (\sa_snapshot[24][7] , \sa_snapshot[24].r.part0[7] );
tran (\sa_snapshot[24][7] , \sa_snapshot[24].f.lower[7] );
tran (\sa_snapshot[24][6] , \sa_snapshot[24].r.part0[6] );
tran (\sa_snapshot[24][6] , \sa_snapshot[24].f.lower[6] );
tran (\sa_snapshot[24][5] , \sa_snapshot[24].r.part0[5] );
tran (\sa_snapshot[24][5] , \sa_snapshot[24].f.lower[5] );
tran (\sa_snapshot[24][4] , \sa_snapshot[24].r.part0[4] );
tran (\sa_snapshot[24][4] , \sa_snapshot[24].f.lower[4] );
tran (\sa_snapshot[24][3] , \sa_snapshot[24].r.part0[3] );
tran (\sa_snapshot[24][3] , \sa_snapshot[24].f.lower[3] );
tran (\sa_snapshot[24][2] , \sa_snapshot[24].r.part0[2] );
tran (\sa_snapshot[24][2] , \sa_snapshot[24].f.lower[2] );
tran (\sa_snapshot[24][1] , \sa_snapshot[24].r.part0[1] );
tran (\sa_snapshot[24][1] , \sa_snapshot[24].f.lower[1] );
tran (\sa_snapshot[24][0] , \sa_snapshot[24].r.part0[0] );
tran (\sa_snapshot[24][0] , \sa_snapshot[24].f.lower[0] );
tran (\sa_snapshot[23][63] , \sa_snapshot[23].r.part1[31] );
tran (\sa_snapshot[23][63] , \sa_snapshot[23].f.unused[13] );
tran (\sa_snapshot[23][62] , \sa_snapshot[23].r.part1[30] );
tran (\sa_snapshot[23][62] , \sa_snapshot[23].f.unused[12] );
tran (\sa_snapshot[23][61] , \sa_snapshot[23].r.part1[29] );
tran (\sa_snapshot[23][61] , \sa_snapshot[23].f.unused[11] );
tran (\sa_snapshot[23][60] , \sa_snapshot[23].r.part1[28] );
tran (\sa_snapshot[23][60] , \sa_snapshot[23].f.unused[10] );
tran (\sa_snapshot[23][59] , \sa_snapshot[23].r.part1[27] );
tran (\sa_snapshot[23][59] , \sa_snapshot[23].f.unused[9] );
tran (\sa_snapshot[23][58] , \sa_snapshot[23].r.part1[26] );
tran (\sa_snapshot[23][58] , \sa_snapshot[23].f.unused[8] );
tran (\sa_snapshot[23][57] , \sa_snapshot[23].r.part1[25] );
tran (\sa_snapshot[23][57] , \sa_snapshot[23].f.unused[7] );
tran (\sa_snapshot[23][56] , \sa_snapshot[23].r.part1[24] );
tran (\sa_snapshot[23][56] , \sa_snapshot[23].f.unused[6] );
tran (\sa_snapshot[23][55] , \sa_snapshot[23].r.part1[23] );
tran (\sa_snapshot[23][55] , \sa_snapshot[23].f.unused[5] );
tran (\sa_snapshot[23][54] , \sa_snapshot[23].r.part1[22] );
tran (\sa_snapshot[23][54] , \sa_snapshot[23].f.unused[4] );
tran (\sa_snapshot[23][53] , \sa_snapshot[23].r.part1[21] );
tran (\sa_snapshot[23][53] , \sa_snapshot[23].f.unused[3] );
tran (\sa_snapshot[23][52] , \sa_snapshot[23].r.part1[20] );
tran (\sa_snapshot[23][52] , \sa_snapshot[23].f.unused[2] );
tran (\sa_snapshot[23][51] , \sa_snapshot[23].r.part1[19] );
tran (\sa_snapshot[23][51] , \sa_snapshot[23].f.unused[1] );
tran (\sa_snapshot[23][50] , \sa_snapshot[23].r.part1[18] );
tran (\sa_snapshot[23][50] , \sa_snapshot[23].f.unused[0] );
tran (\sa_snapshot[23][49] , \sa_snapshot[23].r.part1[17] );
tran (\sa_snapshot[23][49] , \sa_snapshot[23].f.upper[17] );
tran (\sa_snapshot[23][48] , \sa_snapshot[23].r.part1[16] );
tran (\sa_snapshot[23][48] , \sa_snapshot[23].f.upper[16] );
tran (\sa_snapshot[23][47] , \sa_snapshot[23].r.part1[15] );
tran (\sa_snapshot[23][47] , \sa_snapshot[23].f.upper[15] );
tran (\sa_snapshot[23][46] , \sa_snapshot[23].r.part1[14] );
tran (\sa_snapshot[23][46] , \sa_snapshot[23].f.upper[14] );
tran (\sa_snapshot[23][45] , \sa_snapshot[23].r.part1[13] );
tran (\sa_snapshot[23][45] , \sa_snapshot[23].f.upper[13] );
tran (\sa_snapshot[23][44] , \sa_snapshot[23].r.part1[12] );
tran (\sa_snapshot[23][44] , \sa_snapshot[23].f.upper[12] );
tran (\sa_snapshot[23][43] , \sa_snapshot[23].r.part1[11] );
tran (\sa_snapshot[23][43] , \sa_snapshot[23].f.upper[11] );
tran (\sa_snapshot[23][42] , \sa_snapshot[23].r.part1[10] );
tran (\sa_snapshot[23][42] , \sa_snapshot[23].f.upper[10] );
tran (\sa_snapshot[23][41] , \sa_snapshot[23].r.part1[9] );
tran (\sa_snapshot[23][41] , \sa_snapshot[23].f.upper[9] );
tran (\sa_snapshot[23][40] , \sa_snapshot[23].r.part1[8] );
tran (\sa_snapshot[23][40] , \sa_snapshot[23].f.upper[8] );
tran (\sa_snapshot[23][39] , \sa_snapshot[23].r.part1[7] );
tran (\sa_snapshot[23][39] , \sa_snapshot[23].f.upper[7] );
tran (\sa_snapshot[23][38] , \sa_snapshot[23].r.part1[6] );
tran (\sa_snapshot[23][38] , \sa_snapshot[23].f.upper[6] );
tran (\sa_snapshot[23][37] , \sa_snapshot[23].r.part1[5] );
tran (\sa_snapshot[23][37] , \sa_snapshot[23].f.upper[5] );
tran (\sa_snapshot[23][36] , \sa_snapshot[23].r.part1[4] );
tran (\sa_snapshot[23][36] , \sa_snapshot[23].f.upper[4] );
tran (\sa_snapshot[23][35] , \sa_snapshot[23].r.part1[3] );
tran (\sa_snapshot[23][35] , \sa_snapshot[23].f.upper[3] );
tran (\sa_snapshot[23][34] , \sa_snapshot[23].r.part1[2] );
tran (\sa_snapshot[23][34] , \sa_snapshot[23].f.upper[2] );
tran (\sa_snapshot[23][33] , \sa_snapshot[23].r.part1[1] );
tran (\sa_snapshot[23][33] , \sa_snapshot[23].f.upper[1] );
tran (\sa_snapshot[23][32] , \sa_snapshot[23].r.part1[0] );
tran (\sa_snapshot[23][32] , \sa_snapshot[23].f.upper[0] );
tran (\sa_snapshot[23][31] , \sa_snapshot[23].r.part0[31] );
tran (\sa_snapshot[23][31] , \sa_snapshot[23].f.lower[31] );
tran (\sa_snapshot[23][30] , \sa_snapshot[23].r.part0[30] );
tran (\sa_snapshot[23][30] , \sa_snapshot[23].f.lower[30] );
tran (\sa_snapshot[23][29] , \sa_snapshot[23].r.part0[29] );
tran (\sa_snapshot[23][29] , \sa_snapshot[23].f.lower[29] );
tran (\sa_snapshot[23][28] , \sa_snapshot[23].r.part0[28] );
tran (\sa_snapshot[23][28] , \sa_snapshot[23].f.lower[28] );
tran (\sa_snapshot[23][27] , \sa_snapshot[23].r.part0[27] );
tran (\sa_snapshot[23][27] , \sa_snapshot[23].f.lower[27] );
tran (\sa_snapshot[23][26] , \sa_snapshot[23].r.part0[26] );
tran (\sa_snapshot[23][26] , \sa_snapshot[23].f.lower[26] );
tran (\sa_snapshot[23][25] , \sa_snapshot[23].r.part0[25] );
tran (\sa_snapshot[23][25] , \sa_snapshot[23].f.lower[25] );
tran (\sa_snapshot[23][24] , \sa_snapshot[23].r.part0[24] );
tran (\sa_snapshot[23][24] , \sa_snapshot[23].f.lower[24] );
tran (\sa_snapshot[23][23] , \sa_snapshot[23].r.part0[23] );
tran (\sa_snapshot[23][23] , \sa_snapshot[23].f.lower[23] );
tran (\sa_snapshot[23][22] , \sa_snapshot[23].r.part0[22] );
tran (\sa_snapshot[23][22] , \sa_snapshot[23].f.lower[22] );
tran (\sa_snapshot[23][21] , \sa_snapshot[23].r.part0[21] );
tran (\sa_snapshot[23][21] , \sa_snapshot[23].f.lower[21] );
tran (\sa_snapshot[23][20] , \sa_snapshot[23].r.part0[20] );
tran (\sa_snapshot[23][20] , \sa_snapshot[23].f.lower[20] );
tran (\sa_snapshot[23][19] , \sa_snapshot[23].r.part0[19] );
tran (\sa_snapshot[23][19] , \sa_snapshot[23].f.lower[19] );
tran (\sa_snapshot[23][18] , \sa_snapshot[23].r.part0[18] );
tran (\sa_snapshot[23][18] , \sa_snapshot[23].f.lower[18] );
tran (\sa_snapshot[23][17] , \sa_snapshot[23].r.part0[17] );
tran (\sa_snapshot[23][17] , \sa_snapshot[23].f.lower[17] );
tran (\sa_snapshot[23][16] , \sa_snapshot[23].r.part0[16] );
tran (\sa_snapshot[23][16] , \sa_snapshot[23].f.lower[16] );
tran (\sa_snapshot[23][15] , \sa_snapshot[23].r.part0[15] );
tran (\sa_snapshot[23][15] , \sa_snapshot[23].f.lower[15] );
tran (\sa_snapshot[23][14] , \sa_snapshot[23].r.part0[14] );
tran (\sa_snapshot[23][14] , \sa_snapshot[23].f.lower[14] );
tran (\sa_snapshot[23][13] , \sa_snapshot[23].r.part0[13] );
tran (\sa_snapshot[23][13] , \sa_snapshot[23].f.lower[13] );
tran (\sa_snapshot[23][12] , \sa_snapshot[23].r.part0[12] );
tran (\sa_snapshot[23][12] , \sa_snapshot[23].f.lower[12] );
tran (\sa_snapshot[23][11] , \sa_snapshot[23].r.part0[11] );
tran (\sa_snapshot[23][11] , \sa_snapshot[23].f.lower[11] );
tran (\sa_snapshot[23][10] , \sa_snapshot[23].r.part0[10] );
tran (\sa_snapshot[23][10] , \sa_snapshot[23].f.lower[10] );
tran (\sa_snapshot[23][9] , \sa_snapshot[23].r.part0[9] );
tran (\sa_snapshot[23][9] , \sa_snapshot[23].f.lower[9] );
tran (\sa_snapshot[23][8] , \sa_snapshot[23].r.part0[8] );
tran (\sa_snapshot[23][8] , \sa_snapshot[23].f.lower[8] );
tran (\sa_snapshot[23][7] , \sa_snapshot[23].r.part0[7] );
tran (\sa_snapshot[23][7] , \sa_snapshot[23].f.lower[7] );
tran (\sa_snapshot[23][6] , \sa_snapshot[23].r.part0[6] );
tran (\sa_snapshot[23][6] , \sa_snapshot[23].f.lower[6] );
tran (\sa_snapshot[23][5] , \sa_snapshot[23].r.part0[5] );
tran (\sa_snapshot[23][5] , \sa_snapshot[23].f.lower[5] );
tran (\sa_snapshot[23][4] , \sa_snapshot[23].r.part0[4] );
tran (\sa_snapshot[23][4] , \sa_snapshot[23].f.lower[4] );
tran (\sa_snapshot[23][3] , \sa_snapshot[23].r.part0[3] );
tran (\sa_snapshot[23][3] , \sa_snapshot[23].f.lower[3] );
tran (\sa_snapshot[23][2] , \sa_snapshot[23].r.part0[2] );
tran (\sa_snapshot[23][2] , \sa_snapshot[23].f.lower[2] );
tran (\sa_snapshot[23][1] , \sa_snapshot[23].r.part0[1] );
tran (\sa_snapshot[23][1] , \sa_snapshot[23].f.lower[1] );
tran (\sa_snapshot[23][0] , \sa_snapshot[23].r.part0[0] );
tran (\sa_snapshot[23][0] , \sa_snapshot[23].f.lower[0] );
tran (\sa_snapshot[22][63] , \sa_snapshot[22].r.part1[31] );
tran (\sa_snapshot[22][63] , \sa_snapshot[22].f.unused[13] );
tran (\sa_snapshot[22][62] , \sa_snapshot[22].r.part1[30] );
tran (\sa_snapshot[22][62] , \sa_snapshot[22].f.unused[12] );
tran (\sa_snapshot[22][61] , \sa_snapshot[22].r.part1[29] );
tran (\sa_snapshot[22][61] , \sa_snapshot[22].f.unused[11] );
tran (\sa_snapshot[22][60] , \sa_snapshot[22].r.part1[28] );
tran (\sa_snapshot[22][60] , \sa_snapshot[22].f.unused[10] );
tran (\sa_snapshot[22][59] , \sa_snapshot[22].r.part1[27] );
tran (\sa_snapshot[22][59] , \sa_snapshot[22].f.unused[9] );
tran (\sa_snapshot[22][58] , \sa_snapshot[22].r.part1[26] );
tran (\sa_snapshot[22][58] , \sa_snapshot[22].f.unused[8] );
tran (\sa_snapshot[22][57] , \sa_snapshot[22].r.part1[25] );
tran (\sa_snapshot[22][57] , \sa_snapshot[22].f.unused[7] );
tran (\sa_snapshot[22][56] , \sa_snapshot[22].r.part1[24] );
tran (\sa_snapshot[22][56] , \sa_snapshot[22].f.unused[6] );
tran (\sa_snapshot[22][55] , \sa_snapshot[22].r.part1[23] );
tran (\sa_snapshot[22][55] , \sa_snapshot[22].f.unused[5] );
tran (\sa_snapshot[22][54] , \sa_snapshot[22].r.part1[22] );
tran (\sa_snapshot[22][54] , \sa_snapshot[22].f.unused[4] );
tran (\sa_snapshot[22][53] , \sa_snapshot[22].r.part1[21] );
tran (\sa_snapshot[22][53] , \sa_snapshot[22].f.unused[3] );
tran (\sa_snapshot[22][52] , \sa_snapshot[22].r.part1[20] );
tran (\sa_snapshot[22][52] , \sa_snapshot[22].f.unused[2] );
tran (\sa_snapshot[22][51] , \sa_snapshot[22].r.part1[19] );
tran (\sa_snapshot[22][51] , \sa_snapshot[22].f.unused[1] );
tran (\sa_snapshot[22][50] , \sa_snapshot[22].r.part1[18] );
tran (\sa_snapshot[22][50] , \sa_snapshot[22].f.unused[0] );
tran (\sa_snapshot[22][49] , \sa_snapshot[22].r.part1[17] );
tran (\sa_snapshot[22][49] , \sa_snapshot[22].f.upper[17] );
tran (\sa_snapshot[22][48] , \sa_snapshot[22].r.part1[16] );
tran (\sa_snapshot[22][48] , \sa_snapshot[22].f.upper[16] );
tran (\sa_snapshot[22][47] , \sa_snapshot[22].r.part1[15] );
tran (\sa_snapshot[22][47] , \sa_snapshot[22].f.upper[15] );
tran (\sa_snapshot[22][46] , \sa_snapshot[22].r.part1[14] );
tran (\sa_snapshot[22][46] , \sa_snapshot[22].f.upper[14] );
tran (\sa_snapshot[22][45] , \sa_snapshot[22].r.part1[13] );
tran (\sa_snapshot[22][45] , \sa_snapshot[22].f.upper[13] );
tran (\sa_snapshot[22][44] , \sa_snapshot[22].r.part1[12] );
tran (\sa_snapshot[22][44] , \sa_snapshot[22].f.upper[12] );
tran (\sa_snapshot[22][43] , \sa_snapshot[22].r.part1[11] );
tran (\sa_snapshot[22][43] , \sa_snapshot[22].f.upper[11] );
tran (\sa_snapshot[22][42] , \sa_snapshot[22].r.part1[10] );
tran (\sa_snapshot[22][42] , \sa_snapshot[22].f.upper[10] );
tran (\sa_snapshot[22][41] , \sa_snapshot[22].r.part1[9] );
tran (\sa_snapshot[22][41] , \sa_snapshot[22].f.upper[9] );
tran (\sa_snapshot[22][40] , \sa_snapshot[22].r.part1[8] );
tran (\sa_snapshot[22][40] , \sa_snapshot[22].f.upper[8] );
tran (\sa_snapshot[22][39] , \sa_snapshot[22].r.part1[7] );
tran (\sa_snapshot[22][39] , \sa_snapshot[22].f.upper[7] );
tran (\sa_snapshot[22][38] , \sa_snapshot[22].r.part1[6] );
tran (\sa_snapshot[22][38] , \sa_snapshot[22].f.upper[6] );
tran (\sa_snapshot[22][37] , \sa_snapshot[22].r.part1[5] );
tran (\sa_snapshot[22][37] , \sa_snapshot[22].f.upper[5] );
tran (\sa_snapshot[22][36] , \sa_snapshot[22].r.part1[4] );
tran (\sa_snapshot[22][36] , \sa_snapshot[22].f.upper[4] );
tran (\sa_snapshot[22][35] , \sa_snapshot[22].r.part1[3] );
tran (\sa_snapshot[22][35] , \sa_snapshot[22].f.upper[3] );
tran (\sa_snapshot[22][34] , \sa_snapshot[22].r.part1[2] );
tran (\sa_snapshot[22][34] , \sa_snapshot[22].f.upper[2] );
tran (\sa_snapshot[22][33] , \sa_snapshot[22].r.part1[1] );
tran (\sa_snapshot[22][33] , \sa_snapshot[22].f.upper[1] );
tran (\sa_snapshot[22][32] , \sa_snapshot[22].r.part1[0] );
tran (\sa_snapshot[22][32] , \sa_snapshot[22].f.upper[0] );
tran (\sa_snapshot[22][31] , \sa_snapshot[22].r.part0[31] );
tran (\sa_snapshot[22][31] , \sa_snapshot[22].f.lower[31] );
tran (\sa_snapshot[22][30] , \sa_snapshot[22].r.part0[30] );
tran (\sa_snapshot[22][30] , \sa_snapshot[22].f.lower[30] );
tran (\sa_snapshot[22][29] , \sa_snapshot[22].r.part0[29] );
tran (\sa_snapshot[22][29] , \sa_snapshot[22].f.lower[29] );
tran (\sa_snapshot[22][28] , \sa_snapshot[22].r.part0[28] );
tran (\sa_snapshot[22][28] , \sa_snapshot[22].f.lower[28] );
tran (\sa_snapshot[22][27] , \sa_snapshot[22].r.part0[27] );
tran (\sa_snapshot[22][27] , \sa_snapshot[22].f.lower[27] );
tran (\sa_snapshot[22][26] , \sa_snapshot[22].r.part0[26] );
tran (\sa_snapshot[22][26] , \sa_snapshot[22].f.lower[26] );
tran (\sa_snapshot[22][25] , \sa_snapshot[22].r.part0[25] );
tran (\sa_snapshot[22][25] , \sa_snapshot[22].f.lower[25] );
tran (\sa_snapshot[22][24] , \sa_snapshot[22].r.part0[24] );
tran (\sa_snapshot[22][24] , \sa_snapshot[22].f.lower[24] );
tran (\sa_snapshot[22][23] , \sa_snapshot[22].r.part0[23] );
tran (\sa_snapshot[22][23] , \sa_snapshot[22].f.lower[23] );
tran (\sa_snapshot[22][22] , \sa_snapshot[22].r.part0[22] );
tran (\sa_snapshot[22][22] , \sa_snapshot[22].f.lower[22] );
tran (\sa_snapshot[22][21] , \sa_snapshot[22].r.part0[21] );
tran (\sa_snapshot[22][21] , \sa_snapshot[22].f.lower[21] );
tran (\sa_snapshot[22][20] , \sa_snapshot[22].r.part0[20] );
tran (\sa_snapshot[22][20] , \sa_snapshot[22].f.lower[20] );
tran (\sa_snapshot[22][19] , \sa_snapshot[22].r.part0[19] );
tran (\sa_snapshot[22][19] , \sa_snapshot[22].f.lower[19] );
tran (\sa_snapshot[22][18] , \sa_snapshot[22].r.part0[18] );
tran (\sa_snapshot[22][18] , \sa_snapshot[22].f.lower[18] );
tran (\sa_snapshot[22][17] , \sa_snapshot[22].r.part0[17] );
tran (\sa_snapshot[22][17] , \sa_snapshot[22].f.lower[17] );
tran (\sa_snapshot[22][16] , \sa_snapshot[22].r.part0[16] );
tran (\sa_snapshot[22][16] , \sa_snapshot[22].f.lower[16] );
tran (\sa_snapshot[22][15] , \sa_snapshot[22].r.part0[15] );
tran (\sa_snapshot[22][15] , \sa_snapshot[22].f.lower[15] );
tran (\sa_snapshot[22][14] , \sa_snapshot[22].r.part0[14] );
tran (\sa_snapshot[22][14] , \sa_snapshot[22].f.lower[14] );
tran (\sa_snapshot[22][13] , \sa_snapshot[22].r.part0[13] );
tran (\sa_snapshot[22][13] , \sa_snapshot[22].f.lower[13] );
tran (\sa_snapshot[22][12] , \sa_snapshot[22].r.part0[12] );
tran (\sa_snapshot[22][12] , \sa_snapshot[22].f.lower[12] );
tran (\sa_snapshot[22][11] , \sa_snapshot[22].r.part0[11] );
tran (\sa_snapshot[22][11] , \sa_snapshot[22].f.lower[11] );
tran (\sa_snapshot[22][10] , \sa_snapshot[22].r.part0[10] );
tran (\sa_snapshot[22][10] , \sa_snapshot[22].f.lower[10] );
tran (\sa_snapshot[22][9] , \sa_snapshot[22].r.part0[9] );
tran (\sa_snapshot[22][9] , \sa_snapshot[22].f.lower[9] );
tran (\sa_snapshot[22][8] , \sa_snapshot[22].r.part0[8] );
tran (\sa_snapshot[22][8] , \sa_snapshot[22].f.lower[8] );
tran (\sa_snapshot[22][7] , \sa_snapshot[22].r.part0[7] );
tran (\sa_snapshot[22][7] , \sa_snapshot[22].f.lower[7] );
tran (\sa_snapshot[22][6] , \sa_snapshot[22].r.part0[6] );
tran (\sa_snapshot[22][6] , \sa_snapshot[22].f.lower[6] );
tran (\sa_snapshot[22][5] , \sa_snapshot[22].r.part0[5] );
tran (\sa_snapshot[22][5] , \sa_snapshot[22].f.lower[5] );
tran (\sa_snapshot[22][4] , \sa_snapshot[22].r.part0[4] );
tran (\sa_snapshot[22][4] , \sa_snapshot[22].f.lower[4] );
tran (\sa_snapshot[22][3] , \sa_snapshot[22].r.part0[3] );
tran (\sa_snapshot[22][3] , \sa_snapshot[22].f.lower[3] );
tran (\sa_snapshot[22][2] , \sa_snapshot[22].r.part0[2] );
tran (\sa_snapshot[22][2] , \sa_snapshot[22].f.lower[2] );
tran (\sa_snapshot[22][1] , \sa_snapshot[22].r.part0[1] );
tran (\sa_snapshot[22][1] , \sa_snapshot[22].f.lower[1] );
tran (\sa_snapshot[22][0] , \sa_snapshot[22].r.part0[0] );
tran (\sa_snapshot[22][0] , \sa_snapshot[22].f.lower[0] );
tran (\sa_snapshot[21][63] , \sa_snapshot[21].r.part1[31] );
tran (\sa_snapshot[21][63] , \sa_snapshot[21].f.unused[13] );
tran (\sa_snapshot[21][62] , \sa_snapshot[21].r.part1[30] );
tran (\sa_snapshot[21][62] , \sa_snapshot[21].f.unused[12] );
tran (\sa_snapshot[21][61] , \sa_snapshot[21].r.part1[29] );
tran (\sa_snapshot[21][61] , \sa_snapshot[21].f.unused[11] );
tran (\sa_snapshot[21][60] , \sa_snapshot[21].r.part1[28] );
tran (\sa_snapshot[21][60] , \sa_snapshot[21].f.unused[10] );
tran (\sa_snapshot[21][59] , \sa_snapshot[21].r.part1[27] );
tran (\sa_snapshot[21][59] , \sa_snapshot[21].f.unused[9] );
tran (\sa_snapshot[21][58] , \sa_snapshot[21].r.part1[26] );
tran (\sa_snapshot[21][58] , \sa_snapshot[21].f.unused[8] );
tran (\sa_snapshot[21][57] , \sa_snapshot[21].r.part1[25] );
tran (\sa_snapshot[21][57] , \sa_snapshot[21].f.unused[7] );
tran (\sa_snapshot[21][56] , \sa_snapshot[21].r.part1[24] );
tran (\sa_snapshot[21][56] , \sa_snapshot[21].f.unused[6] );
tran (\sa_snapshot[21][55] , \sa_snapshot[21].r.part1[23] );
tran (\sa_snapshot[21][55] , \sa_snapshot[21].f.unused[5] );
tran (\sa_snapshot[21][54] , \sa_snapshot[21].r.part1[22] );
tran (\sa_snapshot[21][54] , \sa_snapshot[21].f.unused[4] );
tran (\sa_snapshot[21][53] , \sa_snapshot[21].r.part1[21] );
tran (\sa_snapshot[21][53] , \sa_snapshot[21].f.unused[3] );
tran (\sa_snapshot[21][52] , \sa_snapshot[21].r.part1[20] );
tran (\sa_snapshot[21][52] , \sa_snapshot[21].f.unused[2] );
tran (\sa_snapshot[21][51] , \sa_snapshot[21].r.part1[19] );
tran (\sa_snapshot[21][51] , \sa_snapshot[21].f.unused[1] );
tran (\sa_snapshot[21][50] , \sa_snapshot[21].r.part1[18] );
tran (\sa_snapshot[21][50] , \sa_snapshot[21].f.unused[0] );
tran (\sa_snapshot[21][49] , \sa_snapshot[21].r.part1[17] );
tran (\sa_snapshot[21][49] , \sa_snapshot[21].f.upper[17] );
tran (\sa_snapshot[21][48] , \sa_snapshot[21].r.part1[16] );
tran (\sa_snapshot[21][48] , \sa_snapshot[21].f.upper[16] );
tran (\sa_snapshot[21][47] , \sa_snapshot[21].r.part1[15] );
tran (\sa_snapshot[21][47] , \sa_snapshot[21].f.upper[15] );
tran (\sa_snapshot[21][46] , \sa_snapshot[21].r.part1[14] );
tran (\sa_snapshot[21][46] , \sa_snapshot[21].f.upper[14] );
tran (\sa_snapshot[21][45] , \sa_snapshot[21].r.part1[13] );
tran (\sa_snapshot[21][45] , \sa_snapshot[21].f.upper[13] );
tran (\sa_snapshot[21][44] , \sa_snapshot[21].r.part1[12] );
tran (\sa_snapshot[21][44] , \sa_snapshot[21].f.upper[12] );
tran (\sa_snapshot[21][43] , \sa_snapshot[21].r.part1[11] );
tran (\sa_snapshot[21][43] , \sa_snapshot[21].f.upper[11] );
tran (\sa_snapshot[21][42] , \sa_snapshot[21].r.part1[10] );
tran (\sa_snapshot[21][42] , \sa_snapshot[21].f.upper[10] );
tran (\sa_snapshot[21][41] , \sa_snapshot[21].r.part1[9] );
tran (\sa_snapshot[21][41] , \sa_snapshot[21].f.upper[9] );
tran (\sa_snapshot[21][40] , \sa_snapshot[21].r.part1[8] );
tran (\sa_snapshot[21][40] , \sa_snapshot[21].f.upper[8] );
tran (\sa_snapshot[21][39] , \sa_snapshot[21].r.part1[7] );
tran (\sa_snapshot[21][39] , \sa_snapshot[21].f.upper[7] );
tran (\sa_snapshot[21][38] , \sa_snapshot[21].r.part1[6] );
tran (\sa_snapshot[21][38] , \sa_snapshot[21].f.upper[6] );
tran (\sa_snapshot[21][37] , \sa_snapshot[21].r.part1[5] );
tran (\sa_snapshot[21][37] , \sa_snapshot[21].f.upper[5] );
tran (\sa_snapshot[21][36] , \sa_snapshot[21].r.part1[4] );
tran (\sa_snapshot[21][36] , \sa_snapshot[21].f.upper[4] );
tran (\sa_snapshot[21][35] , \sa_snapshot[21].r.part1[3] );
tran (\sa_snapshot[21][35] , \sa_snapshot[21].f.upper[3] );
tran (\sa_snapshot[21][34] , \sa_snapshot[21].r.part1[2] );
tran (\sa_snapshot[21][34] , \sa_snapshot[21].f.upper[2] );
tran (\sa_snapshot[21][33] , \sa_snapshot[21].r.part1[1] );
tran (\sa_snapshot[21][33] , \sa_snapshot[21].f.upper[1] );
tran (\sa_snapshot[21][32] , \sa_snapshot[21].r.part1[0] );
tran (\sa_snapshot[21][32] , \sa_snapshot[21].f.upper[0] );
tran (\sa_snapshot[21][31] , \sa_snapshot[21].r.part0[31] );
tran (\sa_snapshot[21][31] , \sa_snapshot[21].f.lower[31] );
tran (\sa_snapshot[21][30] , \sa_snapshot[21].r.part0[30] );
tran (\sa_snapshot[21][30] , \sa_snapshot[21].f.lower[30] );
tran (\sa_snapshot[21][29] , \sa_snapshot[21].r.part0[29] );
tran (\sa_snapshot[21][29] , \sa_snapshot[21].f.lower[29] );
tran (\sa_snapshot[21][28] , \sa_snapshot[21].r.part0[28] );
tran (\sa_snapshot[21][28] , \sa_snapshot[21].f.lower[28] );
tran (\sa_snapshot[21][27] , \sa_snapshot[21].r.part0[27] );
tran (\sa_snapshot[21][27] , \sa_snapshot[21].f.lower[27] );
tran (\sa_snapshot[21][26] , \sa_snapshot[21].r.part0[26] );
tran (\sa_snapshot[21][26] , \sa_snapshot[21].f.lower[26] );
tran (\sa_snapshot[21][25] , \sa_snapshot[21].r.part0[25] );
tran (\sa_snapshot[21][25] , \sa_snapshot[21].f.lower[25] );
tran (\sa_snapshot[21][24] , \sa_snapshot[21].r.part0[24] );
tran (\sa_snapshot[21][24] , \sa_snapshot[21].f.lower[24] );
tran (\sa_snapshot[21][23] , \sa_snapshot[21].r.part0[23] );
tran (\sa_snapshot[21][23] , \sa_snapshot[21].f.lower[23] );
tran (\sa_snapshot[21][22] , \sa_snapshot[21].r.part0[22] );
tran (\sa_snapshot[21][22] , \sa_snapshot[21].f.lower[22] );
tran (\sa_snapshot[21][21] , \sa_snapshot[21].r.part0[21] );
tran (\sa_snapshot[21][21] , \sa_snapshot[21].f.lower[21] );
tran (\sa_snapshot[21][20] , \sa_snapshot[21].r.part0[20] );
tran (\sa_snapshot[21][20] , \sa_snapshot[21].f.lower[20] );
tran (\sa_snapshot[21][19] , \sa_snapshot[21].r.part0[19] );
tran (\sa_snapshot[21][19] , \sa_snapshot[21].f.lower[19] );
tran (\sa_snapshot[21][18] , \sa_snapshot[21].r.part0[18] );
tran (\sa_snapshot[21][18] , \sa_snapshot[21].f.lower[18] );
tran (\sa_snapshot[21][17] , \sa_snapshot[21].r.part0[17] );
tran (\sa_snapshot[21][17] , \sa_snapshot[21].f.lower[17] );
tran (\sa_snapshot[21][16] , \sa_snapshot[21].r.part0[16] );
tran (\sa_snapshot[21][16] , \sa_snapshot[21].f.lower[16] );
tran (\sa_snapshot[21][15] , \sa_snapshot[21].r.part0[15] );
tran (\sa_snapshot[21][15] , \sa_snapshot[21].f.lower[15] );
tran (\sa_snapshot[21][14] , \sa_snapshot[21].r.part0[14] );
tran (\sa_snapshot[21][14] , \sa_snapshot[21].f.lower[14] );
tran (\sa_snapshot[21][13] , \sa_snapshot[21].r.part0[13] );
tran (\sa_snapshot[21][13] , \sa_snapshot[21].f.lower[13] );
tran (\sa_snapshot[21][12] , \sa_snapshot[21].r.part0[12] );
tran (\sa_snapshot[21][12] , \sa_snapshot[21].f.lower[12] );
tran (\sa_snapshot[21][11] , \sa_snapshot[21].r.part0[11] );
tran (\sa_snapshot[21][11] , \sa_snapshot[21].f.lower[11] );
tran (\sa_snapshot[21][10] , \sa_snapshot[21].r.part0[10] );
tran (\sa_snapshot[21][10] , \sa_snapshot[21].f.lower[10] );
tran (\sa_snapshot[21][9] , \sa_snapshot[21].r.part0[9] );
tran (\sa_snapshot[21][9] , \sa_snapshot[21].f.lower[9] );
tran (\sa_snapshot[21][8] , \sa_snapshot[21].r.part0[8] );
tran (\sa_snapshot[21][8] , \sa_snapshot[21].f.lower[8] );
tran (\sa_snapshot[21][7] , \sa_snapshot[21].r.part0[7] );
tran (\sa_snapshot[21][7] , \sa_snapshot[21].f.lower[7] );
tran (\sa_snapshot[21][6] , \sa_snapshot[21].r.part0[6] );
tran (\sa_snapshot[21][6] , \sa_snapshot[21].f.lower[6] );
tran (\sa_snapshot[21][5] , \sa_snapshot[21].r.part0[5] );
tran (\sa_snapshot[21][5] , \sa_snapshot[21].f.lower[5] );
tran (\sa_snapshot[21][4] , \sa_snapshot[21].r.part0[4] );
tran (\sa_snapshot[21][4] , \sa_snapshot[21].f.lower[4] );
tran (\sa_snapshot[21][3] , \sa_snapshot[21].r.part0[3] );
tran (\sa_snapshot[21][3] , \sa_snapshot[21].f.lower[3] );
tran (\sa_snapshot[21][2] , \sa_snapshot[21].r.part0[2] );
tran (\sa_snapshot[21][2] , \sa_snapshot[21].f.lower[2] );
tran (\sa_snapshot[21][1] , \sa_snapshot[21].r.part0[1] );
tran (\sa_snapshot[21][1] , \sa_snapshot[21].f.lower[1] );
tran (\sa_snapshot[21][0] , \sa_snapshot[21].r.part0[0] );
tran (\sa_snapshot[21][0] , \sa_snapshot[21].f.lower[0] );
tran (\sa_snapshot[20][63] , \sa_snapshot[20].r.part1[31] );
tran (\sa_snapshot[20][63] , \sa_snapshot[20].f.unused[13] );
tran (\sa_snapshot[20][62] , \sa_snapshot[20].r.part1[30] );
tran (\sa_snapshot[20][62] , \sa_snapshot[20].f.unused[12] );
tran (\sa_snapshot[20][61] , \sa_snapshot[20].r.part1[29] );
tran (\sa_snapshot[20][61] , \sa_snapshot[20].f.unused[11] );
tran (\sa_snapshot[20][60] , \sa_snapshot[20].r.part1[28] );
tran (\sa_snapshot[20][60] , \sa_snapshot[20].f.unused[10] );
tran (\sa_snapshot[20][59] , \sa_snapshot[20].r.part1[27] );
tran (\sa_snapshot[20][59] , \sa_snapshot[20].f.unused[9] );
tran (\sa_snapshot[20][58] , \sa_snapshot[20].r.part1[26] );
tran (\sa_snapshot[20][58] , \sa_snapshot[20].f.unused[8] );
tran (\sa_snapshot[20][57] , \sa_snapshot[20].r.part1[25] );
tran (\sa_snapshot[20][57] , \sa_snapshot[20].f.unused[7] );
tran (\sa_snapshot[20][56] , \sa_snapshot[20].r.part1[24] );
tran (\sa_snapshot[20][56] , \sa_snapshot[20].f.unused[6] );
tran (\sa_snapshot[20][55] , \sa_snapshot[20].r.part1[23] );
tran (\sa_snapshot[20][55] , \sa_snapshot[20].f.unused[5] );
tran (\sa_snapshot[20][54] , \sa_snapshot[20].r.part1[22] );
tran (\sa_snapshot[20][54] , \sa_snapshot[20].f.unused[4] );
tran (\sa_snapshot[20][53] , \sa_snapshot[20].r.part1[21] );
tran (\sa_snapshot[20][53] , \sa_snapshot[20].f.unused[3] );
tran (\sa_snapshot[20][52] , \sa_snapshot[20].r.part1[20] );
tran (\sa_snapshot[20][52] , \sa_snapshot[20].f.unused[2] );
tran (\sa_snapshot[20][51] , \sa_snapshot[20].r.part1[19] );
tran (\sa_snapshot[20][51] , \sa_snapshot[20].f.unused[1] );
tran (\sa_snapshot[20][50] , \sa_snapshot[20].r.part1[18] );
tran (\sa_snapshot[20][50] , \sa_snapshot[20].f.unused[0] );
tran (\sa_snapshot[20][49] , \sa_snapshot[20].r.part1[17] );
tran (\sa_snapshot[20][49] , \sa_snapshot[20].f.upper[17] );
tran (\sa_snapshot[20][48] , \sa_snapshot[20].r.part1[16] );
tran (\sa_snapshot[20][48] , \sa_snapshot[20].f.upper[16] );
tran (\sa_snapshot[20][47] , \sa_snapshot[20].r.part1[15] );
tran (\sa_snapshot[20][47] , \sa_snapshot[20].f.upper[15] );
tran (\sa_snapshot[20][46] , \sa_snapshot[20].r.part1[14] );
tran (\sa_snapshot[20][46] , \sa_snapshot[20].f.upper[14] );
tran (\sa_snapshot[20][45] , \sa_snapshot[20].r.part1[13] );
tran (\sa_snapshot[20][45] , \sa_snapshot[20].f.upper[13] );
tran (\sa_snapshot[20][44] , \sa_snapshot[20].r.part1[12] );
tran (\sa_snapshot[20][44] , \sa_snapshot[20].f.upper[12] );
tran (\sa_snapshot[20][43] , \sa_snapshot[20].r.part1[11] );
tran (\sa_snapshot[20][43] , \sa_snapshot[20].f.upper[11] );
tran (\sa_snapshot[20][42] , \sa_snapshot[20].r.part1[10] );
tran (\sa_snapshot[20][42] , \sa_snapshot[20].f.upper[10] );
tran (\sa_snapshot[20][41] , \sa_snapshot[20].r.part1[9] );
tran (\sa_snapshot[20][41] , \sa_snapshot[20].f.upper[9] );
tran (\sa_snapshot[20][40] , \sa_snapshot[20].r.part1[8] );
tran (\sa_snapshot[20][40] , \sa_snapshot[20].f.upper[8] );
tran (\sa_snapshot[20][39] , \sa_snapshot[20].r.part1[7] );
tran (\sa_snapshot[20][39] , \sa_snapshot[20].f.upper[7] );
tran (\sa_snapshot[20][38] , \sa_snapshot[20].r.part1[6] );
tran (\sa_snapshot[20][38] , \sa_snapshot[20].f.upper[6] );
tran (\sa_snapshot[20][37] , \sa_snapshot[20].r.part1[5] );
tran (\sa_snapshot[20][37] , \sa_snapshot[20].f.upper[5] );
tran (\sa_snapshot[20][36] , \sa_snapshot[20].r.part1[4] );
tran (\sa_snapshot[20][36] , \sa_snapshot[20].f.upper[4] );
tran (\sa_snapshot[20][35] , \sa_snapshot[20].r.part1[3] );
tran (\sa_snapshot[20][35] , \sa_snapshot[20].f.upper[3] );
tran (\sa_snapshot[20][34] , \sa_snapshot[20].r.part1[2] );
tran (\sa_snapshot[20][34] , \sa_snapshot[20].f.upper[2] );
tran (\sa_snapshot[20][33] , \sa_snapshot[20].r.part1[1] );
tran (\sa_snapshot[20][33] , \sa_snapshot[20].f.upper[1] );
tran (\sa_snapshot[20][32] , \sa_snapshot[20].r.part1[0] );
tran (\sa_snapshot[20][32] , \sa_snapshot[20].f.upper[0] );
tran (\sa_snapshot[20][31] , \sa_snapshot[20].r.part0[31] );
tran (\sa_snapshot[20][31] , \sa_snapshot[20].f.lower[31] );
tran (\sa_snapshot[20][30] , \sa_snapshot[20].r.part0[30] );
tran (\sa_snapshot[20][30] , \sa_snapshot[20].f.lower[30] );
tran (\sa_snapshot[20][29] , \sa_snapshot[20].r.part0[29] );
tran (\sa_snapshot[20][29] , \sa_snapshot[20].f.lower[29] );
tran (\sa_snapshot[20][28] , \sa_snapshot[20].r.part0[28] );
tran (\sa_snapshot[20][28] , \sa_snapshot[20].f.lower[28] );
tran (\sa_snapshot[20][27] , \sa_snapshot[20].r.part0[27] );
tran (\sa_snapshot[20][27] , \sa_snapshot[20].f.lower[27] );
tran (\sa_snapshot[20][26] , \sa_snapshot[20].r.part0[26] );
tran (\sa_snapshot[20][26] , \sa_snapshot[20].f.lower[26] );
tran (\sa_snapshot[20][25] , \sa_snapshot[20].r.part0[25] );
tran (\sa_snapshot[20][25] , \sa_snapshot[20].f.lower[25] );
tran (\sa_snapshot[20][24] , \sa_snapshot[20].r.part0[24] );
tran (\sa_snapshot[20][24] , \sa_snapshot[20].f.lower[24] );
tran (\sa_snapshot[20][23] , \sa_snapshot[20].r.part0[23] );
tran (\sa_snapshot[20][23] , \sa_snapshot[20].f.lower[23] );
tran (\sa_snapshot[20][22] , \sa_snapshot[20].r.part0[22] );
tran (\sa_snapshot[20][22] , \sa_snapshot[20].f.lower[22] );
tran (\sa_snapshot[20][21] , \sa_snapshot[20].r.part0[21] );
tran (\sa_snapshot[20][21] , \sa_snapshot[20].f.lower[21] );
tran (\sa_snapshot[20][20] , \sa_snapshot[20].r.part0[20] );
tran (\sa_snapshot[20][20] , \sa_snapshot[20].f.lower[20] );
tran (\sa_snapshot[20][19] , \sa_snapshot[20].r.part0[19] );
tran (\sa_snapshot[20][19] , \sa_snapshot[20].f.lower[19] );
tran (\sa_snapshot[20][18] , \sa_snapshot[20].r.part0[18] );
tran (\sa_snapshot[20][18] , \sa_snapshot[20].f.lower[18] );
tran (\sa_snapshot[20][17] , \sa_snapshot[20].r.part0[17] );
tran (\sa_snapshot[20][17] , \sa_snapshot[20].f.lower[17] );
tran (\sa_snapshot[20][16] , \sa_snapshot[20].r.part0[16] );
tran (\sa_snapshot[20][16] , \sa_snapshot[20].f.lower[16] );
tran (\sa_snapshot[20][15] , \sa_snapshot[20].r.part0[15] );
tran (\sa_snapshot[20][15] , \sa_snapshot[20].f.lower[15] );
tran (\sa_snapshot[20][14] , \sa_snapshot[20].r.part0[14] );
tran (\sa_snapshot[20][14] , \sa_snapshot[20].f.lower[14] );
tran (\sa_snapshot[20][13] , \sa_snapshot[20].r.part0[13] );
tran (\sa_snapshot[20][13] , \sa_snapshot[20].f.lower[13] );
tran (\sa_snapshot[20][12] , \sa_snapshot[20].r.part0[12] );
tran (\sa_snapshot[20][12] , \sa_snapshot[20].f.lower[12] );
tran (\sa_snapshot[20][11] , \sa_snapshot[20].r.part0[11] );
tran (\sa_snapshot[20][11] , \sa_snapshot[20].f.lower[11] );
tran (\sa_snapshot[20][10] , \sa_snapshot[20].r.part0[10] );
tran (\sa_snapshot[20][10] , \sa_snapshot[20].f.lower[10] );
tran (\sa_snapshot[20][9] , \sa_snapshot[20].r.part0[9] );
tran (\sa_snapshot[20][9] , \sa_snapshot[20].f.lower[9] );
tran (\sa_snapshot[20][8] , \sa_snapshot[20].r.part0[8] );
tran (\sa_snapshot[20][8] , \sa_snapshot[20].f.lower[8] );
tran (\sa_snapshot[20][7] , \sa_snapshot[20].r.part0[7] );
tran (\sa_snapshot[20][7] , \sa_snapshot[20].f.lower[7] );
tran (\sa_snapshot[20][6] , \sa_snapshot[20].r.part0[6] );
tran (\sa_snapshot[20][6] , \sa_snapshot[20].f.lower[6] );
tran (\sa_snapshot[20][5] , \sa_snapshot[20].r.part0[5] );
tran (\sa_snapshot[20][5] , \sa_snapshot[20].f.lower[5] );
tran (\sa_snapshot[20][4] , \sa_snapshot[20].r.part0[4] );
tran (\sa_snapshot[20][4] , \sa_snapshot[20].f.lower[4] );
tran (\sa_snapshot[20][3] , \sa_snapshot[20].r.part0[3] );
tran (\sa_snapshot[20][3] , \sa_snapshot[20].f.lower[3] );
tran (\sa_snapshot[20][2] , \sa_snapshot[20].r.part0[2] );
tran (\sa_snapshot[20][2] , \sa_snapshot[20].f.lower[2] );
tran (\sa_snapshot[20][1] , \sa_snapshot[20].r.part0[1] );
tran (\sa_snapshot[20][1] , \sa_snapshot[20].f.lower[1] );
tran (\sa_snapshot[20][0] , \sa_snapshot[20].r.part0[0] );
tran (\sa_snapshot[20][0] , \sa_snapshot[20].f.lower[0] );
tran (\sa_snapshot[19][63] , \sa_snapshot[19].r.part1[31] );
tran (\sa_snapshot[19][63] , \sa_snapshot[19].f.unused[13] );
tran (\sa_snapshot[19][62] , \sa_snapshot[19].r.part1[30] );
tran (\sa_snapshot[19][62] , \sa_snapshot[19].f.unused[12] );
tran (\sa_snapshot[19][61] , \sa_snapshot[19].r.part1[29] );
tran (\sa_snapshot[19][61] , \sa_snapshot[19].f.unused[11] );
tran (\sa_snapshot[19][60] , \sa_snapshot[19].r.part1[28] );
tran (\sa_snapshot[19][60] , \sa_snapshot[19].f.unused[10] );
tran (\sa_snapshot[19][59] , \sa_snapshot[19].r.part1[27] );
tran (\sa_snapshot[19][59] , \sa_snapshot[19].f.unused[9] );
tran (\sa_snapshot[19][58] , \sa_snapshot[19].r.part1[26] );
tran (\sa_snapshot[19][58] , \sa_snapshot[19].f.unused[8] );
tran (\sa_snapshot[19][57] , \sa_snapshot[19].r.part1[25] );
tran (\sa_snapshot[19][57] , \sa_snapshot[19].f.unused[7] );
tran (\sa_snapshot[19][56] , \sa_snapshot[19].r.part1[24] );
tran (\sa_snapshot[19][56] , \sa_snapshot[19].f.unused[6] );
tran (\sa_snapshot[19][55] , \sa_snapshot[19].r.part1[23] );
tran (\sa_snapshot[19][55] , \sa_snapshot[19].f.unused[5] );
tran (\sa_snapshot[19][54] , \sa_snapshot[19].r.part1[22] );
tran (\sa_snapshot[19][54] , \sa_snapshot[19].f.unused[4] );
tran (\sa_snapshot[19][53] , \sa_snapshot[19].r.part1[21] );
tran (\sa_snapshot[19][53] , \sa_snapshot[19].f.unused[3] );
tran (\sa_snapshot[19][52] , \sa_snapshot[19].r.part1[20] );
tran (\sa_snapshot[19][52] , \sa_snapshot[19].f.unused[2] );
tran (\sa_snapshot[19][51] , \sa_snapshot[19].r.part1[19] );
tran (\sa_snapshot[19][51] , \sa_snapshot[19].f.unused[1] );
tran (\sa_snapshot[19][50] , \sa_snapshot[19].r.part1[18] );
tran (\sa_snapshot[19][50] , \sa_snapshot[19].f.unused[0] );
tran (\sa_snapshot[19][49] , \sa_snapshot[19].r.part1[17] );
tran (\sa_snapshot[19][49] , \sa_snapshot[19].f.upper[17] );
tran (\sa_snapshot[19][48] , \sa_snapshot[19].r.part1[16] );
tran (\sa_snapshot[19][48] , \sa_snapshot[19].f.upper[16] );
tran (\sa_snapshot[19][47] , \sa_snapshot[19].r.part1[15] );
tran (\sa_snapshot[19][47] , \sa_snapshot[19].f.upper[15] );
tran (\sa_snapshot[19][46] , \sa_snapshot[19].r.part1[14] );
tran (\sa_snapshot[19][46] , \sa_snapshot[19].f.upper[14] );
tran (\sa_snapshot[19][45] , \sa_snapshot[19].r.part1[13] );
tran (\sa_snapshot[19][45] , \sa_snapshot[19].f.upper[13] );
tran (\sa_snapshot[19][44] , \sa_snapshot[19].r.part1[12] );
tran (\sa_snapshot[19][44] , \sa_snapshot[19].f.upper[12] );
tran (\sa_snapshot[19][43] , \sa_snapshot[19].r.part1[11] );
tran (\sa_snapshot[19][43] , \sa_snapshot[19].f.upper[11] );
tran (\sa_snapshot[19][42] , \sa_snapshot[19].r.part1[10] );
tran (\sa_snapshot[19][42] , \sa_snapshot[19].f.upper[10] );
tran (\sa_snapshot[19][41] , \sa_snapshot[19].r.part1[9] );
tran (\sa_snapshot[19][41] , \sa_snapshot[19].f.upper[9] );
tran (\sa_snapshot[19][40] , \sa_snapshot[19].r.part1[8] );
tran (\sa_snapshot[19][40] , \sa_snapshot[19].f.upper[8] );
tran (\sa_snapshot[19][39] , \sa_snapshot[19].r.part1[7] );
tran (\sa_snapshot[19][39] , \sa_snapshot[19].f.upper[7] );
tran (\sa_snapshot[19][38] , \sa_snapshot[19].r.part1[6] );
tran (\sa_snapshot[19][38] , \sa_snapshot[19].f.upper[6] );
tran (\sa_snapshot[19][37] , \sa_snapshot[19].r.part1[5] );
tran (\sa_snapshot[19][37] , \sa_snapshot[19].f.upper[5] );
tran (\sa_snapshot[19][36] , \sa_snapshot[19].r.part1[4] );
tran (\sa_snapshot[19][36] , \sa_snapshot[19].f.upper[4] );
tran (\sa_snapshot[19][35] , \sa_snapshot[19].r.part1[3] );
tran (\sa_snapshot[19][35] , \sa_snapshot[19].f.upper[3] );
tran (\sa_snapshot[19][34] , \sa_snapshot[19].r.part1[2] );
tran (\sa_snapshot[19][34] , \sa_snapshot[19].f.upper[2] );
tran (\sa_snapshot[19][33] , \sa_snapshot[19].r.part1[1] );
tran (\sa_snapshot[19][33] , \sa_snapshot[19].f.upper[1] );
tran (\sa_snapshot[19][32] , \sa_snapshot[19].r.part1[0] );
tran (\sa_snapshot[19][32] , \sa_snapshot[19].f.upper[0] );
tran (\sa_snapshot[19][31] , \sa_snapshot[19].r.part0[31] );
tran (\sa_snapshot[19][31] , \sa_snapshot[19].f.lower[31] );
tran (\sa_snapshot[19][30] , \sa_snapshot[19].r.part0[30] );
tran (\sa_snapshot[19][30] , \sa_snapshot[19].f.lower[30] );
tran (\sa_snapshot[19][29] , \sa_snapshot[19].r.part0[29] );
tran (\sa_snapshot[19][29] , \sa_snapshot[19].f.lower[29] );
tran (\sa_snapshot[19][28] , \sa_snapshot[19].r.part0[28] );
tran (\sa_snapshot[19][28] , \sa_snapshot[19].f.lower[28] );
tran (\sa_snapshot[19][27] , \sa_snapshot[19].r.part0[27] );
tran (\sa_snapshot[19][27] , \sa_snapshot[19].f.lower[27] );
tran (\sa_snapshot[19][26] , \sa_snapshot[19].r.part0[26] );
tran (\sa_snapshot[19][26] , \sa_snapshot[19].f.lower[26] );
tran (\sa_snapshot[19][25] , \sa_snapshot[19].r.part0[25] );
tran (\sa_snapshot[19][25] , \sa_snapshot[19].f.lower[25] );
tran (\sa_snapshot[19][24] , \sa_snapshot[19].r.part0[24] );
tran (\sa_snapshot[19][24] , \sa_snapshot[19].f.lower[24] );
tran (\sa_snapshot[19][23] , \sa_snapshot[19].r.part0[23] );
tran (\sa_snapshot[19][23] , \sa_snapshot[19].f.lower[23] );
tran (\sa_snapshot[19][22] , \sa_snapshot[19].r.part0[22] );
tran (\sa_snapshot[19][22] , \sa_snapshot[19].f.lower[22] );
tran (\sa_snapshot[19][21] , \sa_snapshot[19].r.part0[21] );
tran (\sa_snapshot[19][21] , \sa_snapshot[19].f.lower[21] );
tran (\sa_snapshot[19][20] , \sa_snapshot[19].r.part0[20] );
tran (\sa_snapshot[19][20] , \sa_snapshot[19].f.lower[20] );
tran (\sa_snapshot[19][19] , \sa_snapshot[19].r.part0[19] );
tran (\sa_snapshot[19][19] , \sa_snapshot[19].f.lower[19] );
tran (\sa_snapshot[19][18] , \sa_snapshot[19].r.part0[18] );
tran (\sa_snapshot[19][18] , \sa_snapshot[19].f.lower[18] );
tran (\sa_snapshot[19][17] , \sa_snapshot[19].r.part0[17] );
tran (\sa_snapshot[19][17] , \sa_snapshot[19].f.lower[17] );
tran (\sa_snapshot[19][16] , \sa_snapshot[19].r.part0[16] );
tran (\sa_snapshot[19][16] , \sa_snapshot[19].f.lower[16] );
tran (\sa_snapshot[19][15] , \sa_snapshot[19].r.part0[15] );
tran (\sa_snapshot[19][15] , \sa_snapshot[19].f.lower[15] );
tran (\sa_snapshot[19][14] , \sa_snapshot[19].r.part0[14] );
tran (\sa_snapshot[19][14] , \sa_snapshot[19].f.lower[14] );
tran (\sa_snapshot[19][13] , \sa_snapshot[19].r.part0[13] );
tran (\sa_snapshot[19][13] , \sa_snapshot[19].f.lower[13] );
tran (\sa_snapshot[19][12] , \sa_snapshot[19].r.part0[12] );
tran (\sa_snapshot[19][12] , \sa_snapshot[19].f.lower[12] );
tran (\sa_snapshot[19][11] , \sa_snapshot[19].r.part0[11] );
tran (\sa_snapshot[19][11] , \sa_snapshot[19].f.lower[11] );
tran (\sa_snapshot[19][10] , \sa_snapshot[19].r.part0[10] );
tran (\sa_snapshot[19][10] , \sa_snapshot[19].f.lower[10] );
tran (\sa_snapshot[19][9] , \sa_snapshot[19].r.part0[9] );
tran (\sa_snapshot[19][9] , \sa_snapshot[19].f.lower[9] );
tran (\sa_snapshot[19][8] , \sa_snapshot[19].r.part0[8] );
tran (\sa_snapshot[19][8] , \sa_snapshot[19].f.lower[8] );
tran (\sa_snapshot[19][7] , \sa_snapshot[19].r.part0[7] );
tran (\sa_snapshot[19][7] , \sa_snapshot[19].f.lower[7] );
tran (\sa_snapshot[19][6] , \sa_snapshot[19].r.part0[6] );
tran (\sa_snapshot[19][6] , \sa_snapshot[19].f.lower[6] );
tran (\sa_snapshot[19][5] , \sa_snapshot[19].r.part0[5] );
tran (\sa_snapshot[19][5] , \sa_snapshot[19].f.lower[5] );
tran (\sa_snapshot[19][4] , \sa_snapshot[19].r.part0[4] );
tran (\sa_snapshot[19][4] , \sa_snapshot[19].f.lower[4] );
tran (\sa_snapshot[19][3] , \sa_snapshot[19].r.part0[3] );
tran (\sa_snapshot[19][3] , \sa_snapshot[19].f.lower[3] );
tran (\sa_snapshot[19][2] , \sa_snapshot[19].r.part0[2] );
tran (\sa_snapshot[19][2] , \sa_snapshot[19].f.lower[2] );
tran (\sa_snapshot[19][1] , \sa_snapshot[19].r.part0[1] );
tran (\sa_snapshot[19][1] , \sa_snapshot[19].f.lower[1] );
tran (\sa_snapshot[19][0] , \sa_snapshot[19].r.part0[0] );
tran (\sa_snapshot[19][0] , \sa_snapshot[19].f.lower[0] );
tran (\sa_snapshot[18][63] , \sa_snapshot[18].r.part1[31] );
tran (\sa_snapshot[18][63] , \sa_snapshot[18].f.unused[13] );
tran (\sa_snapshot[18][62] , \sa_snapshot[18].r.part1[30] );
tran (\sa_snapshot[18][62] , \sa_snapshot[18].f.unused[12] );
tran (\sa_snapshot[18][61] , \sa_snapshot[18].r.part1[29] );
tran (\sa_snapshot[18][61] , \sa_snapshot[18].f.unused[11] );
tran (\sa_snapshot[18][60] , \sa_snapshot[18].r.part1[28] );
tran (\sa_snapshot[18][60] , \sa_snapshot[18].f.unused[10] );
tran (\sa_snapshot[18][59] , \sa_snapshot[18].r.part1[27] );
tran (\sa_snapshot[18][59] , \sa_snapshot[18].f.unused[9] );
tran (\sa_snapshot[18][58] , \sa_snapshot[18].r.part1[26] );
tran (\sa_snapshot[18][58] , \sa_snapshot[18].f.unused[8] );
tran (\sa_snapshot[18][57] , \sa_snapshot[18].r.part1[25] );
tran (\sa_snapshot[18][57] , \sa_snapshot[18].f.unused[7] );
tran (\sa_snapshot[18][56] , \sa_snapshot[18].r.part1[24] );
tran (\sa_snapshot[18][56] , \sa_snapshot[18].f.unused[6] );
tran (\sa_snapshot[18][55] , \sa_snapshot[18].r.part1[23] );
tran (\sa_snapshot[18][55] , \sa_snapshot[18].f.unused[5] );
tran (\sa_snapshot[18][54] , \sa_snapshot[18].r.part1[22] );
tran (\sa_snapshot[18][54] , \sa_snapshot[18].f.unused[4] );
tran (\sa_snapshot[18][53] , \sa_snapshot[18].r.part1[21] );
tran (\sa_snapshot[18][53] , \sa_snapshot[18].f.unused[3] );
tran (\sa_snapshot[18][52] , \sa_snapshot[18].r.part1[20] );
tran (\sa_snapshot[18][52] , \sa_snapshot[18].f.unused[2] );
tran (\sa_snapshot[18][51] , \sa_snapshot[18].r.part1[19] );
tran (\sa_snapshot[18][51] , \sa_snapshot[18].f.unused[1] );
tran (\sa_snapshot[18][50] , \sa_snapshot[18].r.part1[18] );
tran (\sa_snapshot[18][50] , \sa_snapshot[18].f.unused[0] );
tran (\sa_snapshot[18][49] , \sa_snapshot[18].r.part1[17] );
tran (\sa_snapshot[18][49] , \sa_snapshot[18].f.upper[17] );
tran (\sa_snapshot[18][48] , \sa_snapshot[18].r.part1[16] );
tran (\sa_snapshot[18][48] , \sa_snapshot[18].f.upper[16] );
tran (\sa_snapshot[18][47] , \sa_snapshot[18].r.part1[15] );
tran (\sa_snapshot[18][47] , \sa_snapshot[18].f.upper[15] );
tran (\sa_snapshot[18][46] , \sa_snapshot[18].r.part1[14] );
tran (\sa_snapshot[18][46] , \sa_snapshot[18].f.upper[14] );
tran (\sa_snapshot[18][45] , \sa_snapshot[18].r.part1[13] );
tran (\sa_snapshot[18][45] , \sa_snapshot[18].f.upper[13] );
tran (\sa_snapshot[18][44] , \sa_snapshot[18].r.part1[12] );
tran (\sa_snapshot[18][44] , \sa_snapshot[18].f.upper[12] );
tran (\sa_snapshot[18][43] , \sa_snapshot[18].r.part1[11] );
tran (\sa_snapshot[18][43] , \sa_snapshot[18].f.upper[11] );
tran (\sa_snapshot[18][42] , \sa_snapshot[18].r.part1[10] );
tran (\sa_snapshot[18][42] , \sa_snapshot[18].f.upper[10] );
tran (\sa_snapshot[18][41] , \sa_snapshot[18].r.part1[9] );
tran (\sa_snapshot[18][41] , \sa_snapshot[18].f.upper[9] );
tran (\sa_snapshot[18][40] , \sa_snapshot[18].r.part1[8] );
tran (\sa_snapshot[18][40] , \sa_snapshot[18].f.upper[8] );
tran (\sa_snapshot[18][39] , \sa_snapshot[18].r.part1[7] );
tran (\sa_snapshot[18][39] , \sa_snapshot[18].f.upper[7] );
tran (\sa_snapshot[18][38] , \sa_snapshot[18].r.part1[6] );
tran (\sa_snapshot[18][38] , \sa_snapshot[18].f.upper[6] );
tran (\sa_snapshot[18][37] , \sa_snapshot[18].r.part1[5] );
tran (\sa_snapshot[18][37] , \sa_snapshot[18].f.upper[5] );
tran (\sa_snapshot[18][36] , \sa_snapshot[18].r.part1[4] );
tran (\sa_snapshot[18][36] , \sa_snapshot[18].f.upper[4] );
tran (\sa_snapshot[18][35] , \sa_snapshot[18].r.part1[3] );
tran (\sa_snapshot[18][35] , \sa_snapshot[18].f.upper[3] );
tran (\sa_snapshot[18][34] , \sa_snapshot[18].r.part1[2] );
tran (\sa_snapshot[18][34] , \sa_snapshot[18].f.upper[2] );
tran (\sa_snapshot[18][33] , \sa_snapshot[18].r.part1[1] );
tran (\sa_snapshot[18][33] , \sa_snapshot[18].f.upper[1] );
tran (\sa_snapshot[18][32] , \sa_snapshot[18].r.part1[0] );
tran (\sa_snapshot[18][32] , \sa_snapshot[18].f.upper[0] );
tran (\sa_snapshot[18][31] , \sa_snapshot[18].r.part0[31] );
tran (\sa_snapshot[18][31] , \sa_snapshot[18].f.lower[31] );
tran (\sa_snapshot[18][30] , \sa_snapshot[18].r.part0[30] );
tran (\sa_snapshot[18][30] , \sa_snapshot[18].f.lower[30] );
tran (\sa_snapshot[18][29] , \sa_snapshot[18].r.part0[29] );
tran (\sa_snapshot[18][29] , \sa_snapshot[18].f.lower[29] );
tran (\sa_snapshot[18][28] , \sa_snapshot[18].r.part0[28] );
tran (\sa_snapshot[18][28] , \sa_snapshot[18].f.lower[28] );
tran (\sa_snapshot[18][27] , \sa_snapshot[18].r.part0[27] );
tran (\sa_snapshot[18][27] , \sa_snapshot[18].f.lower[27] );
tran (\sa_snapshot[18][26] , \sa_snapshot[18].r.part0[26] );
tran (\sa_snapshot[18][26] , \sa_snapshot[18].f.lower[26] );
tran (\sa_snapshot[18][25] , \sa_snapshot[18].r.part0[25] );
tran (\sa_snapshot[18][25] , \sa_snapshot[18].f.lower[25] );
tran (\sa_snapshot[18][24] , \sa_snapshot[18].r.part0[24] );
tran (\sa_snapshot[18][24] , \sa_snapshot[18].f.lower[24] );
tran (\sa_snapshot[18][23] , \sa_snapshot[18].r.part0[23] );
tran (\sa_snapshot[18][23] , \sa_snapshot[18].f.lower[23] );
tran (\sa_snapshot[18][22] , \sa_snapshot[18].r.part0[22] );
tran (\sa_snapshot[18][22] , \sa_snapshot[18].f.lower[22] );
tran (\sa_snapshot[18][21] , \sa_snapshot[18].r.part0[21] );
tran (\sa_snapshot[18][21] , \sa_snapshot[18].f.lower[21] );
tran (\sa_snapshot[18][20] , \sa_snapshot[18].r.part0[20] );
tran (\sa_snapshot[18][20] , \sa_snapshot[18].f.lower[20] );
tran (\sa_snapshot[18][19] , \sa_snapshot[18].r.part0[19] );
tran (\sa_snapshot[18][19] , \sa_snapshot[18].f.lower[19] );
tran (\sa_snapshot[18][18] , \sa_snapshot[18].r.part0[18] );
tran (\sa_snapshot[18][18] , \sa_snapshot[18].f.lower[18] );
tran (\sa_snapshot[18][17] , \sa_snapshot[18].r.part0[17] );
tran (\sa_snapshot[18][17] , \sa_snapshot[18].f.lower[17] );
tran (\sa_snapshot[18][16] , \sa_snapshot[18].r.part0[16] );
tran (\sa_snapshot[18][16] , \sa_snapshot[18].f.lower[16] );
tran (\sa_snapshot[18][15] , \sa_snapshot[18].r.part0[15] );
tran (\sa_snapshot[18][15] , \sa_snapshot[18].f.lower[15] );
tran (\sa_snapshot[18][14] , \sa_snapshot[18].r.part0[14] );
tran (\sa_snapshot[18][14] , \sa_snapshot[18].f.lower[14] );
tran (\sa_snapshot[18][13] , \sa_snapshot[18].r.part0[13] );
tran (\sa_snapshot[18][13] , \sa_snapshot[18].f.lower[13] );
tran (\sa_snapshot[18][12] , \sa_snapshot[18].r.part0[12] );
tran (\sa_snapshot[18][12] , \sa_snapshot[18].f.lower[12] );
tran (\sa_snapshot[18][11] , \sa_snapshot[18].r.part0[11] );
tran (\sa_snapshot[18][11] , \sa_snapshot[18].f.lower[11] );
tran (\sa_snapshot[18][10] , \sa_snapshot[18].r.part0[10] );
tran (\sa_snapshot[18][10] , \sa_snapshot[18].f.lower[10] );
tran (\sa_snapshot[18][9] , \sa_snapshot[18].r.part0[9] );
tran (\sa_snapshot[18][9] , \sa_snapshot[18].f.lower[9] );
tran (\sa_snapshot[18][8] , \sa_snapshot[18].r.part0[8] );
tran (\sa_snapshot[18][8] , \sa_snapshot[18].f.lower[8] );
tran (\sa_snapshot[18][7] , \sa_snapshot[18].r.part0[7] );
tran (\sa_snapshot[18][7] , \sa_snapshot[18].f.lower[7] );
tran (\sa_snapshot[18][6] , \sa_snapshot[18].r.part0[6] );
tran (\sa_snapshot[18][6] , \sa_snapshot[18].f.lower[6] );
tran (\sa_snapshot[18][5] , \sa_snapshot[18].r.part0[5] );
tran (\sa_snapshot[18][5] , \sa_snapshot[18].f.lower[5] );
tran (\sa_snapshot[18][4] , \sa_snapshot[18].r.part0[4] );
tran (\sa_snapshot[18][4] , \sa_snapshot[18].f.lower[4] );
tran (\sa_snapshot[18][3] , \sa_snapshot[18].r.part0[3] );
tran (\sa_snapshot[18][3] , \sa_snapshot[18].f.lower[3] );
tran (\sa_snapshot[18][2] , \sa_snapshot[18].r.part0[2] );
tran (\sa_snapshot[18][2] , \sa_snapshot[18].f.lower[2] );
tran (\sa_snapshot[18][1] , \sa_snapshot[18].r.part0[1] );
tran (\sa_snapshot[18][1] , \sa_snapshot[18].f.lower[1] );
tran (\sa_snapshot[18][0] , \sa_snapshot[18].r.part0[0] );
tran (\sa_snapshot[18][0] , \sa_snapshot[18].f.lower[0] );
tran (\sa_snapshot[17][63] , \sa_snapshot[17].r.part1[31] );
tran (\sa_snapshot[17][63] , \sa_snapshot[17].f.unused[13] );
tran (\sa_snapshot[17][62] , \sa_snapshot[17].r.part1[30] );
tran (\sa_snapshot[17][62] , \sa_snapshot[17].f.unused[12] );
tran (\sa_snapshot[17][61] , \sa_snapshot[17].r.part1[29] );
tran (\sa_snapshot[17][61] , \sa_snapshot[17].f.unused[11] );
tran (\sa_snapshot[17][60] , \sa_snapshot[17].r.part1[28] );
tran (\sa_snapshot[17][60] , \sa_snapshot[17].f.unused[10] );
tran (\sa_snapshot[17][59] , \sa_snapshot[17].r.part1[27] );
tran (\sa_snapshot[17][59] , \sa_snapshot[17].f.unused[9] );
tran (\sa_snapshot[17][58] , \sa_snapshot[17].r.part1[26] );
tran (\sa_snapshot[17][58] , \sa_snapshot[17].f.unused[8] );
tran (\sa_snapshot[17][57] , \sa_snapshot[17].r.part1[25] );
tran (\sa_snapshot[17][57] , \sa_snapshot[17].f.unused[7] );
tran (\sa_snapshot[17][56] , \sa_snapshot[17].r.part1[24] );
tran (\sa_snapshot[17][56] , \sa_snapshot[17].f.unused[6] );
tran (\sa_snapshot[17][55] , \sa_snapshot[17].r.part1[23] );
tran (\sa_snapshot[17][55] , \sa_snapshot[17].f.unused[5] );
tran (\sa_snapshot[17][54] , \sa_snapshot[17].r.part1[22] );
tran (\sa_snapshot[17][54] , \sa_snapshot[17].f.unused[4] );
tran (\sa_snapshot[17][53] , \sa_snapshot[17].r.part1[21] );
tran (\sa_snapshot[17][53] , \sa_snapshot[17].f.unused[3] );
tran (\sa_snapshot[17][52] , \sa_snapshot[17].r.part1[20] );
tran (\sa_snapshot[17][52] , \sa_snapshot[17].f.unused[2] );
tran (\sa_snapshot[17][51] , \sa_snapshot[17].r.part1[19] );
tran (\sa_snapshot[17][51] , \sa_snapshot[17].f.unused[1] );
tran (\sa_snapshot[17][50] , \sa_snapshot[17].r.part1[18] );
tran (\sa_snapshot[17][50] , \sa_snapshot[17].f.unused[0] );
tran (\sa_snapshot[17][49] , \sa_snapshot[17].r.part1[17] );
tran (\sa_snapshot[17][49] , \sa_snapshot[17].f.upper[17] );
tran (\sa_snapshot[17][48] , \sa_snapshot[17].r.part1[16] );
tran (\sa_snapshot[17][48] , \sa_snapshot[17].f.upper[16] );
tran (\sa_snapshot[17][47] , \sa_snapshot[17].r.part1[15] );
tran (\sa_snapshot[17][47] , \sa_snapshot[17].f.upper[15] );
tran (\sa_snapshot[17][46] , \sa_snapshot[17].r.part1[14] );
tran (\sa_snapshot[17][46] , \sa_snapshot[17].f.upper[14] );
tran (\sa_snapshot[17][45] , \sa_snapshot[17].r.part1[13] );
tran (\sa_snapshot[17][45] , \sa_snapshot[17].f.upper[13] );
tran (\sa_snapshot[17][44] , \sa_snapshot[17].r.part1[12] );
tran (\sa_snapshot[17][44] , \sa_snapshot[17].f.upper[12] );
tran (\sa_snapshot[17][43] , \sa_snapshot[17].r.part1[11] );
tran (\sa_snapshot[17][43] , \sa_snapshot[17].f.upper[11] );
tran (\sa_snapshot[17][42] , \sa_snapshot[17].r.part1[10] );
tran (\sa_snapshot[17][42] , \sa_snapshot[17].f.upper[10] );
tran (\sa_snapshot[17][41] , \sa_snapshot[17].r.part1[9] );
tran (\sa_snapshot[17][41] , \sa_snapshot[17].f.upper[9] );
tran (\sa_snapshot[17][40] , \sa_snapshot[17].r.part1[8] );
tran (\sa_snapshot[17][40] , \sa_snapshot[17].f.upper[8] );
tran (\sa_snapshot[17][39] , \sa_snapshot[17].r.part1[7] );
tran (\sa_snapshot[17][39] , \sa_snapshot[17].f.upper[7] );
tran (\sa_snapshot[17][38] , \sa_snapshot[17].r.part1[6] );
tran (\sa_snapshot[17][38] , \sa_snapshot[17].f.upper[6] );
tran (\sa_snapshot[17][37] , \sa_snapshot[17].r.part1[5] );
tran (\sa_snapshot[17][37] , \sa_snapshot[17].f.upper[5] );
tran (\sa_snapshot[17][36] , \sa_snapshot[17].r.part1[4] );
tran (\sa_snapshot[17][36] , \sa_snapshot[17].f.upper[4] );
tran (\sa_snapshot[17][35] , \sa_snapshot[17].r.part1[3] );
tran (\sa_snapshot[17][35] , \sa_snapshot[17].f.upper[3] );
tran (\sa_snapshot[17][34] , \sa_snapshot[17].r.part1[2] );
tran (\sa_snapshot[17][34] , \sa_snapshot[17].f.upper[2] );
tran (\sa_snapshot[17][33] , \sa_snapshot[17].r.part1[1] );
tran (\sa_snapshot[17][33] , \sa_snapshot[17].f.upper[1] );
tran (\sa_snapshot[17][32] , \sa_snapshot[17].r.part1[0] );
tran (\sa_snapshot[17][32] , \sa_snapshot[17].f.upper[0] );
tran (\sa_snapshot[17][31] , \sa_snapshot[17].r.part0[31] );
tran (\sa_snapshot[17][31] , \sa_snapshot[17].f.lower[31] );
tran (\sa_snapshot[17][30] , \sa_snapshot[17].r.part0[30] );
tran (\sa_snapshot[17][30] , \sa_snapshot[17].f.lower[30] );
tran (\sa_snapshot[17][29] , \sa_snapshot[17].r.part0[29] );
tran (\sa_snapshot[17][29] , \sa_snapshot[17].f.lower[29] );
tran (\sa_snapshot[17][28] , \sa_snapshot[17].r.part0[28] );
tran (\sa_snapshot[17][28] , \sa_snapshot[17].f.lower[28] );
tran (\sa_snapshot[17][27] , \sa_snapshot[17].r.part0[27] );
tran (\sa_snapshot[17][27] , \sa_snapshot[17].f.lower[27] );
tran (\sa_snapshot[17][26] , \sa_snapshot[17].r.part0[26] );
tran (\sa_snapshot[17][26] , \sa_snapshot[17].f.lower[26] );
tran (\sa_snapshot[17][25] , \sa_snapshot[17].r.part0[25] );
tran (\sa_snapshot[17][25] , \sa_snapshot[17].f.lower[25] );
tran (\sa_snapshot[17][24] , \sa_snapshot[17].r.part0[24] );
tran (\sa_snapshot[17][24] , \sa_snapshot[17].f.lower[24] );
tran (\sa_snapshot[17][23] , \sa_snapshot[17].r.part0[23] );
tran (\sa_snapshot[17][23] , \sa_snapshot[17].f.lower[23] );
tran (\sa_snapshot[17][22] , \sa_snapshot[17].r.part0[22] );
tran (\sa_snapshot[17][22] , \sa_snapshot[17].f.lower[22] );
tran (\sa_snapshot[17][21] , \sa_snapshot[17].r.part0[21] );
tran (\sa_snapshot[17][21] , \sa_snapshot[17].f.lower[21] );
tran (\sa_snapshot[17][20] , \sa_snapshot[17].r.part0[20] );
tran (\sa_snapshot[17][20] , \sa_snapshot[17].f.lower[20] );
tran (\sa_snapshot[17][19] , \sa_snapshot[17].r.part0[19] );
tran (\sa_snapshot[17][19] , \sa_snapshot[17].f.lower[19] );
tran (\sa_snapshot[17][18] , \sa_snapshot[17].r.part0[18] );
tran (\sa_snapshot[17][18] , \sa_snapshot[17].f.lower[18] );
tran (\sa_snapshot[17][17] , \sa_snapshot[17].r.part0[17] );
tran (\sa_snapshot[17][17] , \sa_snapshot[17].f.lower[17] );
tran (\sa_snapshot[17][16] , \sa_snapshot[17].r.part0[16] );
tran (\sa_snapshot[17][16] , \sa_snapshot[17].f.lower[16] );
tran (\sa_snapshot[17][15] , \sa_snapshot[17].r.part0[15] );
tran (\sa_snapshot[17][15] , \sa_snapshot[17].f.lower[15] );
tran (\sa_snapshot[17][14] , \sa_snapshot[17].r.part0[14] );
tran (\sa_snapshot[17][14] , \sa_snapshot[17].f.lower[14] );
tran (\sa_snapshot[17][13] , \sa_snapshot[17].r.part0[13] );
tran (\sa_snapshot[17][13] , \sa_snapshot[17].f.lower[13] );
tran (\sa_snapshot[17][12] , \sa_snapshot[17].r.part0[12] );
tran (\sa_snapshot[17][12] , \sa_snapshot[17].f.lower[12] );
tran (\sa_snapshot[17][11] , \sa_snapshot[17].r.part0[11] );
tran (\sa_snapshot[17][11] , \sa_snapshot[17].f.lower[11] );
tran (\sa_snapshot[17][10] , \sa_snapshot[17].r.part0[10] );
tran (\sa_snapshot[17][10] , \sa_snapshot[17].f.lower[10] );
tran (\sa_snapshot[17][9] , \sa_snapshot[17].r.part0[9] );
tran (\sa_snapshot[17][9] , \sa_snapshot[17].f.lower[9] );
tran (\sa_snapshot[17][8] , \sa_snapshot[17].r.part0[8] );
tran (\sa_snapshot[17][8] , \sa_snapshot[17].f.lower[8] );
tran (\sa_snapshot[17][7] , \sa_snapshot[17].r.part0[7] );
tran (\sa_snapshot[17][7] , \sa_snapshot[17].f.lower[7] );
tran (\sa_snapshot[17][6] , \sa_snapshot[17].r.part0[6] );
tran (\sa_snapshot[17][6] , \sa_snapshot[17].f.lower[6] );
tran (\sa_snapshot[17][5] , \sa_snapshot[17].r.part0[5] );
tran (\sa_snapshot[17][5] , \sa_snapshot[17].f.lower[5] );
tran (\sa_snapshot[17][4] , \sa_snapshot[17].r.part0[4] );
tran (\sa_snapshot[17][4] , \sa_snapshot[17].f.lower[4] );
tran (\sa_snapshot[17][3] , \sa_snapshot[17].r.part0[3] );
tran (\sa_snapshot[17][3] , \sa_snapshot[17].f.lower[3] );
tran (\sa_snapshot[17][2] , \sa_snapshot[17].r.part0[2] );
tran (\sa_snapshot[17][2] , \sa_snapshot[17].f.lower[2] );
tran (\sa_snapshot[17][1] , \sa_snapshot[17].r.part0[1] );
tran (\sa_snapshot[17][1] , \sa_snapshot[17].f.lower[1] );
tran (\sa_snapshot[17][0] , \sa_snapshot[17].r.part0[0] );
tran (\sa_snapshot[17][0] , \sa_snapshot[17].f.lower[0] );
tran (\sa_snapshot[16][63] , \sa_snapshot[16].r.part1[31] );
tran (\sa_snapshot[16][63] , \sa_snapshot[16].f.unused[13] );
tran (\sa_snapshot[16][62] , \sa_snapshot[16].r.part1[30] );
tran (\sa_snapshot[16][62] , \sa_snapshot[16].f.unused[12] );
tran (\sa_snapshot[16][61] , \sa_snapshot[16].r.part1[29] );
tran (\sa_snapshot[16][61] , \sa_snapshot[16].f.unused[11] );
tran (\sa_snapshot[16][60] , \sa_snapshot[16].r.part1[28] );
tran (\sa_snapshot[16][60] , \sa_snapshot[16].f.unused[10] );
tran (\sa_snapshot[16][59] , \sa_snapshot[16].r.part1[27] );
tran (\sa_snapshot[16][59] , \sa_snapshot[16].f.unused[9] );
tran (\sa_snapshot[16][58] , \sa_snapshot[16].r.part1[26] );
tran (\sa_snapshot[16][58] , \sa_snapshot[16].f.unused[8] );
tran (\sa_snapshot[16][57] , \sa_snapshot[16].r.part1[25] );
tran (\sa_snapshot[16][57] , \sa_snapshot[16].f.unused[7] );
tran (\sa_snapshot[16][56] , \sa_snapshot[16].r.part1[24] );
tran (\sa_snapshot[16][56] , \sa_snapshot[16].f.unused[6] );
tran (\sa_snapshot[16][55] , \sa_snapshot[16].r.part1[23] );
tran (\sa_snapshot[16][55] , \sa_snapshot[16].f.unused[5] );
tran (\sa_snapshot[16][54] , \sa_snapshot[16].r.part1[22] );
tran (\sa_snapshot[16][54] , \sa_snapshot[16].f.unused[4] );
tran (\sa_snapshot[16][53] , \sa_snapshot[16].r.part1[21] );
tran (\sa_snapshot[16][53] , \sa_snapshot[16].f.unused[3] );
tran (\sa_snapshot[16][52] , \sa_snapshot[16].r.part1[20] );
tran (\sa_snapshot[16][52] , \sa_snapshot[16].f.unused[2] );
tran (\sa_snapshot[16][51] , \sa_snapshot[16].r.part1[19] );
tran (\sa_snapshot[16][51] , \sa_snapshot[16].f.unused[1] );
tran (\sa_snapshot[16][50] , \sa_snapshot[16].r.part1[18] );
tran (\sa_snapshot[16][50] , \sa_snapshot[16].f.unused[0] );
tran (\sa_snapshot[16][49] , \sa_snapshot[16].r.part1[17] );
tran (\sa_snapshot[16][49] , \sa_snapshot[16].f.upper[17] );
tran (\sa_snapshot[16][48] , \sa_snapshot[16].r.part1[16] );
tran (\sa_snapshot[16][48] , \sa_snapshot[16].f.upper[16] );
tran (\sa_snapshot[16][47] , \sa_snapshot[16].r.part1[15] );
tran (\sa_snapshot[16][47] , \sa_snapshot[16].f.upper[15] );
tran (\sa_snapshot[16][46] , \sa_snapshot[16].r.part1[14] );
tran (\sa_snapshot[16][46] , \sa_snapshot[16].f.upper[14] );
tran (\sa_snapshot[16][45] , \sa_snapshot[16].r.part1[13] );
tran (\sa_snapshot[16][45] , \sa_snapshot[16].f.upper[13] );
tran (\sa_snapshot[16][44] , \sa_snapshot[16].r.part1[12] );
tran (\sa_snapshot[16][44] , \sa_snapshot[16].f.upper[12] );
tran (\sa_snapshot[16][43] , \sa_snapshot[16].r.part1[11] );
tran (\sa_snapshot[16][43] , \sa_snapshot[16].f.upper[11] );
tran (\sa_snapshot[16][42] , \sa_snapshot[16].r.part1[10] );
tran (\sa_snapshot[16][42] , \sa_snapshot[16].f.upper[10] );
tran (\sa_snapshot[16][41] , \sa_snapshot[16].r.part1[9] );
tran (\sa_snapshot[16][41] , \sa_snapshot[16].f.upper[9] );
tran (\sa_snapshot[16][40] , \sa_snapshot[16].r.part1[8] );
tran (\sa_snapshot[16][40] , \sa_snapshot[16].f.upper[8] );
tran (\sa_snapshot[16][39] , \sa_snapshot[16].r.part1[7] );
tran (\sa_snapshot[16][39] , \sa_snapshot[16].f.upper[7] );
tran (\sa_snapshot[16][38] , \sa_snapshot[16].r.part1[6] );
tran (\sa_snapshot[16][38] , \sa_snapshot[16].f.upper[6] );
tran (\sa_snapshot[16][37] , \sa_snapshot[16].r.part1[5] );
tran (\sa_snapshot[16][37] , \sa_snapshot[16].f.upper[5] );
tran (\sa_snapshot[16][36] , \sa_snapshot[16].r.part1[4] );
tran (\sa_snapshot[16][36] , \sa_snapshot[16].f.upper[4] );
tran (\sa_snapshot[16][35] , \sa_snapshot[16].r.part1[3] );
tran (\sa_snapshot[16][35] , \sa_snapshot[16].f.upper[3] );
tran (\sa_snapshot[16][34] , \sa_snapshot[16].r.part1[2] );
tran (\sa_snapshot[16][34] , \sa_snapshot[16].f.upper[2] );
tran (\sa_snapshot[16][33] , \sa_snapshot[16].r.part1[1] );
tran (\sa_snapshot[16][33] , \sa_snapshot[16].f.upper[1] );
tran (\sa_snapshot[16][32] , \sa_snapshot[16].r.part1[0] );
tran (\sa_snapshot[16][32] , \sa_snapshot[16].f.upper[0] );
tran (\sa_snapshot[16][31] , \sa_snapshot[16].r.part0[31] );
tran (\sa_snapshot[16][31] , \sa_snapshot[16].f.lower[31] );
tran (\sa_snapshot[16][30] , \sa_snapshot[16].r.part0[30] );
tran (\sa_snapshot[16][30] , \sa_snapshot[16].f.lower[30] );
tran (\sa_snapshot[16][29] , \sa_snapshot[16].r.part0[29] );
tran (\sa_snapshot[16][29] , \sa_snapshot[16].f.lower[29] );
tran (\sa_snapshot[16][28] , \sa_snapshot[16].r.part0[28] );
tran (\sa_snapshot[16][28] , \sa_snapshot[16].f.lower[28] );
tran (\sa_snapshot[16][27] , \sa_snapshot[16].r.part0[27] );
tran (\sa_snapshot[16][27] , \sa_snapshot[16].f.lower[27] );
tran (\sa_snapshot[16][26] , \sa_snapshot[16].r.part0[26] );
tran (\sa_snapshot[16][26] , \sa_snapshot[16].f.lower[26] );
tran (\sa_snapshot[16][25] , \sa_snapshot[16].r.part0[25] );
tran (\sa_snapshot[16][25] , \sa_snapshot[16].f.lower[25] );
tran (\sa_snapshot[16][24] , \sa_snapshot[16].r.part0[24] );
tran (\sa_snapshot[16][24] , \sa_snapshot[16].f.lower[24] );
tran (\sa_snapshot[16][23] , \sa_snapshot[16].r.part0[23] );
tran (\sa_snapshot[16][23] , \sa_snapshot[16].f.lower[23] );
tran (\sa_snapshot[16][22] , \sa_snapshot[16].r.part0[22] );
tran (\sa_snapshot[16][22] , \sa_snapshot[16].f.lower[22] );
tran (\sa_snapshot[16][21] , \sa_snapshot[16].r.part0[21] );
tran (\sa_snapshot[16][21] , \sa_snapshot[16].f.lower[21] );
tran (\sa_snapshot[16][20] , \sa_snapshot[16].r.part0[20] );
tran (\sa_snapshot[16][20] , \sa_snapshot[16].f.lower[20] );
tran (\sa_snapshot[16][19] , \sa_snapshot[16].r.part0[19] );
tran (\sa_snapshot[16][19] , \sa_snapshot[16].f.lower[19] );
tran (\sa_snapshot[16][18] , \sa_snapshot[16].r.part0[18] );
tran (\sa_snapshot[16][18] , \sa_snapshot[16].f.lower[18] );
tran (\sa_snapshot[16][17] , \sa_snapshot[16].r.part0[17] );
tran (\sa_snapshot[16][17] , \sa_snapshot[16].f.lower[17] );
tran (\sa_snapshot[16][16] , \sa_snapshot[16].r.part0[16] );
tran (\sa_snapshot[16][16] , \sa_snapshot[16].f.lower[16] );
tran (\sa_snapshot[16][15] , \sa_snapshot[16].r.part0[15] );
tran (\sa_snapshot[16][15] , \sa_snapshot[16].f.lower[15] );
tran (\sa_snapshot[16][14] , \sa_snapshot[16].r.part0[14] );
tran (\sa_snapshot[16][14] , \sa_snapshot[16].f.lower[14] );
tran (\sa_snapshot[16][13] , \sa_snapshot[16].r.part0[13] );
tran (\sa_snapshot[16][13] , \sa_snapshot[16].f.lower[13] );
tran (\sa_snapshot[16][12] , \sa_snapshot[16].r.part0[12] );
tran (\sa_snapshot[16][12] , \sa_snapshot[16].f.lower[12] );
tran (\sa_snapshot[16][11] , \sa_snapshot[16].r.part0[11] );
tran (\sa_snapshot[16][11] , \sa_snapshot[16].f.lower[11] );
tran (\sa_snapshot[16][10] , \sa_snapshot[16].r.part0[10] );
tran (\sa_snapshot[16][10] , \sa_snapshot[16].f.lower[10] );
tran (\sa_snapshot[16][9] , \sa_snapshot[16].r.part0[9] );
tran (\sa_snapshot[16][9] , \sa_snapshot[16].f.lower[9] );
tran (\sa_snapshot[16][8] , \sa_snapshot[16].r.part0[8] );
tran (\sa_snapshot[16][8] , \sa_snapshot[16].f.lower[8] );
tran (\sa_snapshot[16][7] , \sa_snapshot[16].r.part0[7] );
tran (\sa_snapshot[16][7] , \sa_snapshot[16].f.lower[7] );
tran (\sa_snapshot[16][6] , \sa_snapshot[16].r.part0[6] );
tran (\sa_snapshot[16][6] , \sa_snapshot[16].f.lower[6] );
tran (\sa_snapshot[16][5] , \sa_snapshot[16].r.part0[5] );
tran (\sa_snapshot[16][5] , \sa_snapshot[16].f.lower[5] );
tran (\sa_snapshot[16][4] , \sa_snapshot[16].r.part0[4] );
tran (\sa_snapshot[16][4] , \sa_snapshot[16].f.lower[4] );
tran (\sa_snapshot[16][3] , \sa_snapshot[16].r.part0[3] );
tran (\sa_snapshot[16][3] , \sa_snapshot[16].f.lower[3] );
tran (\sa_snapshot[16][2] , \sa_snapshot[16].r.part0[2] );
tran (\sa_snapshot[16][2] , \sa_snapshot[16].f.lower[2] );
tran (\sa_snapshot[16][1] , \sa_snapshot[16].r.part0[1] );
tran (\sa_snapshot[16][1] , \sa_snapshot[16].f.lower[1] );
tran (\sa_snapshot[16][0] , \sa_snapshot[16].r.part0[0] );
tran (\sa_snapshot[16][0] , \sa_snapshot[16].f.lower[0] );
tran (\sa_snapshot[15][63] , \sa_snapshot[15].r.part1[31] );
tran (\sa_snapshot[15][63] , \sa_snapshot[15].f.unused[13] );
tran (\sa_snapshot[15][62] , \sa_snapshot[15].r.part1[30] );
tran (\sa_snapshot[15][62] , \sa_snapshot[15].f.unused[12] );
tran (\sa_snapshot[15][61] , \sa_snapshot[15].r.part1[29] );
tran (\sa_snapshot[15][61] , \sa_snapshot[15].f.unused[11] );
tran (\sa_snapshot[15][60] , \sa_snapshot[15].r.part1[28] );
tran (\sa_snapshot[15][60] , \sa_snapshot[15].f.unused[10] );
tran (\sa_snapshot[15][59] , \sa_snapshot[15].r.part1[27] );
tran (\sa_snapshot[15][59] , \sa_snapshot[15].f.unused[9] );
tran (\sa_snapshot[15][58] , \sa_snapshot[15].r.part1[26] );
tran (\sa_snapshot[15][58] , \sa_snapshot[15].f.unused[8] );
tran (\sa_snapshot[15][57] , \sa_snapshot[15].r.part1[25] );
tran (\sa_snapshot[15][57] , \sa_snapshot[15].f.unused[7] );
tran (\sa_snapshot[15][56] , \sa_snapshot[15].r.part1[24] );
tran (\sa_snapshot[15][56] , \sa_snapshot[15].f.unused[6] );
tran (\sa_snapshot[15][55] , \sa_snapshot[15].r.part1[23] );
tran (\sa_snapshot[15][55] , \sa_snapshot[15].f.unused[5] );
tran (\sa_snapshot[15][54] , \sa_snapshot[15].r.part1[22] );
tran (\sa_snapshot[15][54] , \sa_snapshot[15].f.unused[4] );
tran (\sa_snapshot[15][53] , \sa_snapshot[15].r.part1[21] );
tran (\sa_snapshot[15][53] , \sa_snapshot[15].f.unused[3] );
tran (\sa_snapshot[15][52] , \sa_snapshot[15].r.part1[20] );
tran (\sa_snapshot[15][52] , \sa_snapshot[15].f.unused[2] );
tran (\sa_snapshot[15][51] , \sa_snapshot[15].r.part1[19] );
tran (\sa_snapshot[15][51] , \sa_snapshot[15].f.unused[1] );
tran (\sa_snapshot[15][50] , \sa_snapshot[15].r.part1[18] );
tran (\sa_snapshot[15][50] , \sa_snapshot[15].f.unused[0] );
tran (\sa_snapshot[15][49] , \sa_snapshot[15].r.part1[17] );
tran (\sa_snapshot[15][49] , \sa_snapshot[15].f.upper[17] );
tran (\sa_snapshot[15][48] , \sa_snapshot[15].r.part1[16] );
tran (\sa_snapshot[15][48] , \sa_snapshot[15].f.upper[16] );
tran (\sa_snapshot[15][47] , \sa_snapshot[15].r.part1[15] );
tran (\sa_snapshot[15][47] , \sa_snapshot[15].f.upper[15] );
tran (\sa_snapshot[15][46] , \sa_snapshot[15].r.part1[14] );
tran (\sa_snapshot[15][46] , \sa_snapshot[15].f.upper[14] );
tran (\sa_snapshot[15][45] , \sa_snapshot[15].r.part1[13] );
tran (\sa_snapshot[15][45] , \sa_snapshot[15].f.upper[13] );
tran (\sa_snapshot[15][44] , \sa_snapshot[15].r.part1[12] );
tran (\sa_snapshot[15][44] , \sa_snapshot[15].f.upper[12] );
tran (\sa_snapshot[15][43] , \sa_snapshot[15].r.part1[11] );
tran (\sa_snapshot[15][43] , \sa_snapshot[15].f.upper[11] );
tran (\sa_snapshot[15][42] , \sa_snapshot[15].r.part1[10] );
tran (\sa_snapshot[15][42] , \sa_snapshot[15].f.upper[10] );
tran (\sa_snapshot[15][41] , \sa_snapshot[15].r.part1[9] );
tran (\sa_snapshot[15][41] , \sa_snapshot[15].f.upper[9] );
tran (\sa_snapshot[15][40] , \sa_snapshot[15].r.part1[8] );
tran (\sa_snapshot[15][40] , \sa_snapshot[15].f.upper[8] );
tran (\sa_snapshot[15][39] , \sa_snapshot[15].r.part1[7] );
tran (\sa_snapshot[15][39] , \sa_snapshot[15].f.upper[7] );
tran (\sa_snapshot[15][38] , \sa_snapshot[15].r.part1[6] );
tran (\sa_snapshot[15][38] , \sa_snapshot[15].f.upper[6] );
tran (\sa_snapshot[15][37] , \sa_snapshot[15].r.part1[5] );
tran (\sa_snapshot[15][37] , \sa_snapshot[15].f.upper[5] );
tran (\sa_snapshot[15][36] , \sa_snapshot[15].r.part1[4] );
tran (\sa_snapshot[15][36] , \sa_snapshot[15].f.upper[4] );
tran (\sa_snapshot[15][35] , \sa_snapshot[15].r.part1[3] );
tran (\sa_snapshot[15][35] , \sa_snapshot[15].f.upper[3] );
tran (\sa_snapshot[15][34] , \sa_snapshot[15].r.part1[2] );
tran (\sa_snapshot[15][34] , \sa_snapshot[15].f.upper[2] );
tran (\sa_snapshot[15][33] , \sa_snapshot[15].r.part1[1] );
tran (\sa_snapshot[15][33] , \sa_snapshot[15].f.upper[1] );
tran (\sa_snapshot[15][32] , \sa_snapshot[15].r.part1[0] );
tran (\sa_snapshot[15][32] , \sa_snapshot[15].f.upper[0] );
tran (\sa_snapshot[15][31] , \sa_snapshot[15].r.part0[31] );
tran (\sa_snapshot[15][31] , \sa_snapshot[15].f.lower[31] );
tran (\sa_snapshot[15][30] , \sa_snapshot[15].r.part0[30] );
tran (\sa_snapshot[15][30] , \sa_snapshot[15].f.lower[30] );
tran (\sa_snapshot[15][29] , \sa_snapshot[15].r.part0[29] );
tran (\sa_snapshot[15][29] , \sa_snapshot[15].f.lower[29] );
tran (\sa_snapshot[15][28] , \sa_snapshot[15].r.part0[28] );
tran (\sa_snapshot[15][28] , \sa_snapshot[15].f.lower[28] );
tran (\sa_snapshot[15][27] , \sa_snapshot[15].r.part0[27] );
tran (\sa_snapshot[15][27] , \sa_snapshot[15].f.lower[27] );
tran (\sa_snapshot[15][26] , \sa_snapshot[15].r.part0[26] );
tran (\sa_snapshot[15][26] , \sa_snapshot[15].f.lower[26] );
tran (\sa_snapshot[15][25] , \sa_snapshot[15].r.part0[25] );
tran (\sa_snapshot[15][25] , \sa_snapshot[15].f.lower[25] );
tran (\sa_snapshot[15][24] , \sa_snapshot[15].r.part0[24] );
tran (\sa_snapshot[15][24] , \sa_snapshot[15].f.lower[24] );
tran (\sa_snapshot[15][23] , \sa_snapshot[15].r.part0[23] );
tran (\sa_snapshot[15][23] , \sa_snapshot[15].f.lower[23] );
tran (\sa_snapshot[15][22] , \sa_snapshot[15].r.part0[22] );
tran (\sa_snapshot[15][22] , \sa_snapshot[15].f.lower[22] );
tran (\sa_snapshot[15][21] , \sa_snapshot[15].r.part0[21] );
tran (\sa_snapshot[15][21] , \sa_snapshot[15].f.lower[21] );
tran (\sa_snapshot[15][20] , \sa_snapshot[15].r.part0[20] );
tran (\sa_snapshot[15][20] , \sa_snapshot[15].f.lower[20] );
tran (\sa_snapshot[15][19] , \sa_snapshot[15].r.part0[19] );
tran (\sa_snapshot[15][19] , \sa_snapshot[15].f.lower[19] );
tran (\sa_snapshot[15][18] , \sa_snapshot[15].r.part0[18] );
tran (\sa_snapshot[15][18] , \sa_snapshot[15].f.lower[18] );
tran (\sa_snapshot[15][17] , \sa_snapshot[15].r.part0[17] );
tran (\sa_snapshot[15][17] , \sa_snapshot[15].f.lower[17] );
tran (\sa_snapshot[15][16] , \sa_snapshot[15].r.part0[16] );
tran (\sa_snapshot[15][16] , \sa_snapshot[15].f.lower[16] );
tran (\sa_snapshot[15][15] , \sa_snapshot[15].r.part0[15] );
tran (\sa_snapshot[15][15] , \sa_snapshot[15].f.lower[15] );
tran (\sa_snapshot[15][14] , \sa_snapshot[15].r.part0[14] );
tran (\sa_snapshot[15][14] , \sa_snapshot[15].f.lower[14] );
tran (\sa_snapshot[15][13] , \sa_snapshot[15].r.part0[13] );
tran (\sa_snapshot[15][13] , \sa_snapshot[15].f.lower[13] );
tran (\sa_snapshot[15][12] , \sa_snapshot[15].r.part0[12] );
tran (\sa_snapshot[15][12] , \sa_snapshot[15].f.lower[12] );
tran (\sa_snapshot[15][11] , \sa_snapshot[15].r.part0[11] );
tran (\sa_snapshot[15][11] , \sa_snapshot[15].f.lower[11] );
tran (\sa_snapshot[15][10] , \sa_snapshot[15].r.part0[10] );
tran (\sa_snapshot[15][10] , \sa_snapshot[15].f.lower[10] );
tran (\sa_snapshot[15][9] , \sa_snapshot[15].r.part0[9] );
tran (\sa_snapshot[15][9] , \sa_snapshot[15].f.lower[9] );
tran (\sa_snapshot[15][8] , \sa_snapshot[15].r.part0[8] );
tran (\sa_snapshot[15][8] , \sa_snapshot[15].f.lower[8] );
tran (\sa_snapshot[15][7] , \sa_snapshot[15].r.part0[7] );
tran (\sa_snapshot[15][7] , \sa_snapshot[15].f.lower[7] );
tran (\sa_snapshot[15][6] , \sa_snapshot[15].r.part0[6] );
tran (\sa_snapshot[15][6] , \sa_snapshot[15].f.lower[6] );
tran (\sa_snapshot[15][5] , \sa_snapshot[15].r.part0[5] );
tran (\sa_snapshot[15][5] , \sa_snapshot[15].f.lower[5] );
tran (\sa_snapshot[15][4] , \sa_snapshot[15].r.part0[4] );
tran (\sa_snapshot[15][4] , \sa_snapshot[15].f.lower[4] );
tran (\sa_snapshot[15][3] , \sa_snapshot[15].r.part0[3] );
tran (\sa_snapshot[15][3] , \sa_snapshot[15].f.lower[3] );
tran (\sa_snapshot[15][2] , \sa_snapshot[15].r.part0[2] );
tran (\sa_snapshot[15][2] , \sa_snapshot[15].f.lower[2] );
tran (\sa_snapshot[15][1] , \sa_snapshot[15].r.part0[1] );
tran (\sa_snapshot[15][1] , \sa_snapshot[15].f.lower[1] );
tran (\sa_snapshot[15][0] , \sa_snapshot[15].r.part0[0] );
tran (\sa_snapshot[15][0] , \sa_snapshot[15].f.lower[0] );
tran (\sa_snapshot[14][63] , \sa_snapshot[14].r.part1[31] );
tran (\sa_snapshot[14][63] , \sa_snapshot[14].f.unused[13] );
tran (\sa_snapshot[14][62] , \sa_snapshot[14].r.part1[30] );
tran (\sa_snapshot[14][62] , \sa_snapshot[14].f.unused[12] );
tran (\sa_snapshot[14][61] , \sa_snapshot[14].r.part1[29] );
tran (\sa_snapshot[14][61] , \sa_snapshot[14].f.unused[11] );
tran (\sa_snapshot[14][60] , \sa_snapshot[14].r.part1[28] );
tran (\sa_snapshot[14][60] , \sa_snapshot[14].f.unused[10] );
tran (\sa_snapshot[14][59] , \sa_snapshot[14].r.part1[27] );
tran (\sa_snapshot[14][59] , \sa_snapshot[14].f.unused[9] );
tran (\sa_snapshot[14][58] , \sa_snapshot[14].r.part1[26] );
tran (\sa_snapshot[14][58] , \sa_snapshot[14].f.unused[8] );
tran (\sa_snapshot[14][57] , \sa_snapshot[14].r.part1[25] );
tran (\sa_snapshot[14][57] , \sa_snapshot[14].f.unused[7] );
tran (\sa_snapshot[14][56] , \sa_snapshot[14].r.part1[24] );
tran (\sa_snapshot[14][56] , \sa_snapshot[14].f.unused[6] );
tran (\sa_snapshot[14][55] , \sa_snapshot[14].r.part1[23] );
tran (\sa_snapshot[14][55] , \sa_snapshot[14].f.unused[5] );
tran (\sa_snapshot[14][54] , \sa_snapshot[14].r.part1[22] );
tran (\sa_snapshot[14][54] , \sa_snapshot[14].f.unused[4] );
tran (\sa_snapshot[14][53] , \sa_snapshot[14].r.part1[21] );
tran (\sa_snapshot[14][53] , \sa_snapshot[14].f.unused[3] );
tran (\sa_snapshot[14][52] , \sa_snapshot[14].r.part1[20] );
tran (\sa_snapshot[14][52] , \sa_snapshot[14].f.unused[2] );
tran (\sa_snapshot[14][51] , \sa_snapshot[14].r.part1[19] );
tran (\sa_snapshot[14][51] , \sa_snapshot[14].f.unused[1] );
tran (\sa_snapshot[14][50] , \sa_snapshot[14].r.part1[18] );
tran (\sa_snapshot[14][50] , \sa_snapshot[14].f.unused[0] );
tran (\sa_snapshot[14][49] , \sa_snapshot[14].r.part1[17] );
tran (\sa_snapshot[14][49] , \sa_snapshot[14].f.upper[17] );
tran (\sa_snapshot[14][48] , \sa_snapshot[14].r.part1[16] );
tran (\sa_snapshot[14][48] , \sa_snapshot[14].f.upper[16] );
tran (\sa_snapshot[14][47] , \sa_snapshot[14].r.part1[15] );
tran (\sa_snapshot[14][47] , \sa_snapshot[14].f.upper[15] );
tran (\sa_snapshot[14][46] , \sa_snapshot[14].r.part1[14] );
tran (\sa_snapshot[14][46] , \sa_snapshot[14].f.upper[14] );
tran (\sa_snapshot[14][45] , \sa_snapshot[14].r.part1[13] );
tran (\sa_snapshot[14][45] , \sa_snapshot[14].f.upper[13] );
tran (\sa_snapshot[14][44] , \sa_snapshot[14].r.part1[12] );
tran (\sa_snapshot[14][44] , \sa_snapshot[14].f.upper[12] );
tran (\sa_snapshot[14][43] , \sa_snapshot[14].r.part1[11] );
tran (\sa_snapshot[14][43] , \sa_snapshot[14].f.upper[11] );
tran (\sa_snapshot[14][42] , \sa_snapshot[14].r.part1[10] );
tran (\sa_snapshot[14][42] , \sa_snapshot[14].f.upper[10] );
tran (\sa_snapshot[14][41] , \sa_snapshot[14].r.part1[9] );
tran (\sa_snapshot[14][41] , \sa_snapshot[14].f.upper[9] );
tran (\sa_snapshot[14][40] , \sa_snapshot[14].r.part1[8] );
tran (\sa_snapshot[14][40] , \sa_snapshot[14].f.upper[8] );
tran (\sa_snapshot[14][39] , \sa_snapshot[14].r.part1[7] );
tran (\sa_snapshot[14][39] , \sa_snapshot[14].f.upper[7] );
tran (\sa_snapshot[14][38] , \sa_snapshot[14].r.part1[6] );
tran (\sa_snapshot[14][38] , \sa_snapshot[14].f.upper[6] );
tran (\sa_snapshot[14][37] , \sa_snapshot[14].r.part1[5] );
tran (\sa_snapshot[14][37] , \sa_snapshot[14].f.upper[5] );
tran (\sa_snapshot[14][36] , \sa_snapshot[14].r.part1[4] );
tran (\sa_snapshot[14][36] , \sa_snapshot[14].f.upper[4] );
tran (\sa_snapshot[14][35] , \sa_snapshot[14].r.part1[3] );
tran (\sa_snapshot[14][35] , \sa_snapshot[14].f.upper[3] );
tran (\sa_snapshot[14][34] , \sa_snapshot[14].r.part1[2] );
tran (\sa_snapshot[14][34] , \sa_snapshot[14].f.upper[2] );
tran (\sa_snapshot[14][33] , \sa_snapshot[14].r.part1[1] );
tran (\sa_snapshot[14][33] , \sa_snapshot[14].f.upper[1] );
tran (\sa_snapshot[14][32] , \sa_snapshot[14].r.part1[0] );
tran (\sa_snapshot[14][32] , \sa_snapshot[14].f.upper[0] );
tran (\sa_snapshot[14][31] , \sa_snapshot[14].r.part0[31] );
tran (\sa_snapshot[14][31] , \sa_snapshot[14].f.lower[31] );
tran (\sa_snapshot[14][30] , \sa_snapshot[14].r.part0[30] );
tran (\sa_snapshot[14][30] , \sa_snapshot[14].f.lower[30] );
tran (\sa_snapshot[14][29] , \sa_snapshot[14].r.part0[29] );
tran (\sa_snapshot[14][29] , \sa_snapshot[14].f.lower[29] );
tran (\sa_snapshot[14][28] , \sa_snapshot[14].r.part0[28] );
tran (\sa_snapshot[14][28] , \sa_snapshot[14].f.lower[28] );
tran (\sa_snapshot[14][27] , \sa_snapshot[14].r.part0[27] );
tran (\sa_snapshot[14][27] , \sa_snapshot[14].f.lower[27] );
tran (\sa_snapshot[14][26] , \sa_snapshot[14].r.part0[26] );
tran (\sa_snapshot[14][26] , \sa_snapshot[14].f.lower[26] );
tran (\sa_snapshot[14][25] , \sa_snapshot[14].r.part0[25] );
tran (\sa_snapshot[14][25] , \sa_snapshot[14].f.lower[25] );
tran (\sa_snapshot[14][24] , \sa_snapshot[14].r.part0[24] );
tran (\sa_snapshot[14][24] , \sa_snapshot[14].f.lower[24] );
tran (\sa_snapshot[14][23] , \sa_snapshot[14].r.part0[23] );
tran (\sa_snapshot[14][23] , \sa_snapshot[14].f.lower[23] );
tran (\sa_snapshot[14][22] , \sa_snapshot[14].r.part0[22] );
tran (\sa_snapshot[14][22] , \sa_snapshot[14].f.lower[22] );
tran (\sa_snapshot[14][21] , \sa_snapshot[14].r.part0[21] );
tran (\sa_snapshot[14][21] , \sa_snapshot[14].f.lower[21] );
tran (\sa_snapshot[14][20] , \sa_snapshot[14].r.part0[20] );
tran (\sa_snapshot[14][20] , \sa_snapshot[14].f.lower[20] );
tran (\sa_snapshot[14][19] , \sa_snapshot[14].r.part0[19] );
tran (\sa_snapshot[14][19] , \sa_snapshot[14].f.lower[19] );
tran (\sa_snapshot[14][18] , \sa_snapshot[14].r.part0[18] );
tran (\sa_snapshot[14][18] , \sa_snapshot[14].f.lower[18] );
tran (\sa_snapshot[14][17] , \sa_snapshot[14].r.part0[17] );
tran (\sa_snapshot[14][17] , \sa_snapshot[14].f.lower[17] );
tran (\sa_snapshot[14][16] , \sa_snapshot[14].r.part0[16] );
tran (\sa_snapshot[14][16] , \sa_snapshot[14].f.lower[16] );
tran (\sa_snapshot[14][15] , \sa_snapshot[14].r.part0[15] );
tran (\sa_snapshot[14][15] , \sa_snapshot[14].f.lower[15] );
tran (\sa_snapshot[14][14] , \sa_snapshot[14].r.part0[14] );
tran (\sa_snapshot[14][14] , \sa_snapshot[14].f.lower[14] );
tran (\sa_snapshot[14][13] , \sa_snapshot[14].r.part0[13] );
tran (\sa_snapshot[14][13] , \sa_snapshot[14].f.lower[13] );
tran (\sa_snapshot[14][12] , \sa_snapshot[14].r.part0[12] );
tran (\sa_snapshot[14][12] , \sa_snapshot[14].f.lower[12] );
tran (\sa_snapshot[14][11] , \sa_snapshot[14].r.part0[11] );
tran (\sa_snapshot[14][11] , \sa_snapshot[14].f.lower[11] );
tran (\sa_snapshot[14][10] , \sa_snapshot[14].r.part0[10] );
tran (\sa_snapshot[14][10] , \sa_snapshot[14].f.lower[10] );
tran (\sa_snapshot[14][9] , \sa_snapshot[14].r.part0[9] );
tran (\sa_snapshot[14][9] , \sa_snapshot[14].f.lower[9] );
tran (\sa_snapshot[14][8] , \sa_snapshot[14].r.part0[8] );
tran (\sa_snapshot[14][8] , \sa_snapshot[14].f.lower[8] );
tran (\sa_snapshot[14][7] , \sa_snapshot[14].r.part0[7] );
tran (\sa_snapshot[14][7] , \sa_snapshot[14].f.lower[7] );
tran (\sa_snapshot[14][6] , \sa_snapshot[14].r.part0[6] );
tran (\sa_snapshot[14][6] , \sa_snapshot[14].f.lower[6] );
tran (\sa_snapshot[14][5] , \sa_snapshot[14].r.part0[5] );
tran (\sa_snapshot[14][5] , \sa_snapshot[14].f.lower[5] );
tran (\sa_snapshot[14][4] , \sa_snapshot[14].r.part0[4] );
tran (\sa_snapshot[14][4] , \sa_snapshot[14].f.lower[4] );
tran (\sa_snapshot[14][3] , \sa_snapshot[14].r.part0[3] );
tran (\sa_snapshot[14][3] , \sa_snapshot[14].f.lower[3] );
tran (\sa_snapshot[14][2] , \sa_snapshot[14].r.part0[2] );
tran (\sa_snapshot[14][2] , \sa_snapshot[14].f.lower[2] );
tran (\sa_snapshot[14][1] , \sa_snapshot[14].r.part0[1] );
tran (\sa_snapshot[14][1] , \sa_snapshot[14].f.lower[1] );
tran (\sa_snapshot[14][0] , \sa_snapshot[14].r.part0[0] );
tran (\sa_snapshot[14][0] , \sa_snapshot[14].f.lower[0] );
tran (\sa_snapshot[13][63] , \sa_snapshot[13].r.part1[31] );
tran (\sa_snapshot[13][63] , \sa_snapshot[13].f.unused[13] );
tran (\sa_snapshot[13][62] , \sa_snapshot[13].r.part1[30] );
tran (\sa_snapshot[13][62] , \sa_snapshot[13].f.unused[12] );
tran (\sa_snapshot[13][61] , \sa_snapshot[13].r.part1[29] );
tran (\sa_snapshot[13][61] , \sa_snapshot[13].f.unused[11] );
tran (\sa_snapshot[13][60] , \sa_snapshot[13].r.part1[28] );
tran (\sa_snapshot[13][60] , \sa_snapshot[13].f.unused[10] );
tran (\sa_snapshot[13][59] , \sa_snapshot[13].r.part1[27] );
tran (\sa_snapshot[13][59] , \sa_snapshot[13].f.unused[9] );
tran (\sa_snapshot[13][58] , \sa_snapshot[13].r.part1[26] );
tran (\sa_snapshot[13][58] , \sa_snapshot[13].f.unused[8] );
tran (\sa_snapshot[13][57] , \sa_snapshot[13].r.part1[25] );
tran (\sa_snapshot[13][57] , \sa_snapshot[13].f.unused[7] );
tran (\sa_snapshot[13][56] , \sa_snapshot[13].r.part1[24] );
tran (\sa_snapshot[13][56] , \sa_snapshot[13].f.unused[6] );
tran (\sa_snapshot[13][55] , \sa_snapshot[13].r.part1[23] );
tran (\sa_snapshot[13][55] , \sa_snapshot[13].f.unused[5] );
tran (\sa_snapshot[13][54] , \sa_snapshot[13].r.part1[22] );
tran (\sa_snapshot[13][54] , \sa_snapshot[13].f.unused[4] );
tran (\sa_snapshot[13][53] , \sa_snapshot[13].r.part1[21] );
tran (\sa_snapshot[13][53] , \sa_snapshot[13].f.unused[3] );
tran (\sa_snapshot[13][52] , \sa_snapshot[13].r.part1[20] );
tran (\sa_snapshot[13][52] , \sa_snapshot[13].f.unused[2] );
tran (\sa_snapshot[13][51] , \sa_snapshot[13].r.part1[19] );
tran (\sa_snapshot[13][51] , \sa_snapshot[13].f.unused[1] );
tran (\sa_snapshot[13][50] , \sa_snapshot[13].r.part1[18] );
tran (\sa_snapshot[13][50] , \sa_snapshot[13].f.unused[0] );
tran (\sa_snapshot[13][49] , \sa_snapshot[13].r.part1[17] );
tran (\sa_snapshot[13][49] , \sa_snapshot[13].f.upper[17] );
tran (\sa_snapshot[13][48] , \sa_snapshot[13].r.part1[16] );
tran (\sa_snapshot[13][48] , \sa_snapshot[13].f.upper[16] );
tran (\sa_snapshot[13][47] , \sa_snapshot[13].r.part1[15] );
tran (\sa_snapshot[13][47] , \sa_snapshot[13].f.upper[15] );
tran (\sa_snapshot[13][46] , \sa_snapshot[13].r.part1[14] );
tran (\sa_snapshot[13][46] , \sa_snapshot[13].f.upper[14] );
tran (\sa_snapshot[13][45] , \sa_snapshot[13].r.part1[13] );
tran (\sa_snapshot[13][45] , \sa_snapshot[13].f.upper[13] );
tran (\sa_snapshot[13][44] , \sa_snapshot[13].r.part1[12] );
tran (\sa_snapshot[13][44] , \sa_snapshot[13].f.upper[12] );
tran (\sa_snapshot[13][43] , \sa_snapshot[13].r.part1[11] );
tran (\sa_snapshot[13][43] , \sa_snapshot[13].f.upper[11] );
tran (\sa_snapshot[13][42] , \sa_snapshot[13].r.part1[10] );
tran (\sa_snapshot[13][42] , \sa_snapshot[13].f.upper[10] );
tran (\sa_snapshot[13][41] , \sa_snapshot[13].r.part1[9] );
tran (\sa_snapshot[13][41] , \sa_snapshot[13].f.upper[9] );
tran (\sa_snapshot[13][40] , \sa_snapshot[13].r.part1[8] );
tran (\sa_snapshot[13][40] , \sa_snapshot[13].f.upper[8] );
tran (\sa_snapshot[13][39] , \sa_snapshot[13].r.part1[7] );
tran (\sa_snapshot[13][39] , \sa_snapshot[13].f.upper[7] );
tran (\sa_snapshot[13][38] , \sa_snapshot[13].r.part1[6] );
tran (\sa_snapshot[13][38] , \sa_snapshot[13].f.upper[6] );
tran (\sa_snapshot[13][37] , \sa_snapshot[13].r.part1[5] );
tran (\sa_snapshot[13][37] , \sa_snapshot[13].f.upper[5] );
tran (\sa_snapshot[13][36] , \sa_snapshot[13].r.part1[4] );
tran (\sa_snapshot[13][36] , \sa_snapshot[13].f.upper[4] );
tran (\sa_snapshot[13][35] , \sa_snapshot[13].r.part1[3] );
tran (\sa_snapshot[13][35] , \sa_snapshot[13].f.upper[3] );
tran (\sa_snapshot[13][34] , \sa_snapshot[13].r.part1[2] );
tran (\sa_snapshot[13][34] , \sa_snapshot[13].f.upper[2] );
tran (\sa_snapshot[13][33] , \sa_snapshot[13].r.part1[1] );
tran (\sa_snapshot[13][33] , \sa_snapshot[13].f.upper[1] );
tran (\sa_snapshot[13][32] , \sa_snapshot[13].r.part1[0] );
tran (\sa_snapshot[13][32] , \sa_snapshot[13].f.upper[0] );
tran (\sa_snapshot[13][31] , \sa_snapshot[13].r.part0[31] );
tran (\sa_snapshot[13][31] , \sa_snapshot[13].f.lower[31] );
tran (\sa_snapshot[13][30] , \sa_snapshot[13].r.part0[30] );
tran (\sa_snapshot[13][30] , \sa_snapshot[13].f.lower[30] );
tran (\sa_snapshot[13][29] , \sa_snapshot[13].r.part0[29] );
tran (\sa_snapshot[13][29] , \sa_snapshot[13].f.lower[29] );
tran (\sa_snapshot[13][28] , \sa_snapshot[13].r.part0[28] );
tran (\sa_snapshot[13][28] , \sa_snapshot[13].f.lower[28] );
tran (\sa_snapshot[13][27] , \sa_snapshot[13].r.part0[27] );
tran (\sa_snapshot[13][27] , \sa_snapshot[13].f.lower[27] );
tran (\sa_snapshot[13][26] , \sa_snapshot[13].r.part0[26] );
tran (\sa_snapshot[13][26] , \sa_snapshot[13].f.lower[26] );
tran (\sa_snapshot[13][25] , \sa_snapshot[13].r.part0[25] );
tran (\sa_snapshot[13][25] , \sa_snapshot[13].f.lower[25] );
tran (\sa_snapshot[13][24] , \sa_snapshot[13].r.part0[24] );
tran (\sa_snapshot[13][24] , \sa_snapshot[13].f.lower[24] );
tran (\sa_snapshot[13][23] , \sa_snapshot[13].r.part0[23] );
tran (\sa_snapshot[13][23] , \sa_snapshot[13].f.lower[23] );
tran (\sa_snapshot[13][22] , \sa_snapshot[13].r.part0[22] );
tran (\sa_snapshot[13][22] , \sa_snapshot[13].f.lower[22] );
tran (\sa_snapshot[13][21] , \sa_snapshot[13].r.part0[21] );
tran (\sa_snapshot[13][21] , \sa_snapshot[13].f.lower[21] );
tran (\sa_snapshot[13][20] , \sa_snapshot[13].r.part0[20] );
tran (\sa_snapshot[13][20] , \sa_snapshot[13].f.lower[20] );
tran (\sa_snapshot[13][19] , \sa_snapshot[13].r.part0[19] );
tran (\sa_snapshot[13][19] , \sa_snapshot[13].f.lower[19] );
tran (\sa_snapshot[13][18] , \sa_snapshot[13].r.part0[18] );
tran (\sa_snapshot[13][18] , \sa_snapshot[13].f.lower[18] );
tran (\sa_snapshot[13][17] , \sa_snapshot[13].r.part0[17] );
tran (\sa_snapshot[13][17] , \sa_snapshot[13].f.lower[17] );
tran (\sa_snapshot[13][16] , \sa_snapshot[13].r.part0[16] );
tran (\sa_snapshot[13][16] , \sa_snapshot[13].f.lower[16] );
tran (\sa_snapshot[13][15] , \sa_snapshot[13].r.part0[15] );
tran (\sa_snapshot[13][15] , \sa_snapshot[13].f.lower[15] );
tran (\sa_snapshot[13][14] , \sa_snapshot[13].r.part0[14] );
tran (\sa_snapshot[13][14] , \sa_snapshot[13].f.lower[14] );
tran (\sa_snapshot[13][13] , \sa_snapshot[13].r.part0[13] );
tran (\sa_snapshot[13][13] , \sa_snapshot[13].f.lower[13] );
tran (\sa_snapshot[13][12] , \sa_snapshot[13].r.part0[12] );
tran (\sa_snapshot[13][12] , \sa_snapshot[13].f.lower[12] );
tran (\sa_snapshot[13][11] , \sa_snapshot[13].r.part0[11] );
tran (\sa_snapshot[13][11] , \sa_snapshot[13].f.lower[11] );
tran (\sa_snapshot[13][10] , \sa_snapshot[13].r.part0[10] );
tran (\sa_snapshot[13][10] , \sa_snapshot[13].f.lower[10] );
tran (\sa_snapshot[13][9] , \sa_snapshot[13].r.part0[9] );
tran (\sa_snapshot[13][9] , \sa_snapshot[13].f.lower[9] );
tran (\sa_snapshot[13][8] , \sa_snapshot[13].r.part0[8] );
tran (\sa_snapshot[13][8] , \sa_snapshot[13].f.lower[8] );
tran (\sa_snapshot[13][7] , \sa_snapshot[13].r.part0[7] );
tran (\sa_snapshot[13][7] , \sa_snapshot[13].f.lower[7] );
tran (\sa_snapshot[13][6] , \sa_snapshot[13].r.part0[6] );
tran (\sa_snapshot[13][6] , \sa_snapshot[13].f.lower[6] );
tran (\sa_snapshot[13][5] , \sa_snapshot[13].r.part0[5] );
tran (\sa_snapshot[13][5] , \sa_snapshot[13].f.lower[5] );
tran (\sa_snapshot[13][4] , \sa_snapshot[13].r.part0[4] );
tran (\sa_snapshot[13][4] , \sa_snapshot[13].f.lower[4] );
tran (\sa_snapshot[13][3] , \sa_snapshot[13].r.part0[3] );
tran (\sa_snapshot[13][3] , \sa_snapshot[13].f.lower[3] );
tran (\sa_snapshot[13][2] , \sa_snapshot[13].r.part0[2] );
tran (\sa_snapshot[13][2] , \sa_snapshot[13].f.lower[2] );
tran (\sa_snapshot[13][1] , \sa_snapshot[13].r.part0[1] );
tran (\sa_snapshot[13][1] , \sa_snapshot[13].f.lower[1] );
tran (\sa_snapshot[13][0] , \sa_snapshot[13].r.part0[0] );
tran (\sa_snapshot[13][0] , \sa_snapshot[13].f.lower[0] );
tran (\sa_snapshot[12][63] , \sa_snapshot[12].r.part1[31] );
tran (\sa_snapshot[12][63] , \sa_snapshot[12].f.unused[13] );
tran (\sa_snapshot[12][62] , \sa_snapshot[12].r.part1[30] );
tran (\sa_snapshot[12][62] , \sa_snapshot[12].f.unused[12] );
tran (\sa_snapshot[12][61] , \sa_snapshot[12].r.part1[29] );
tran (\sa_snapshot[12][61] , \sa_snapshot[12].f.unused[11] );
tran (\sa_snapshot[12][60] , \sa_snapshot[12].r.part1[28] );
tran (\sa_snapshot[12][60] , \sa_snapshot[12].f.unused[10] );
tran (\sa_snapshot[12][59] , \sa_snapshot[12].r.part1[27] );
tran (\sa_snapshot[12][59] , \sa_snapshot[12].f.unused[9] );
tran (\sa_snapshot[12][58] , \sa_snapshot[12].r.part1[26] );
tran (\sa_snapshot[12][58] , \sa_snapshot[12].f.unused[8] );
tran (\sa_snapshot[12][57] , \sa_snapshot[12].r.part1[25] );
tran (\sa_snapshot[12][57] , \sa_snapshot[12].f.unused[7] );
tran (\sa_snapshot[12][56] , \sa_snapshot[12].r.part1[24] );
tran (\sa_snapshot[12][56] , \sa_snapshot[12].f.unused[6] );
tran (\sa_snapshot[12][55] , \sa_snapshot[12].r.part1[23] );
tran (\sa_snapshot[12][55] , \sa_snapshot[12].f.unused[5] );
tran (\sa_snapshot[12][54] , \sa_snapshot[12].r.part1[22] );
tran (\sa_snapshot[12][54] , \sa_snapshot[12].f.unused[4] );
tran (\sa_snapshot[12][53] , \sa_snapshot[12].r.part1[21] );
tran (\sa_snapshot[12][53] , \sa_snapshot[12].f.unused[3] );
tran (\sa_snapshot[12][52] , \sa_snapshot[12].r.part1[20] );
tran (\sa_snapshot[12][52] , \sa_snapshot[12].f.unused[2] );
tran (\sa_snapshot[12][51] , \sa_snapshot[12].r.part1[19] );
tran (\sa_snapshot[12][51] , \sa_snapshot[12].f.unused[1] );
tran (\sa_snapshot[12][50] , \sa_snapshot[12].r.part1[18] );
tran (\sa_snapshot[12][50] , \sa_snapshot[12].f.unused[0] );
tran (\sa_snapshot[12][49] , \sa_snapshot[12].r.part1[17] );
tran (\sa_snapshot[12][49] , \sa_snapshot[12].f.upper[17] );
tran (\sa_snapshot[12][48] , \sa_snapshot[12].r.part1[16] );
tran (\sa_snapshot[12][48] , \sa_snapshot[12].f.upper[16] );
tran (\sa_snapshot[12][47] , \sa_snapshot[12].r.part1[15] );
tran (\sa_snapshot[12][47] , \sa_snapshot[12].f.upper[15] );
tran (\sa_snapshot[12][46] , \sa_snapshot[12].r.part1[14] );
tran (\sa_snapshot[12][46] , \sa_snapshot[12].f.upper[14] );
tran (\sa_snapshot[12][45] , \sa_snapshot[12].r.part1[13] );
tran (\sa_snapshot[12][45] , \sa_snapshot[12].f.upper[13] );
tran (\sa_snapshot[12][44] , \sa_snapshot[12].r.part1[12] );
tran (\sa_snapshot[12][44] , \sa_snapshot[12].f.upper[12] );
tran (\sa_snapshot[12][43] , \sa_snapshot[12].r.part1[11] );
tran (\sa_snapshot[12][43] , \sa_snapshot[12].f.upper[11] );
tran (\sa_snapshot[12][42] , \sa_snapshot[12].r.part1[10] );
tran (\sa_snapshot[12][42] , \sa_snapshot[12].f.upper[10] );
tran (\sa_snapshot[12][41] , \sa_snapshot[12].r.part1[9] );
tran (\sa_snapshot[12][41] , \sa_snapshot[12].f.upper[9] );
tran (\sa_snapshot[12][40] , \sa_snapshot[12].r.part1[8] );
tran (\sa_snapshot[12][40] , \sa_snapshot[12].f.upper[8] );
tran (\sa_snapshot[12][39] , \sa_snapshot[12].r.part1[7] );
tran (\sa_snapshot[12][39] , \sa_snapshot[12].f.upper[7] );
tran (\sa_snapshot[12][38] , \sa_snapshot[12].r.part1[6] );
tran (\sa_snapshot[12][38] , \sa_snapshot[12].f.upper[6] );
tran (\sa_snapshot[12][37] , \sa_snapshot[12].r.part1[5] );
tran (\sa_snapshot[12][37] , \sa_snapshot[12].f.upper[5] );
tran (\sa_snapshot[12][36] , \sa_snapshot[12].r.part1[4] );
tran (\sa_snapshot[12][36] , \sa_snapshot[12].f.upper[4] );
tran (\sa_snapshot[12][35] , \sa_snapshot[12].r.part1[3] );
tran (\sa_snapshot[12][35] , \sa_snapshot[12].f.upper[3] );
tran (\sa_snapshot[12][34] , \sa_snapshot[12].r.part1[2] );
tran (\sa_snapshot[12][34] , \sa_snapshot[12].f.upper[2] );
tran (\sa_snapshot[12][33] , \sa_snapshot[12].r.part1[1] );
tran (\sa_snapshot[12][33] , \sa_snapshot[12].f.upper[1] );
tran (\sa_snapshot[12][32] , \sa_snapshot[12].r.part1[0] );
tran (\sa_snapshot[12][32] , \sa_snapshot[12].f.upper[0] );
tran (\sa_snapshot[12][31] , \sa_snapshot[12].r.part0[31] );
tran (\sa_snapshot[12][31] , \sa_snapshot[12].f.lower[31] );
tran (\sa_snapshot[12][30] , \sa_snapshot[12].r.part0[30] );
tran (\sa_snapshot[12][30] , \sa_snapshot[12].f.lower[30] );
tran (\sa_snapshot[12][29] , \sa_snapshot[12].r.part0[29] );
tran (\sa_snapshot[12][29] , \sa_snapshot[12].f.lower[29] );
tran (\sa_snapshot[12][28] , \sa_snapshot[12].r.part0[28] );
tran (\sa_snapshot[12][28] , \sa_snapshot[12].f.lower[28] );
tran (\sa_snapshot[12][27] , \sa_snapshot[12].r.part0[27] );
tran (\sa_snapshot[12][27] , \sa_snapshot[12].f.lower[27] );
tran (\sa_snapshot[12][26] , \sa_snapshot[12].r.part0[26] );
tran (\sa_snapshot[12][26] , \sa_snapshot[12].f.lower[26] );
tran (\sa_snapshot[12][25] , \sa_snapshot[12].r.part0[25] );
tran (\sa_snapshot[12][25] , \sa_snapshot[12].f.lower[25] );
tran (\sa_snapshot[12][24] , \sa_snapshot[12].r.part0[24] );
tran (\sa_snapshot[12][24] , \sa_snapshot[12].f.lower[24] );
tran (\sa_snapshot[12][23] , \sa_snapshot[12].r.part0[23] );
tran (\sa_snapshot[12][23] , \sa_snapshot[12].f.lower[23] );
tran (\sa_snapshot[12][22] , \sa_snapshot[12].r.part0[22] );
tran (\sa_snapshot[12][22] , \sa_snapshot[12].f.lower[22] );
tran (\sa_snapshot[12][21] , \sa_snapshot[12].r.part0[21] );
tran (\sa_snapshot[12][21] , \sa_snapshot[12].f.lower[21] );
tran (\sa_snapshot[12][20] , \sa_snapshot[12].r.part0[20] );
tran (\sa_snapshot[12][20] , \sa_snapshot[12].f.lower[20] );
tran (\sa_snapshot[12][19] , \sa_snapshot[12].r.part0[19] );
tran (\sa_snapshot[12][19] , \sa_snapshot[12].f.lower[19] );
tran (\sa_snapshot[12][18] , \sa_snapshot[12].r.part0[18] );
tran (\sa_snapshot[12][18] , \sa_snapshot[12].f.lower[18] );
tran (\sa_snapshot[12][17] , \sa_snapshot[12].r.part0[17] );
tran (\sa_snapshot[12][17] , \sa_snapshot[12].f.lower[17] );
tran (\sa_snapshot[12][16] , \sa_snapshot[12].r.part0[16] );
tran (\sa_snapshot[12][16] , \sa_snapshot[12].f.lower[16] );
tran (\sa_snapshot[12][15] , \sa_snapshot[12].r.part0[15] );
tran (\sa_snapshot[12][15] , \sa_snapshot[12].f.lower[15] );
tran (\sa_snapshot[12][14] , \sa_snapshot[12].r.part0[14] );
tran (\sa_snapshot[12][14] , \sa_snapshot[12].f.lower[14] );
tran (\sa_snapshot[12][13] , \sa_snapshot[12].r.part0[13] );
tran (\sa_snapshot[12][13] , \sa_snapshot[12].f.lower[13] );
tran (\sa_snapshot[12][12] , \sa_snapshot[12].r.part0[12] );
tran (\sa_snapshot[12][12] , \sa_snapshot[12].f.lower[12] );
tran (\sa_snapshot[12][11] , \sa_snapshot[12].r.part0[11] );
tran (\sa_snapshot[12][11] , \sa_snapshot[12].f.lower[11] );
tran (\sa_snapshot[12][10] , \sa_snapshot[12].r.part0[10] );
tran (\sa_snapshot[12][10] , \sa_snapshot[12].f.lower[10] );
tran (\sa_snapshot[12][9] , \sa_snapshot[12].r.part0[9] );
tran (\sa_snapshot[12][9] , \sa_snapshot[12].f.lower[9] );
tran (\sa_snapshot[12][8] , \sa_snapshot[12].r.part0[8] );
tran (\sa_snapshot[12][8] , \sa_snapshot[12].f.lower[8] );
tran (\sa_snapshot[12][7] , \sa_snapshot[12].r.part0[7] );
tran (\sa_snapshot[12][7] , \sa_snapshot[12].f.lower[7] );
tran (\sa_snapshot[12][6] , \sa_snapshot[12].r.part0[6] );
tran (\sa_snapshot[12][6] , \sa_snapshot[12].f.lower[6] );
tran (\sa_snapshot[12][5] , \sa_snapshot[12].r.part0[5] );
tran (\sa_snapshot[12][5] , \sa_snapshot[12].f.lower[5] );
tran (\sa_snapshot[12][4] , \sa_snapshot[12].r.part0[4] );
tran (\sa_snapshot[12][4] , \sa_snapshot[12].f.lower[4] );
tran (\sa_snapshot[12][3] , \sa_snapshot[12].r.part0[3] );
tran (\sa_snapshot[12][3] , \sa_snapshot[12].f.lower[3] );
tran (\sa_snapshot[12][2] , \sa_snapshot[12].r.part0[2] );
tran (\sa_snapshot[12][2] , \sa_snapshot[12].f.lower[2] );
tran (\sa_snapshot[12][1] , \sa_snapshot[12].r.part0[1] );
tran (\sa_snapshot[12][1] , \sa_snapshot[12].f.lower[1] );
tran (\sa_snapshot[12][0] , \sa_snapshot[12].r.part0[0] );
tran (\sa_snapshot[12][0] , \sa_snapshot[12].f.lower[0] );
tran (\sa_snapshot[11][63] , \sa_snapshot[11].r.part1[31] );
tran (\sa_snapshot[11][63] , \sa_snapshot[11].f.unused[13] );
tran (\sa_snapshot[11][62] , \sa_snapshot[11].r.part1[30] );
tran (\sa_snapshot[11][62] , \sa_snapshot[11].f.unused[12] );
tran (\sa_snapshot[11][61] , \sa_snapshot[11].r.part1[29] );
tran (\sa_snapshot[11][61] , \sa_snapshot[11].f.unused[11] );
tran (\sa_snapshot[11][60] , \sa_snapshot[11].r.part1[28] );
tran (\sa_snapshot[11][60] , \sa_snapshot[11].f.unused[10] );
tran (\sa_snapshot[11][59] , \sa_snapshot[11].r.part1[27] );
tran (\sa_snapshot[11][59] , \sa_snapshot[11].f.unused[9] );
tran (\sa_snapshot[11][58] , \sa_snapshot[11].r.part1[26] );
tran (\sa_snapshot[11][58] , \sa_snapshot[11].f.unused[8] );
tran (\sa_snapshot[11][57] , \sa_snapshot[11].r.part1[25] );
tran (\sa_snapshot[11][57] , \sa_snapshot[11].f.unused[7] );
tran (\sa_snapshot[11][56] , \sa_snapshot[11].r.part1[24] );
tran (\sa_snapshot[11][56] , \sa_snapshot[11].f.unused[6] );
tran (\sa_snapshot[11][55] , \sa_snapshot[11].r.part1[23] );
tran (\sa_snapshot[11][55] , \sa_snapshot[11].f.unused[5] );
tran (\sa_snapshot[11][54] , \sa_snapshot[11].r.part1[22] );
tran (\sa_snapshot[11][54] , \sa_snapshot[11].f.unused[4] );
tran (\sa_snapshot[11][53] , \sa_snapshot[11].r.part1[21] );
tran (\sa_snapshot[11][53] , \sa_snapshot[11].f.unused[3] );
tran (\sa_snapshot[11][52] , \sa_snapshot[11].r.part1[20] );
tran (\sa_snapshot[11][52] , \sa_snapshot[11].f.unused[2] );
tran (\sa_snapshot[11][51] , \sa_snapshot[11].r.part1[19] );
tran (\sa_snapshot[11][51] , \sa_snapshot[11].f.unused[1] );
tran (\sa_snapshot[11][50] , \sa_snapshot[11].r.part1[18] );
tran (\sa_snapshot[11][50] , \sa_snapshot[11].f.unused[0] );
tran (\sa_snapshot[11][49] , \sa_snapshot[11].r.part1[17] );
tran (\sa_snapshot[11][49] , \sa_snapshot[11].f.upper[17] );
tran (\sa_snapshot[11][48] , \sa_snapshot[11].r.part1[16] );
tran (\sa_snapshot[11][48] , \sa_snapshot[11].f.upper[16] );
tran (\sa_snapshot[11][47] , \sa_snapshot[11].r.part1[15] );
tran (\sa_snapshot[11][47] , \sa_snapshot[11].f.upper[15] );
tran (\sa_snapshot[11][46] , \sa_snapshot[11].r.part1[14] );
tran (\sa_snapshot[11][46] , \sa_snapshot[11].f.upper[14] );
tran (\sa_snapshot[11][45] , \sa_snapshot[11].r.part1[13] );
tran (\sa_snapshot[11][45] , \sa_snapshot[11].f.upper[13] );
tran (\sa_snapshot[11][44] , \sa_snapshot[11].r.part1[12] );
tran (\sa_snapshot[11][44] , \sa_snapshot[11].f.upper[12] );
tran (\sa_snapshot[11][43] , \sa_snapshot[11].r.part1[11] );
tran (\sa_snapshot[11][43] , \sa_snapshot[11].f.upper[11] );
tran (\sa_snapshot[11][42] , \sa_snapshot[11].r.part1[10] );
tran (\sa_snapshot[11][42] , \sa_snapshot[11].f.upper[10] );
tran (\sa_snapshot[11][41] , \sa_snapshot[11].r.part1[9] );
tran (\sa_snapshot[11][41] , \sa_snapshot[11].f.upper[9] );
tran (\sa_snapshot[11][40] , \sa_snapshot[11].r.part1[8] );
tran (\sa_snapshot[11][40] , \sa_snapshot[11].f.upper[8] );
tran (\sa_snapshot[11][39] , \sa_snapshot[11].r.part1[7] );
tran (\sa_snapshot[11][39] , \sa_snapshot[11].f.upper[7] );
tran (\sa_snapshot[11][38] , \sa_snapshot[11].r.part1[6] );
tran (\sa_snapshot[11][38] , \sa_snapshot[11].f.upper[6] );
tran (\sa_snapshot[11][37] , \sa_snapshot[11].r.part1[5] );
tran (\sa_snapshot[11][37] , \sa_snapshot[11].f.upper[5] );
tran (\sa_snapshot[11][36] , \sa_snapshot[11].r.part1[4] );
tran (\sa_snapshot[11][36] , \sa_snapshot[11].f.upper[4] );
tran (\sa_snapshot[11][35] , \sa_snapshot[11].r.part1[3] );
tran (\sa_snapshot[11][35] , \sa_snapshot[11].f.upper[3] );
tran (\sa_snapshot[11][34] , \sa_snapshot[11].r.part1[2] );
tran (\sa_snapshot[11][34] , \sa_snapshot[11].f.upper[2] );
tran (\sa_snapshot[11][33] , \sa_snapshot[11].r.part1[1] );
tran (\sa_snapshot[11][33] , \sa_snapshot[11].f.upper[1] );
tran (\sa_snapshot[11][32] , \sa_snapshot[11].r.part1[0] );
tran (\sa_snapshot[11][32] , \sa_snapshot[11].f.upper[0] );
tran (\sa_snapshot[11][31] , \sa_snapshot[11].r.part0[31] );
tran (\sa_snapshot[11][31] , \sa_snapshot[11].f.lower[31] );
tran (\sa_snapshot[11][30] , \sa_snapshot[11].r.part0[30] );
tran (\sa_snapshot[11][30] , \sa_snapshot[11].f.lower[30] );
tran (\sa_snapshot[11][29] , \sa_snapshot[11].r.part0[29] );
tran (\sa_snapshot[11][29] , \sa_snapshot[11].f.lower[29] );
tran (\sa_snapshot[11][28] , \sa_snapshot[11].r.part0[28] );
tran (\sa_snapshot[11][28] , \sa_snapshot[11].f.lower[28] );
tran (\sa_snapshot[11][27] , \sa_snapshot[11].r.part0[27] );
tran (\sa_snapshot[11][27] , \sa_snapshot[11].f.lower[27] );
tran (\sa_snapshot[11][26] , \sa_snapshot[11].r.part0[26] );
tran (\sa_snapshot[11][26] , \sa_snapshot[11].f.lower[26] );
tran (\sa_snapshot[11][25] , \sa_snapshot[11].r.part0[25] );
tran (\sa_snapshot[11][25] , \sa_snapshot[11].f.lower[25] );
tran (\sa_snapshot[11][24] , \sa_snapshot[11].r.part0[24] );
tran (\sa_snapshot[11][24] , \sa_snapshot[11].f.lower[24] );
tran (\sa_snapshot[11][23] , \sa_snapshot[11].r.part0[23] );
tran (\sa_snapshot[11][23] , \sa_snapshot[11].f.lower[23] );
tran (\sa_snapshot[11][22] , \sa_snapshot[11].r.part0[22] );
tran (\sa_snapshot[11][22] , \sa_snapshot[11].f.lower[22] );
tran (\sa_snapshot[11][21] , \sa_snapshot[11].r.part0[21] );
tran (\sa_snapshot[11][21] , \sa_snapshot[11].f.lower[21] );
tran (\sa_snapshot[11][20] , \sa_snapshot[11].r.part0[20] );
tran (\sa_snapshot[11][20] , \sa_snapshot[11].f.lower[20] );
tran (\sa_snapshot[11][19] , \sa_snapshot[11].r.part0[19] );
tran (\sa_snapshot[11][19] , \sa_snapshot[11].f.lower[19] );
tran (\sa_snapshot[11][18] , \sa_snapshot[11].r.part0[18] );
tran (\sa_snapshot[11][18] , \sa_snapshot[11].f.lower[18] );
tran (\sa_snapshot[11][17] , \sa_snapshot[11].r.part0[17] );
tran (\sa_snapshot[11][17] , \sa_snapshot[11].f.lower[17] );
tran (\sa_snapshot[11][16] , \sa_snapshot[11].r.part0[16] );
tran (\sa_snapshot[11][16] , \sa_snapshot[11].f.lower[16] );
tran (\sa_snapshot[11][15] , \sa_snapshot[11].r.part0[15] );
tran (\sa_snapshot[11][15] , \sa_snapshot[11].f.lower[15] );
tran (\sa_snapshot[11][14] , \sa_snapshot[11].r.part0[14] );
tran (\sa_snapshot[11][14] , \sa_snapshot[11].f.lower[14] );
tran (\sa_snapshot[11][13] , \sa_snapshot[11].r.part0[13] );
tran (\sa_snapshot[11][13] , \sa_snapshot[11].f.lower[13] );
tran (\sa_snapshot[11][12] , \sa_snapshot[11].r.part0[12] );
tran (\sa_snapshot[11][12] , \sa_snapshot[11].f.lower[12] );
tran (\sa_snapshot[11][11] , \sa_snapshot[11].r.part0[11] );
tran (\sa_snapshot[11][11] , \sa_snapshot[11].f.lower[11] );
tran (\sa_snapshot[11][10] , \sa_snapshot[11].r.part0[10] );
tran (\sa_snapshot[11][10] , \sa_snapshot[11].f.lower[10] );
tran (\sa_snapshot[11][9] , \sa_snapshot[11].r.part0[9] );
tran (\sa_snapshot[11][9] , \sa_snapshot[11].f.lower[9] );
tran (\sa_snapshot[11][8] , \sa_snapshot[11].r.part0[8] );
tran (\sa_snapshot[11][8] , \sa_snapshot[11].f.lower[8] );
tran (\sa_snapshot[11][7] , \sa_snapshot[11].r.part0[7] );
tran (\sa_snapshot[11][7] , \sa_snapshot[11].f.lower[7] );
tran (\sa_snapshot[11][6] , \sa_snapshot[11].r.part0[6] );
tran (\sa_snapshot[11][6] , \sa_snapshot[11].f.lower[6] );
tran (\sa_snapshot[11][5] , \sa_snapshot[11].r.part0[5] );
tran (\sa_snapshot[11][5] , \sa_snapshot[11].f.lower[5] );
tran (\sa_snapshot[11][4] , \sa_snapshot[11].r.part0[4] );
tran (\sa_snapshot[11][4] , \sa_snapshot[11].f.lower[4] );
tran (\sa_snapshot[11][3] , \sa_snapshot[11].r.part0[3] );
tran (\sa_snapshot[11][3] , \sa_snapshot[11].f.lower[3] );
tran (\sa_snapshot[11][2] , \sa_snapshot[11].r.part0[2] );
tran (\sa_snapshot[11][2] , \sa_snapshot[11].f.lower[2] );
tran (\sa_snapshot[11][1] , \sa_snapshot[11].r.part0[1] );
tran (\sa_snapshot[11][1] , \sa_snapshot[11].f.lower[1] );
tran (\sa_snapshot[11][0] , \sa_snapshot[11].r.part0[0] );
tran (\sa_snapshot[11][0] , \sa_snapshot[11].f.lower[0] );
tran (\sa_snapshot[10][63] , \sa_snapshot[10].r.part1[31] );
tran (\sa_snapshot[10][63] , \sa_snapshot[10].f.unused[13] );
tran (\sa_snapshot[10][62] , \sa_snapshot[10].r.part1[30] );
tran (\sa_snapshot[10][62] , \sa_snapshot[10].f.unused[12] );
tran (\sa_snapshot[10][61] , \sa_snapshot[10].r.part1[29] );
tran (\sa_snapshot[10][61] , \sa_snapshot[10].f.unused[11] );
tran (\sa_snapshot[10][60] , \sa_snapshot[10].r.part1[28] );
tran (\sa_snapshot[10][60] , \sa_snapshot[10].f.unused[10] );
tran (\sa_snapshot[10][59] , \sa_snapshot[10].r.part1[27] );
tran (\sa_snapshot[10][59] , \sa_snapshot[10].f.unused[9] );
tran (\sa_snapshot[10][58] , \sa_snapshot[10].r.part1[26] );
tran (\sa_snapshot[10][58] , \sa_snapshot[10].f.unused[8] );
tran (\sa_snapshot[10][57] , \sa_snapshot[10].r.part1[25] );
tran (\sa_snapshot[10][57] , \sa_snapshot[10].f.unused[7] );
tran (\sa_snapshot[10][56] , \sa_snapshot[10].r.part1[24] );
tran (\sa_snapshot[10][56] , \sa_snapshot[10].f.unused[6] );
tran (\sa_snapshot[10][55] , \sa_snapshot[10].r.part1[23] );
tran (\sa_snapshot[10][55] , \sa_snapshot[10].f.unused[5] );
tran (\sa_snapshot[10][54] , \sa_snapshot[10].r.part1[22] );
tran (\sa_snapshot[10][54] , \sa_snapshot[10].f.unused[4] );
tran (\sa_snapshot[10][53] , \sa_snapshot[10].r.part1[21] );
tran (\sa_snapshot[10][53] , \sa_snapshot[10].f.unused[3] );
tran (\sa_snapshot[10][52] , \sa_snapshot[10].r.part1[20] );
tran (\sa_snapshot[10][52] , \sa_snapshot[10].f.unused[2] );
tran (\sa_snapshot[10][51] , \sa_snapshot[10].r.part1[19] );
tran (\sa_snapshot[10][51] , \sa_snapshot[10].f.unused[1] );
tran (\sa_snapshot[10][50] , \sa_snapshot[10].r.part1[18] );
tran (\sa_snapshot[10][50] , \sa_snapshot[10].f.unused[0] );
tran (\sa_snapshot[10][49] , \sa_snapshot[10].r.part1[17] );
tran (\sa_snapshot[10][49] , \sa_snapshot[10].f.upper[17] );
tran (\sa_snapshot[10][48] , \sa_snapshot[10].r.part1[16] );
tran (\sa_snapshot[10][48] , \sa_snapshot[10].f.upper[16] );
tran (\sa_snapshot[10][47] , \sa_snapshot[10].r.part1[15] );
tran (\sa_snapshot[10][47] , \sa_snapshot[10].f.upper[15] );
tran (\sa_snapshot[10][46] , \sa_snapshot[10].r.part1[14] );
tran (\sa_snapshot[10][46] , \sa_snapshot[10].f.upper[14] );
tran (\sa_snapshot[10][45] , \sa_snapshot[10].r.part1[13] );
tran (\sa_snapshot[10][45] , \sa_snapshot[10].f.upper[13] );
tran (\sa_snapshot[10][44] , \sa_snapshot[10].r.part1[12] );
tran (\sa_snapshot[10][44] , \sa_snapshot[10].f.upper[12] );
tran (\sa_snapshot[10][43] , \sa_snapshot[10].r.part1[11] );
tran (\sa_snapshot[10][43] , \sa_snapshot[10].f.upper[11] );
tran (\sa_snapshot[10][42] , \sa_snapshot[10].r.part1[10] );
tran (\sa_snapshot[10][42] , \sa_snapshot[10].f.upper[10] );
tran (\sa_snapshot[10][41] , \sa_snapshot[10].r.part1[9] );
tran (\sa_snapshot[10][41] , \sa_snapshot[10].f.upper[9] );
tran (\sa_snapshot[10][40] , \sa_snapshot[10].r.part1[8] );
tran (\sa_snapshot[10][40] , \sa_snapshot[10].f.upper[8] );
tran (\sa_snapshot[10][39] , \sa_snapshot[10].r.part1[7] );
tran (\sa_snapshot[10][39] , \sa_snapshot[10].f.upper[7] );
tran (\sa_snapshot[10][38] , \sa_snapshot[10].r.part1[6] );
tran (\sa_snapshot[10][38] , \sa_snapshot[10].f.upper[6] );
tran (\sa_snapshot[10][37] , \sa_snapshot[10].r.part1[5] );
tran (\sa_snapshot[10][37] , \sa_snapshot[10].f.upper[5] );
tran (\sa_snapshot[10][36] , \sa_snapshot[10].r.part1[4] );
tran (\sa_snapshot[10][36] , \sa_snapshot[10].f.upper[4] );
tran (\sa_snapshot[10][35] , \sa_snapshot[10].r.part1[3] );
tran (\sa_snapshot[10][35] , \sa_snapshot[10].f.upper[3] );
tran (\sa_snapshot[10][34] , \sa_snapshot[10].r.part1[2] );
tran (\sa_snapshot[10][34] , \sa_snapshot[10].f.upper[2] );
tran (\sa_snapshot[10][33] , \sa_snapshot[10].r.part1[1] );
tran (\sa_snapshot[10][33] , \sa_snapshot[10].f.upper[1] );
tran (\sa_snapshot[10][32] , \sa_snapshot[10].r.part1[0] );
tran (\sa_snapshot[10][32] , \sa_snapshot[10].f.upper[0] );
tran (\sa_snapshot[10][31] , \sa_snapshot[10].r.part0[31] );
tran (\sa_snapshot[10][31] , \sa_snapshot[10].f.lower[31] );
tran (\sa_snapshot[10][30] , \sa_snapshot[10].r.part0[30] );
tran (\sa_snapshot[10][30] , \sa_snapshot[10].f.lower[30] );
tran (\sa_snapshot[10][29] , \sa_snapshot[10].r.part0[29] );
tran (\sa_snapshot[10][29] , \sa_snapshot[10].f.lower[29] );
tran (\sa_snapshot[10][28] , \sa_snapshot[10].r.part0[28] );
tran (\sa_snapshot[10][28] , \sa_snapshot[10].f.lower[28] );
tran (\sa_snapshot[10][27] , \sa_snapshot[10].r.part0[27] );
tran (\sa_snapshot[10][27] , \sa_snapshot[10].f.lower[27] );
tran (\sa_snapshot[10][26] , \sa_snapshot[10].r.part0[26] );
tran (\sa_snapshot[10][26] , \sa_snapshot[10].f.lower[26] );
tran (\sa_snapshot[10][25] , \sa_snapshot[10].r.part0[25] );
tran (\sa_snapshot[10][25] , \sa_snapshot[10].f.lower[25] );
tran (\sa_snapshot[10][24] , \sa_snapshot[10].r.part0[24] );
tran (\sa_snapshot[10][24] , \sa_snapshot[10].f.lower[24] );
tran (\sa_snapshot[10][23] , \sa_snapshot[10].r.part0[23] );
tran (\sa_snapshot[10][23] , \sa_snapshot[10].f.lower[23] );
tran (\sa_snapshot[10][22] , \sa_snapshot[10].r.part0[22] );
tran (\sa_snapshot[10][22] , \sa_snapshot[10].f.lower[22] );
tran (\sa_snapshot[10][21] , \sa_snapshot[10].r.part0[21] );
tran (\sa_snapshot[10][21] , \sa_snapshot[10].f.lower[21] );
tran (\sa_snapshot[10][20] , \sa_snapshot[10].r.part0[20] );
tran (\sa_snapshot[10][20] , \sa_snapshot[10].f.lower[20] );
tran (\sa_snapshot[10][19] , \sa_snapshot[10].r.part0[19] );
tran (\sa_snapshot[10][19] , \sa_snapshot[10].f.lower[19] );
tran (\sa_snapshot[10][18] , \sa_snapshot[10].r.part0[18] );
tran (\sa_snapshot[10][18] , \sa_snapshot[10].f.lower[18] );
tran (\sa_snapshot[10][17] , \sa_snapshot[10].r.part0[17] );
tran (\sa_snapshot[10][17] , \sa_snapshot[10].f.lower[17] );
tran (\sa_snapshot[10][16] , \sa_snapshot[10].r.part0[16] );
tran (\sa_snapshot[10][16] , \sa_snapshot[10].f.lower[16] );
tran (\sa_snapshot[10][15] , \sa_snapshot[10].r.part0[15] );
tran (\sa_snapshot[10][15] , \sa_snapshot[10].f.lower[15] );
tran (\sa_snapshot[10][14] , \sa_snapshot[10].r.part0[14] );
tran (\sa_snapshot[10][14] , \sa_snapshot[10].f.lower[14] );
tran (\sa_snapshot[10][13] , \sa_snapshot[10].r.part0[13] );
tran (\sa_snapshot[10][13] , \sa_snapshot[10].f.lower[13] );
tran (\sa_snapshot[10][12] , \sa_snapshot[10].r.part0[12] );
tran (\sa_snapshot[10][12] , \sa_snapshot[10].f.lower[12] );
tran (\sa_snapshot[10][11] , \sa_snapshot[10].r.part0[11] );
tran (\sa_snapshot[10][11] , \sa_snapshot[10].f.lower[11] );
tran (\sa_snapshot[10][10] , \sa_snapshot[10].r.part0[10] );
tran (\sa_snapshot[10][10] , \sa_snapshot[10].f.lower[10] );
tran (\sa_snapshot[10][9] , \sa_snapshot[10].r.part0[9] );
tran (\sa_snapshot[10][9] , \sa_snapshot[10].f.lower[9] );
tran (\sa_snapshot[10][8] , \sa_snapshot[10].r.part0[8] );
tran (\sa_snapshot[10][8] , \sa_snapshot[10].f.lower[8] );
tran (\sa_snapshot[10][7] , \sa_snapshot[10].r.part0[7] );
tran (\sa_snapshot[10][7] , \sa_snapshot[10].f.lower[7] );
tran (\sa_snapshot[10][6] , \sa_snapshot[10].r.part0[6] );
tran (\sa_snapshot[10][6] , \sa_snapshot[10].f.lower[6] );
tran (\sa_snapshot[10][5] , \sa_snapshot[10].r.part0[5] );
tran (\sa_snapshot[10][5] , \sa_snapshot[10].f.lower[5] );
tran (\sa_snapshot[10][4] , \sa_snapshot[10].r.part0[4] );
tran (\sa_snapshot[10][4] , \sa_snapshot[10].f.lower[4] );
tran (\sa_snapshot[10][3] , \sa_snapshot[10].r.part0[3] );
tran (\sa_snapshot[10][3] , \sa_snapshot[10].f.lower[3] );
tran (\sa_snapshot[10][2] , \sa_snapshot[10].r.part0[2] );
tran (\sa_snapshot[10][2] , \sa_snapshot[10].f.lower[2] );
tran (\sa_snapshot[10][1] , \sa_snapshot[10].r.part0[1] );
tran (\sa_snapshot[10][1] , \sa_snapshot[10].f.lower[1] );
tran (\sa_snapshot[10][0] , \sa_snapshot[10].r.part0[0] );
tran (\sa_snapshot[10][0] , \sa_snapshot[10].f.lower[0] );
tran (\sa_snapshot[9][63] , \sa_snapshot[9].r.part1[31] );
tran (\sa_snapshot[9][63] , \sa_snapshot[9].f.unused[13] );
tran (\sa_snapshot[9][62] , \sa_snapshot[9].r.part1[30] );
tran (\sa_snapshot[9][62] , \sa_snapshot[9].f.unused[12] );
tran (\sa_snapshot[9][61] , \sa_snapshot[9].r.part1[29] );
tran (\sa_snapshot[9][61] , \sa_snapshot[9].f.unused[11] );
tran (\sa_snapshot[9][60] , \sa_snapshot[9].r.part1[28] );
tran (\sa_snapshot[9][60] , \sa_snapshot[9].f.unused[10] );
tran (\sa_snapshot[9][59] , \sa_snapshot[9].r.part1[27] );
tran (\sa_snapshot[9][59] , \sa_snapshot[9].f.unused[9] );
tran (\sa_snapshot[9][58] , \sa_snapshot[9].r.part1[26] );
tran (\sa_snapshot[9][58] , \sa_snapshot[9].f.unused[8] );
tran (\sa_snapshot[9][57] , \sa_snapshot[9].r.part1[25] );
tran (\sa_snapshot[9][57] , \sa_snapshot[9].f.unused[7] );
tran (\sa_snapshot[9][56] , \sa_snapshot[9].r.part1[24] );
tran (\sa_snapshot[9][56] , \sa_snapshot[9].f.unused[6] );
tran (\sa_snapshot[9][55] , \sa_snapshot[9].r.part1[23] );
tran (\sa_snapshot[9][55] , \sa_snapshot[9].f.unused[5] );
tran (\sa_snapshot[9][54] , \sa_snapshot[9].r.part1[22] );
tran (\sa_snapshot[9][54] , \sa_snapshot[9].f.unused[4] );
tran (\sa_snapshot[9][53] , \sa_snapshot[9].r.part1[21] );
tran (\sa_snapshot[9][53] , \sa_snapshot[9].f.unused[3] );
tran (\sa_snapshot[9][52] , \sa_snapshot[9].r.part1[20] );
tran (\sa_snapshot[9][52] , \sa_snapshot[9].f.unused[2] );
tran (\sa_snapshot[9][51] , \sa_snapshot[9].r.part1[19] );
tran (\sa_snapshot[9][51] , \sa_snapshot[9].f.unused[1] );
tran (\sa_snapshot[9][50] , \sa_snapshot[9].r.part1[18] );
tran (\sa_snapshot[9][50] , \sa_snapshot[9].f.unused[0] );
tran (\sa_snapshot[9][49] , \sa_snapshot[9].r.part1[17] );
tran (\sa_snapshot[9][49] , \sa_snapshot[9].f.upper[17] );
tran (\sa_snapshot[9][48] , \sa_snapshot[9].r.part1[16] );
tran (\sa_snapshot[9][48] , \sa_snapshot[9].f.upper[16] );
tran (\sa_snapshot[9][47] , \sa_snapshot[9].r.part1[15] );
tran (\sa_snapshot[9][47] , \sa_snapshot[9].f.upper[15] );
tran (\sa_snapshot[9][46] , \sa_snapshot[9].r.part1[14] );
tran (\sa_snapshot[9][46] , \sa_snapshot[9].f.upper[14] );
tran (\sa_snapshot[9][45] , \sa_snapshot[9].r.part1[13] );
tran (\sa_snapshot[9][45] , \sa_snapshot[9].f.upper[13] );
tran (\sa_snapshot[9][44] , \sa_snapshot[9].r.part1[12] );
tran (\sa_snapshot[9][44] , \sa_snapshot[9].f.upper[12] );
tran (\sa_snapshot[9][43] , \sa_snapshot[9].r.part1[11] );
tran (\sa_snapshot[9][43] , \sa_snapshot[9].f.upper[11] );
tran (\sa_snapshot[9][42] , \sa_snapshot[9].r.part1[10] );
tran (\sa_snapshot[9][42] , \sa_snapshot[9].f.upper[10] );
tran (\sa_snapshot[9][41] , \sa_snapshot[9].r.part1[9] );
tran (\sa_snapshot[9][41] , \sa_snapshot[9].f.upper[9] );
tran (\sa_snapshot[9][40] , \sa_snapshot[9].r.part1[8] );
tran (\sa_snapshot[9][40] , \sa_snapshot[9].f.upper[8] );
tran (\sa_snapshot[9][39] , \sa_snapshot[9].r.part1[7] );
tran (\sa_snapshot[9][39] , \sa_snapshot[9].f.upper[7] );
tran (\sa_snapshot[9][38] , \sa_snapshot[9].r.part1[6] );
tran (\sa_snapshot[9][38] , \sa_snapshot[9].f.upper[6] );
tran (\sa_snapshot[9][37] , \sa_snapshot[9].r.part1[5] );
tran (\sa_snapshot[9][37] , \sa_snapshot[9].f.upper[5] );
tran (\sa_snapshot[9][36] , \sa_snapshot[9].r.part1[4] );
tran (\sa_snapshot[9][36] , \sa_snapshot[9].f.upper[4] );
tran (\sa_snapshot[9][35] , \sa_snapshot[9].r.part1[3] );
tran (\sa_snapshot[9][35] , \sa_snapshot[9].f.upper[3] );
tran (\sa_snapshot[9][34] , \sa_snapshot[9].r.part1[2] );
tran (\sa_snapshot[9][34] , \sa_snapshot[9].f.upper[2] );
tran (\sa_snapshot[9][33] , \sa_snapshot[9].r.part1[1] );
tran (\sa_snapshot[9][33] , \sa_snapshot[9].f.upper[1] );
tran (\sa_snapshot[9][32] , \sa_snapshot[9].r.part1[0] );
tran (\sa_snapshot[9][32] , \sa_snapshot[9].f.upper[0] );
tran (\sa_snapshot[9][31] , \sa_snapshot[9].r.part0[31] );
tran (\sa_snapshot[9][31] , \sa_snapshot[9].f.lower[31] );
tran (\sa_snapshot[9][30] , \sa_snapshot[9].r.part0[30] );
tran (\sa_snapshot[9][30] , \sa_snapshot[9].f.lower[30] );
tran (\sa_snapshot[9][29] , \sa_snapshot[9].r.part0[29] );
tran (\sa_snapshot[9][29] , \sa_snapshot[9].f.lower[29] );
tran (\sa_snapshot[9][28] , \sa_snapshot[9].r.part0[28] );
tran (\sa_snapshot[9][28] , \sa_snapshot[9].f.lower[28] );
tran (\sa_snapshot[9][27] , \sa_snapshot[9].r.part0[27] );
tran (\sa_snapshot[9][27] , \sa_snapshot[9].f.lower[27] );
tran (\sa_snapshot[9][26] , \sa_snapshot[9].r.part0[26] );
tran (\sa_snapshot[9][26] , \sa_snapshot[9].f.lower[26] );
tran (\sa_snapshot[9][25] , \sa_snapshot[9].r.part0[25] );
tran (\sa_snapshot[9][25] , \sa_snapshot[9].f.lower[25] );
tran (\sa_snapshot[9][24] , \sa_snapshot[9].r.part0[24] );
tran (\sa_snapshot[9][24] , \sa_snapshot[9].f.lower[24] );
tran (\sa_snapshot[9][23] , \sa_snapshot[9].r.part0[23] );
tran (\sa_snapshot[9][23] , \sa_snapshot[9].f.lower[23] );
tran (\sa_snapshot[9][22] , \sa_snapshot[9].r.part0[22] );
tran (\sa_snapshot[9][22] , \sa_snapshot[9].f.lower[22] );
tran (\sa_snapshot[9][21] , \sa_snapshot[9].r.part0[21] );
tran (\sa_snapshot[9][21] , \sa_snapshot[9].f.lower[21] );
tran (\sa_snapshot[9][20] , \sa_snapshot[9].r.part0[20] );
tran (\sa_snapshot[9][20] , \sa_snapshot[9].f.lower[20] );
tran (\sa_snapshot[9][19] , \sa_snapshot[9].r.part0[19] );
tran (\sa_snapshot[9][19] , \sa_snapshot[9].f.lower[19] );
tran (\sa_snapshot[9][18] , \sa_snapshot[9].r.part0[18] );
tran (\sa_snapshot[9][18] , \sa_snapshot[9].f.lower[18] );
tran (\sa_snapshot[9][17] , \sa_snapshot[9].r.part0[17] );
tran (\sa_snapshot[9][17] , \sa_snapshot[9].f.lower[17] );
tran (\sa_snapshot[9][16] , \sa_snapshot[9].r.part0[16] );
tran (\sa_snapshot[9][16] , \sa_snapshot[9].f.lower[16] );
tran (\sa_snapshot[9][15] , \sa_snapshot[9].r.part0[15] );
tran (\sa_snapshot[9][15] , \sa_snapshot[9].f.lower[15] );
tran (\sa_snapshot[9][14] , \sa_snapshot[9].r.part0[14] );
tran (\sa_snapshot[9][14] , \sa_snapshot[9].f.lower[14] );
tran (\sa_snapshot[9][13] , \sa_snapshot[9].r.part0[13] );
tran (\sa_snapshot[9][13] , \sa_snapshot[9].f.lower[13] );
tran (\sa_snapshot[9][12] , \sa_snapshot[9].r.part0[12] );
tran (\sa_snapshot[9][12] , \sa_snapshot[9].f.lower[12] );
tran (\sa_snapshot[9][11] , \sa_snapshot[9].r.part0[11] );
tran (\sa_snapshot[9][11] , \sa_snapshot[9].f.lower[11] );
tran (\sa_snapshot[9][10] , \sa_snapshot[9].r.part0[10] );
tran (\sa_snapshot[9][10] , \sa_snapshot[9].f.lower[10] );
tran (\sa_snapshot[9][9] , \sa_snapshot[9].r.part0[9] );
tran (\sa_snapshot[9][9] , \sa_snapshot[9].f.lower[9] );
tran (\sa_snapshot[9][8] , \sa_snapshot[9].r.part0[8] );
tran (\sa_snapshot[9][8] , \sa_snapshot[9].f.lower[8] );
tran (\sa_snapshot[9][7] , \sa_snapshot[9].r.part0[7] );
tran (\sa_snapshot[9][7] , \sa_snapshot[9].f.lower[7] );
tran (\sa_snapshot[9][6] , \sa_snapshot[9].r.part0[6] );
tran (\sa_snapshot[9][6] , \sa_snapshot[9].f.lower[6] );
tran (\sa_snapshot[9][5] , \sa_snapshot[9].r.part0[5] );
tran (\sa_snapshot[9][5] , \sa_snapshot[9].f.lower[5] );
tran (\sa_snapshot[9][4] , \sa_snapshot[9].r.part0[4] );
tran (\sa_snapshot[9][4] , \sa_snapshot[9].f.lower[4] );
tran (\sa_snapshot[9][3] , \sa_snapshot[9].r.part0[3] );
tran (\sa_snapshot[9][3] , \sa_snapshot[9].f.lower[3] );
tran (\sa_snapshot[9][2] , \sa_snapshot[9].r.part0[2] );
tran (\sa_snapshot[9][2] , \sa_snapshot[9].f.lower[2] );
tran (\sa_snapshot[9][1] , \sa_snapshot[9].r.part0[1] );
tran (\sa_snapshot[9][1] , \sa_snapshot[9].f.lower[1] );
tran (\sa_snapshot[9][0] , \sa_snapshot[9].r.part0[0] );
tran (\sa_snapshot[9][0] , \sa_snapshot[9].f.lower[0] );
tran (\sa_snapshot[8][63] , \sa_snapshot[8].r.part1[31] );
tran (\sa_snapshot[8][63] , \sa_snapshot[8].f.unused[13] );
tran (\sa_snapshot[8][62] , \sa_snapshot[8].r.part1[30] );
tran (\sa_snapshot[8][62] , \sa_snapshot[8].f.unused[12] );
tran (\sa_snapshot[8][61] , \sa_snapshot[8].r.part1[29] );
tran (\sa_snapshot[8][61] , \sa_snapshot[8].f.unused[11] );
tran (\sa_snapshot[8][60] , \sa_snapshot[8].r.part1[28] );
tran (\sa_snapshot[8][60] , \sa_snapshot[8].f.unused[10] );
tran (\sa_snapshot[8][59] , \sa_snapshot[8].r.part1[27] );
tran (\sa_snapshot[8][59] , \sa_snapshot[8].f.unused[9] );
tran (\sa_snapshot[8][58] , \sa_snapshot[8].r.part1[26] );
tran (\sa_snapshot[8][58] , \sa_snapshot[8].f.unused[8] );
tran (\sa_snapshot[8][57] , \sa_snapshot[8].r.part1[25] );
tran (\sa_snapshot[8][57] , \sa_snapshot[8].f.unused[7] );
tran (\sa_snapshot[8][56] , \sa_snapshot[8].r.part1[24] );
tran (\sa_snapshot[8][56] , \sa_snapshot[8].f.unused[6] );
tran (\sa_snapshot[8][55] , \sa_snapshot[8].r.part1[23] );
tran (\sa_snapshot[8][55] , \sa_snapshot[8].f.unused[5] );
tran (\sa_snapshot[8][54] , \sa_snapshot[8].r.part1[22] );
tran (\sa_snapshot[8][54] , \sa_snapshot[8].f.unused[4] );
tran (\sa_snapshot[8][53] , \sa_snapshot[8].r.part1[21] );
tran (\sa_snapshot[8][53] , \sa_snapshot[8].f.unused[3] );
tran (\sa_snapshot[8][52] , \sa_snapshot[8].r.part1[20] );
tran (\sa_snapshot[8][52] , \sa_snapshot[8].f.unused[2] );
tran (\sa_snapshot[8][51] , \sa_snapshot[8].r.part1[19] );
tran (\sa_snapshot[8][51] , \sa_snapshot[8].f.unused[1] );
tran (\sa_snapshot[8][50] , \sa_snapshot[8].r.part1[18] );
tran (\sa_snapshot[8][50] , \sa_snapshot[8].f.unused[0] );
tran (\sa_snapshot[8][49] , \sa_snapshot[8].r.part1[17] );
tran (\sa_snapshot[8][49] , \sa_snapshot[8].f.upper[17] );
tran (\sa_snapshot[8][48] , \sa_snapshot[8].r.part1[16] );
tran (\sa_snapshot[8][48] , \sa_snapshot[8].f.upper[16] );
tran (\sa_snapshot[8][47] , \sa_snapshot[8].r.part1[15] );
tran (\sa_snapshot[8][47] , \sa_snapshot[8].f.upper[15] );
tran (\sa_snapshot[8][46] , \sa_snapshot[8].r.part1[14] );
tran (\sa_snapshot[8][46] , \sa_snapshot[8].f.upper[14] );
tran (\sa_snapshot[8][45] , \sa_snapshot[8].r.part1[13] );
tran (\sa_snapshot[8][45] , \sa_snapshot[8].f.upper[13] );
tran (\sa_snapshot[8][44] , \sa_snapshot[8].r.part1[12] );
tran (\sa_snapshot[8][44] , \sa_snapshot[8].f.upper[12] );
tran (\sa_snapshot[8][43] , \sa_snapshot[8].r.part1[11] );
tran (\sa_snapshot[8][43] , \sa_snapshot[8].f.upper[11] );
tran (\sa_snapshot[8][42] , \sa_snapshot[8].r.part1[10] );
tran (\sa_snapshot[8][42] , \sa_snapshot[8].f.upper[10] );
tran (\sa_snapshot[8][41] , \sa_snapshot[8].r.part1[9] );
tran (\sa_snapshot[8][41] , \sa_snapshot[8].f.upper[9] );
tran (\sa_snapshot[8][40] , \sa_snapshot[8].r.part1[8] );
tran (\sa_snapshot[8][40] , \sa_snapshot[8].f.upper[8] );
tran (\sa_snapshot[8][39] , \sa_snapshot[8].r.part1[7] );
tran (\sa_snapshot[8][39] , \sa_snapshot[8].f.upper[7] );
tran (\sa_snapshot[8][38] , \sa_snapshot[8].r.part1[6] );
tran (\sa_snapshot[8][38] , \sa_snapshot[8].f.upper[6] );
tran (\sa_snapshot[8][37] , \sa_snapshot[8].r.part1[5] );
tran (\sa_snapshot[8][37] , \sa_snapshot[8].f.upper[5] );
tran (\sa_snapshot[8][36] , \sa_snapshot[8].r.part1[4] );
tran (\sa_snapshot[8][36] , \sa_snapshot[8].f.upper[4] );
tran (\sa_snapshot[8][35] , \sa_snapshot[8].r.part1[3] );
tran (\sa_snapshot[8][35] , \sa_snapshot[8].f.upper[3] );
tran (\sa_snapshot[8][34] , \sa_snapshot[8].r.part1[2] );
tran (\sa_snapshot[8][34] , \sa_snapshot[8].f.upper[2] );
tran (\sa_snapshot[8][33] , \sa_snapshot[8].r.part1[1] );
tran (\sa_snapshot[8][33] , \sa_snapshot[8].f.upper[1] );
tran (\sa_snapshot[8][32] , \sa_snapshot[8].r.part1[0] );
tran (\sa_snapshot[8][32] , \sa_snapshot[8].f.upper[0] );
tran (\sa_snapshot[8][31] , \sa_snapshot[8].r.part0[31] );
tran (\sa_snapshot[8][31] , \sa_snapshot[8].f.lower[31] );
tran (\sa_snapshot[8][30] , \sa_snapshot[8].r.part0[30] );
tran (\sa_snapshot[8][30] , \sa_snapshot[8].f.lower[30] );
tran (\sa_snapshot[8][29] , \sa_snapshot[8].r.part0[29] );
tran (\sa_snapshot[8][29] , \sa_snapshot[8].f.lower[29] );
tran (\sa_snapshot[8][28] , \sa_snapshot[8].r.part0[28] );
tran (\sa_snapshot[8][28] , \sa_snapshot[8].f.lower[28] );
tran (\sa_snapshot[8][27] , \sa_snapshot[8].r.part0[27] );
tran (\sa_snapshot[8][27] , \sa_snapshot[8].f.lower[27] );
tran (\sa_snapshot[8][26] , \sa_snapshot[8].r.part0[26] );
tran (\sa_snapshot[8][26] , \sa_snapshot[8].f.lower[26] );
tran (\sa_snapshot[8][25] , \sa_snapshot[8].r.part0[25] );
tran (\sa_snapshot[8][25] , \sa_snapshot[8].f.lower[25] );
tran (\sa_snapshot[8][24] , \sa_snapshot[8].r.part0[24] );
tran (\sa_snapshot[8][24] , \sa_snapshot[8].f.lower[24] );
tran (\sa_snapshot[8][23] , \sa_snapshot[8].r.part0[23] );
tran (\sa_snapshot[8][23] , \sa_snapshot[8].f.lower[23] );
tran (\sa_snapshot[8][22] , \sa_snapshot[8].r.part0[22] );
tran (\sa_snapshot[8][22] , \sa_snapshot[8].f.lower[22] );
tran (\sa_snapshot[8][21] , \sa_snapshot[8].r.part0[21] );
tran (\sa_snapshot[8][21] , \sa_snapshot[8].f.lower[21] );
tran (\sa_snapshot[8][20] , \sa_snapshot[8].r.part0[20] );
tran (\sa_snapshot[8][20] , \sa_snapshot[8].f.lower[20] );
tran (\sa_snapshot[8][19] , \sa_snapshot[8].r.part0[19] );
tran (\sa_snapshot[8][19] , \sa_snapshot[8].f.lower[19] );
tran (\sa_snapshot[8][18] , \sa_snapshot[8].r.part0[18] );
tran (\sa_snapshot[8][18] , \sa_snapshot[8].f.lower[18] );
tran (\sa_snapshot[8][17] , \sa_snapshot[8].r.part0[17] );
tran (\sa_snapshot[8][17] , \sa_snapshot[8].f.lower[17] );
tran (\sa_snapshot[8][16] , \sa_snapshot[8].r.part0[16] );
tran (\sa_snapshot[8][16] , \sa_snapshot[8].f.lower[16] );
tran (\sa_snapshot[8][15] , \sa_snapshot[8].r.part0[15] );
tran (\sa_snapshot[8][15] , \sa_snapshot[8].f.lower[15] );
tran (\sa_snapshot[8][14] , \sa_snapshot[8].r.part0[14] );
tran (\sa_snapshot[8][14] , \sa_snapshot[8].f.lower[14] );
tran (\sa_snapshot[8][13] , \sa_snapshot[8].r.part0[13] );
tran (\sa_snapshot[8][13] , \sa_snapshot[8].f.lower[13] );
tran (\sa_snapshot[8][12] , \sa_snapshot[8].r.part0[12] );
tran (\sa_snapshot[8][12] , \sa_snapshot[8].f.lower[12] );
tran (\sa_snapshot[8][11] , \sa_snapshot[8].r.part0[11] );
tran (\sa_snapshot[8][11] , \sa_snapshot[8].f.lower[11] );
tran (\sa_snapshot[8][10] , \sa_snapshot[8].r.part0[10] );
tran (\sa_snapshot[8][10] , \sa_snapshot[8].f.lower[10] );
tran (\sa_snapshot[8][9] , \sa_snapshot[8].r.part0[9] );
tran (\sa_snapshot[8][9] , \sa_snapshot[8].f.lower[9] );
tran (\sa_snapshot[8][8] , \sa_snapshot[8].r.part0[8] );
tran (\sa_snapshot[8][8] , \sa_snapshot[8].f.lower[8] );
tran (\sa_snapshot[8][7] , \sa_snapshot[8].r.part0[7] );
tran (\sa_snapshot[8][7] , \sa_snapshot[8].f.lower[7] );
tran (\sa_snapshot[8][6] , \sa_snapshot[8].r.part0[6] );
tran (\sa_snapshot[8][6] , \sa_snapshot[8].f.lower[6] );
tran (\sa_snapshot[8][5] , \sa_snapshot[8].r.part0[5] );
tran (\sa_snapshot[8][5] , \sa_snapshot[8].f.lower[5] );
tran (\sa_snapshot[8][4] , \sa_snapshot[8].r.part0[4] );
tran (\sa_snapshot[8][4] , \sa_snapshot[8].f.lower[4] );
tran (\sa_snapshot[8][3] , \sa_snapshot[8].r.part0[3] );
tran (\sa_snapshot[8][3] , \sa_snapshot[8].f.lower[3] );
tran (\sa_snapshot[8][2] , \sa_snapshot[8].r.part0[2] );
tran (\sa_snapshot[8][2] , \sa_snapshot[8].f.lower[2] );
tran (\sa_snapshot[8][1] , \sa_snapshot[8].r.part0[1] );
tran (\sa_snapshot[8][1] , \sa_snapshot[8].f.lower[1] );
tran (\sa_snapshot[8][0] , \sa_snapshot[8].r.part0[0] );
tran (\sa_snapshot[8][0] , \sa_snapshot[8].f.lower[0] );
tran (\sa_snapshot[7][63] , \sa_snapshot[7].r.part1[31] );
tran (\sa_snapshot[7][63] , \sa_snapshot[7].f.unused[13] );
tran (\sa_snapshot[7][62] , \sa_snapshot[7].r.part1[30] );
tran (\sa_snapshot[7][62] , \sa_snapshot[7].f.unused[12] );
tran (\sa_snapshot[7][61] , \sa_snapshot[7].r.part1[29] );
tran (\sa_snapshot[7][61] , \sa_snapshot[7].f.unused[11] );
tran (\sa_snapshot[7][60] , \sa_snapshot[7].r.part1[28] );
tran (\sa_snapshot[7][60] , \sa_snapshot[7].f.unused[10] );
tran (\sa_snapshot[7][59] , \sa_snapshot[7].r.part1[27] );
tran (\sa_snapshot[7][59] , \sa_snapshot[7].f.unused[9] );
tran (\sa_snapshot[7][58] , \sa_snapshot[7].r.part1[26] );
tran (\sa_snapshot[7][58] , \sa_snapshot[7].f.unused[8] );
tran (\sa_snapshot[7][57] , \sa_snapshot[7].r.part1[25] );
tran (\sa_snapshot[7][57] , \sa_snapshot[7].f.unused[7] );
tran (\sa_snapshot[7][56] , \sa_snapshot[7].r.part1[24] );
tran (\sa_snapshot[7][56] , \sa_snapshot[7].f.unused[6] );
tran (\sa_snapshot[7][55] , \sa_snapshot[7].r.part1[23] );
tran (\sa_snapshot[7][55] , \sa_snapshot[7].f.unused[5] );
tran (\sa_snapshot[7][54] , \sa_snapshot[7].r.part1[22] );
tran (\sa_snapshot[7][54] , \sa_snapshot[7].f.unused[4] );
tran (\sa_snapshot[7][53] , \sa_snapshot[7].r.part1[21] );
tran (\sa_snapshot[7][53] , \sa_snapshot[7].f.unused[3] );
tran (\sa_snapshot[7][52] , \sa_snapshot[7].r.part1[20] );
tran (\sa_snapshot[7][52] , \sa_snapshot[7].f.unused[2] );
tran (\sa_snapshot[7][51] , \sa_snapshot[7].r.part1[19] );
tran (\sa_snapshot[7][51] , \sa_snapshot[7].f.unused[1] );
tran (\sa_snapshot[7][50] , \sa_snapshot[7].r.part1[18] );
tran (\sa_snapshot[7][50] , \sa_snapshot[7].f.unused[0] );
tran (\sa_snapshot[7][49] , \sa_snapshot[7].r.part1[17] );
tran (\sa_snapshot[7][49] , \sa_snapshot[7].f.upper[17] );
tran (\sa_snapshot[7][48] , \sa_snapshot[7].r.part1[16] );
tran (\sa_snapshot[7][48] , \sa_snapshot[7].f.upper[16] );
tran (\sa_snapshot[7][47] , \sa_snapshot[7].r.part1[15] );
tran (\sa_snapshot[7][47] , \sa_snapshot[7].f.upper[15] );
tran (\sa_snapshot[7][46] , \sa_snapshot[7].r.part1[14] );
tran (\sa_snapshot[7][46] , \sa_snapshot[7].f.upper[14] );
tran (\sa_snapshot[7][45] , \sa_snapshot[7].r.part1[13] );
tran (\sa_snapshot[7][45] , \sa_snapshot[7].f.upper[13] );
tran (\sa_snapshot[7][44] , \sa_snapshot[7].r.part1[12] );
tran (\sa_snapshot[7][44] , \sa_snapshot[7].f.upper[12] );
tran (\sa_snapshot[7][43] , \sa_snapshot[7].r.part1[11] );
tran (\sa_snapshot[7][43] , \sa_snapshot[7].f.upper[11] );
tran (\sa_snapshot[7][42] , \sa_snapshot[7].r.part1[10] );
tran (\sa_snapshot[7][42] , \sa_snapshot[7].f.upper[10] );
tran (\sa_snapshot[7][41] , \sa_snapshot[7].r.part1[9] );
tran (\sa_snapshot[7][41] , \sa_snapshot[7].f.upper[9] );
tran (\sa_snapshot[7][40] , \sa_snapshot[7].r.part1[8] );
tran (\sa_snapshot[7][40] , \sa_snapshot[7].f.upper[8] );
tran (\sa_snapshot[7][39] , \sa_snapshot[7].r.part1[7] );
tran (\sa_snapshot[7][39] , \sa_snapshot[7].f.upper[7] );
tran (\sa_snapshot[7][38] , \sa_snapshot[7].r.part1[6] );
tran (\sa_snapshot[7][38] , \sa_snapshot[7].f.upper[6] );
tran (\sa_snapshot[7][37] , \sa_snapshot[7].r.part1[5] );
tran (\sa_snapshot[7][37] , \sa_snapshot[7].f.upper[5] );
tran (\sa_snapshot[7][36] , \sa_snapshot[7].r.part1[4] );
tran (\sa_snapshot[7][36] , \sa_snapshot[7].f.upper[4] );
tran (\sa_snapshot[7][35] , \sa_snapshot[7].r.part1[3] );
tran (\sa_snapshot[7][35] , \sa_snapshot[7].f.upper[3] );
tran (\sa_snapshot[7][34] , \sa_snapshot[7].r.part1[2] );
tran (\sa_snapshot[7][34] , \sa_snapshot[7].f.upper[2] );
tran (\sa_snapshot[7][33] , \sa_snapshot[7].r.part1[1] );
tran (\sa_snapshot[7][33] , \sa_snapshot[7].f.upper[1] );
tran (\sa_snapshot[7][32] , \sa_snapshot[7].r.part1[0] );
tran (\sa_snapshot[7][32] , \sa_snapshot[7].f.upper[0] );
tran (\sa_snapshot[7][31] , \sa_snapshot[7].r.part0[31] );
tran (\sa_snapshot[7][31] , \sa_snapshot[7].f.lower[31] );
tran (\sa_snapshot[7][30] , \sa_snapshot[7].r.part0[30] );
tran (\sa_snapshot[7][30] , \sa_snapshot[7].f.lower[30] );
tran (\sa_snapshot[7][29] , \sa_snapshot[7].r.part0[29] );
tran (\sa_snapshot[7][29] , \sa_snapshot[7].f.lower[29] );
tran (\sa_snapshot[7][28] , \sa_snapshot[7].r.part0[28] );
tran (\sa_snapshot[7][28] , \sa_snapshot[7].f.lower[28] );
tran (\sa_snapshot[7][27] , \sa_snapshot[7].r.part0[27] );
tran (\sa_snapshot[7][27] , \sa_snapshot[7].f.lower[27] );
tran (\sa_snapshot[7][26] , \sa_snapshot[7].r.part0[26] );
tran (\sa_snapshot[7][26] , \sa_snapshot[7].f.lower[26] );
tran (\sa_snapshot[7][25] , \sa_snapshot[7].r.part0[25] );
tran (\sa_snapshot[7][25] , \sa_snapshot[7].f.lower[25] );
tran (\sa_snapshot[7][24] , \sa_snapshot[7].r.part0[24] );
tran (\sa_snapshot[7][24] , \sa_snapshot[7].f.lower[24] );
tran (\sa_snapshot[7][23] , \sa_snapshot[7].r.part0[23] );
tran (\sa_snapshot[7][23] , \sa_snapshot[7].f.lower[23] );
tran (\sa_snapshot[7][22] , \sa_snapshot[7].r.part0[22] );
tran (\sa_snapshot[7][22] , \sa_snapshot[7].f.lower[22] );
tran (\sa_snapshot[7][21] , \sa_snapshot[7].r.part0[21] );
tran (\sa_snapshot[7][21] , \sa_snapshot[7].f.lower[21] );
tran (\sa_snapshot[7][20] , \sa_snapshot[7].r.part0[20] );
tran (\sa_snapshot[7][20] , \sa_snapshot[7].f.lower[20] );
tran (\sa_snapshot[7][19] , \sa_snapshot[7].r.part0[19] );
tran (\sa_snapshot[7][19] , \sa_snapshot[7].f.lower[19] );
tran (\sa_snapshot[7][18] , \sa_snapshot[7].r.part0[18] );
tran (\sa_snapshot[7][18] , \sa_snapshot[7].f.lower[18] );
tran (\sa_snapshot[7][17] , \sa_snapshot[7].r.part0[17] );
tran (\sa_snapshot[7][17] , \sa_snapshot[7].f.lower[17] );
tran (\sa_snapshot[7][16] , \sa_snapshot[7].r.part0[16] );
tran (\sa_snapshot[7][16] , \sa_snapshot[7].f.lower[16] );
tran (\sa_snapshot[7][15] , \sa_snapshot[7].r.part0[15] );
tran (\sa_snapshot[7][15] , \sa_snapshot[7].f.lower[15] );
tran (\sa_snapshot[7][14] , \sa_snapshot[7].r.part0[14] );
tran (\sa_snapshot[7][14] , \sa_snapshot[7].f.lower[14] );
tran (\sa_snapshot[7][13] , \sa_snapshot[7].r.part0[13] );
tran (\sa_snapshot[7][13] , \sa_snapshot[7].f.lower[13] );
tran (\sa_snapshot[7][12] , \sa_snapshot[7].r.part0[12] );
tran (\sa_snapshot[7][12] , \sa_snapshot[7].f.lower[12] );
tran (\sa_snapshot[7][11] , \sa_snapshot[7].r.part0[11] );
tran (\sa_snapshot[7][11] , \sa_snapshot[7].f.lower[11] );
tran (\sa_snapshot[7][10] , \sa_snapshot[7].r.part0[10] );
tran (\sa_snapshot[7][10] , \sa_snapshot[7].f.lower[10] );
tran (\sa_snapshot[7][9] , \sa_snapshot[7].r.part0[9] );
tran (\sa_snapshot[7][9] , \sa_snapshot[7].f.lower[9] );
tran (\sa_snapshot[7][8] , \sa_snapshot[7].r.part0[8] );
tran (\sa_snapshot[7][8] , \sa_snapshot[7].f.lower[8] );
tran (\sa_snapshot[7][7] , \sa_snapshot[7].r.part0[7] );
tran (\sa_snapshot[7][7] , \sa_snapshot[7].f.lower[7] );
tran (\sa_snapshot[7][6] , \sa_snapshot[7].r.part0[6] );
tran (\sa_snapshot[7][6] , \sa_snapshot[7].f.lower[6] );
tran (\sa_snapshot[7][5] , \sa_snapshot[7].r.part0[5] );
tran (\sa_snapshot[7][5] , \sa_snapshot[7].f.lower[5] );
tran (\sa_snapshot[7][4] , \sa_snapshot[7].r.part0[4] );
tran (\sa_snapshot[7][4] , \sa_snapshot[7].f.lower[4] );
tran (\sa_snapshot[7][3] , \sa_snapshot[7].r.part0[3] );
tran (\sa_snapshot[7][3] , \sa_snapshot[7].f.lower[3] );
tran (\sa_snapshot[7][2] , \sa_snapshot[7].r.part0[2] );
tran (\sa_snapshot[7][2] , \sa_snapshot[7].f.lower[2] );
tran (\sa_snapshot[7][1] , \sa_snapshot[7].r.part0[1] );
tran (\sa_snapshot[7][1] , \sa_snapshot[7].f.lower[1] );
tran (\sa_snapshot[7][0] , \sa_snapshot[7].r.part0[0] );
tran (\sa_snapshot[7][0] , \sa_snapshot[7].f.lower[0] );
tran (\sa_snapshot[6][63] , \sa_snapshot[6].r.part1[31] );
tran (\sa_snapshot[6][63] , \sa_snapshot[6].f.unused[13] );
tran (\sa_snapshot[6][62] , \sa_snapshot[6].r.part1[30] );
tran (\sa_snapshot[6][62] , \sa_snapshot[6].f.unused[12] );
tran (\sa_snapshot[6][61] , \sa_snapshot[6].r.part1[29] );
tran (\sa_snapshot[6][61] , \sa_snapshot[6].f.unused[11] );
tran (\sa_snapshot[6][60] , \sa_snapshot[6].r.part1[28] );
tran (\sa_snapshot[6][60] , \sa_snapshot[6].f.unused[10] );
tran (\sa_snapshot[6][59] , \sa_snapshot[6].r.part1[27] );
tran (\sa_snapshot[6][59] , \sa_snapshot[6].f.unused[9] );
tran (\sa_snapshot[6][58] , \sa_snapshot[6].r.part1[26] );
tran (\sa_snapshot[6][58] , \sa_snapshot[6].f.unused[8] );
tran (\sa_snapshot[6][57] , \sa_snapshot[6].r.part1[25] );
tran (\sa_snapshot[6][57] , \sa_snapshot[6].f.unused[7] );
tran (\sa_snapshot[6][56] , \sa_snapshot[6].r.part1[24] );
tran (\sa_snapshot[6][56] , \sa_snapshot[6].f.unused[6] );
tran (\sa_snapshot[6][55] , \sa_snapshot[6].r.part1[23] );
tran (\sa_snapshot[6][55] , \sa_snapshot[6].f.unused[5] );
tran (\sa_snapshot[6][54] , \sa_snapshot[6].r.part1[22] );
tran (\sa_snapshot[6][54] , \sa_snapshot[6].f.unused[4] );
tran (\sa_snapshot[6][53] , \sa_snapshot[6].r.part1[21] );
tran (\sa_snapshot[6][53] , \sa_snapshot[6].f.unused[3] );
tran (\sa_snapshot[6][52] , \sa_snapshot[6].r.part1[20] );
tran (\sa_snapshot[6][52] , \sa_snapshot[6].f.unused[2] );
tran (\sa_snapshot[6][51] , \sa_snapshot[6].r.part1[19] );
tran (\sa_snapshot[6][51] , \sa_snapshot[6].f.unused[1] );
tran (\sa_snapshot[6][50] , \sa_snapshot[6].r.part1[18] );
tran (\sa_snapshot[6][50] , \sa_snapshot[6].f.unused[0] );
tran (\sa_snapshot[6][49] , \sa_snapshot[6].r.part1[17] );
tran (\sa_snapshot[6][49] , \sa_snapshot[6].f.upper[17] );
tran (\sa_snapshot[6][48] , \sa_snapshot[6].r.part1[16] );
tran (\sa_snapshot[6][48] , \sa_snapshot[6].f.upper[16] );
tran (\sa_snapshot[6][47] , \sa_snapshot[6].r.part1[15] );
tran (\sa_snapshot[6][47] , \sa_snapshot[6].f.upper[15] );
tran (\sa_snapshot[6][46] , \sa_snapshot[6].r.part1[14] );
tran (\sa_snapshot[6][46] , \sa_snapshot[6].f.upper[14] );
tran (\sa_snapshot[6][45] , \sa_snapshot[6].r.part1[13] );
tran (\sa_snapshot[6][45] , \sa_snapshot[6].f.upper[13] );
tran (\sa_snapshot[6][44] , \sa_snapshot[6].r.part1[12] );
tran (\sa_snapshot[6][44] , \sa_snapshot[6].f.upper[12] );
tran (\sa_snapshot[6][43] , \sa_snapshot[6].r.part1[11] );
tran (\sa_snapshot[6][43] , \sa_snapshot[6].f.upper[11] );
tran (\sa_snapshot[6][42] , \sa_snapshot[6].r.part1[10] );
tran (\sa_snapshot[6][42] , \sa_snapshot[6].f.upper[10] );
tran (\sa_snapshot[6][41] , \sa_snapshot[6].r.part1[9] );
tran (\sa_snapshot[6][41] , \sa_snapshot[6].f.upper[9] );
tran (\sa_snapshot[6][40] , \sa_snapshot[6].r.part1[8] );
tran (\sa_snapshot[6][40] , \sa_snapshot[6].f.upper[8] );
tran (\sa_snapshot[6][39] , \sa_snapshot[6].r.part1[7] );
tran (\sa_snapshot[6][39] , \sa_snapshot[6].f.upper[7] );
tran (\sa_snapshot[6][38] , \sa_snapshot[6].r.part1[6] );
tran (\sa_snapshot[6][38] , \sa_snapshot[6].f.upper[6] );
tran (\sa_snapshot[6][37] , \sa_snapshot[6].r.part1[5] );
tran (\sa_snapshot[6][37] , \sa_snapshot[6].f.upper[5] );
tran (\sa_snapshot[6][36] , \sa_snapshot[6].r.part1[4] );
tran (\sa_snapshot[6][36] , \sa_snapshot[6].f.upper[4] );
tran (\sa_snapshot[6][35] , \sa_snapshot[6].r.part1[3] );
tran (\sa_snapshot[6][35] , \sa_snapshot[6].f.upper[3] );
tran (\sa_snapshot[6][34] , \sa_snapshot[6].r.part1[2] );
tran (\sa_snapshot[6][34] , \sa_snapshot[6].f.upper[2] );
tran (\sa_snapshot[6][33] , \sa_snapshot[6].r.part1[1] );
tran (\sa_snapshot[6][33] , \sa_snapshot[6].f.upper[1] );
tran (\sa_snapshot[6][32] , \sa_snapshot[6].r.part1[0] );
tran (\sa_snapshot[6][32] , \sa_snapshot[6].f.upper[0] );
tran (\sa_snapshot[6][31] , \sa_snapshot[6].r.part0[31] );
tran (\sa_snapshot[6][31] , \sa_snapshot[6].f.lower[31] );
tran (\sa_snapshot[6][30] , \sa_snapshot[6].r.part0[30] );
tran (\sa_snapshot[6][30] , \sa_snapshot[6].f.lower[30] );
tran (\sa_snapshot[6][29] , \sa_snapshot[6].r.part0[29] );
tran (\sa_snapshot[6][29] , \sa_snapshot[6].f.lower[29] );
tran (\sa_snapshot[6][28] , \sa_snapshot[6].r.part0[28] );
tran (\sa_snapshot[6][28] , \sa_snapshot[6].f.lower[28] );
tran (\sa_snapshot[6][27] , \sa_snapshot[6].r.part0[27] );
tran (\sa_snapshot[6][27] , \sa_snapshot[6].f.lower[27] );
tran (\sa_snapshot[6][26] , \sa_snapshot[6].r.part0[26] );
tran (\sa_snapshot[6][26] , \sa_snapshot[6].f.lower[26] );
tran (\sa_snapshot[6][25] , \sa_snapshot[6].r.part0[25] );
tran (\sa_snapshot[6][25] , \sa_snapshot[6].f.lower[25] );
tran (\sa_snapshot[6][24] , \sa_snapshot[6].r.part0[24] );
tran (\sa_snapshot[6][24] , \sa_snapshot[6].f.lower[24] );
tran (\sa_snapshot[6][23] , \sa_snapshot[6].r.part0[23] );
tran (\sa_snapshot[6][23] , \sa_snapshot[6].f.lower[23] );
tran (\sa_snapshot[6][22] , \sa_snapshot[6].r.part0[22] );
tran (\sa_snapshot[6][22] , \sa_snapshot[6].f.lower[22] );
tran (\sa_snapshot[6][21] , \sa_snapshot[6].r.part0[21] );
tran (\sa_snapshot[6][21] , \sa_snapshot[6].f.lower[21] );
tran (\sa_snapshot[6][20] , \sa_snapshot[6].r.part0[20] );
tran (\sa_snapshot[6][20] , \sa_snapshot[6].f.lower[20] );
tran (\sa_snapshot[6][19] , \sa_snapshot[6].r.part0[19] );
tran (\sa_snapshot[6][19] , \sa_snapshot[6].f.lower[19] );
tran (\sa_snapshot[6][18] , \sa_snapshot[6].r.part0[18] );
tran (\sa_snapshot[6][18] , \sa_snapshot[6].f.lower[18] );
tran (\sa_snapshot[6][17] , \sa_snapshot[6].r.part0[17] );
tran (\sa_snapshot[6][17] , \sa_snapshot[6].f.lower[17] );
tran (\sa_snapshot[6][16] , \sa_snapshot[6].r.part0[16] );
tran (\sa_snapshot[6][16] , \sa_snapshot[6].f.lower[16] );
tran (\sa_snapshot[6][15] , \sa_snapshot[6].r.part0[15] );
tran (\sa_snapshot[6][15] , \sa_snapshot[6].f.lower[15] );
tran (\sa_snapshot[6][14] , \sa_snapshot[6].r.part0[14] );
tran (\sa_snapshot[6][14] , \sa_snapshot[6].f.lower[14] );
tran (\sa_snapshot[6][13] , \sa_snapshot[6].r.part0[13] );
tran (\sa_snapshot[6][13] , \sa_snapshot[6].f.lower[13] );
tran (\sa_snapshot[6][12] , \sa_snapshot[6].r.part0[12] );
tran (\sa_snapshot[6][12] , \sa_snapshot[6].f.lower[12] );
tran (\sa_snapshot[6][11] , \sa_snapshot[6].r.part0[11] );
tran (\sa_snapshot[6][11] , \sa_snapshot[6].f.lower[11] );
tran (\sa_snapshot[6][10] , \sa_snapshot[6].r.part0[10] );
tran (\sa_snapshot[6][10] , \sa_snapshot[6].f.lower[10] );
tran (\sa_snapshot[6][9] , \sa_snapshot[6].r.part0[9] );
tran (\sa_snapshot[6][9] , \sa_snapshot[6].f.lower[9] );
tran (\sa_snapshot[6][8] , \sa_snapshot[6].r.part0[8] );
tran (\sa_snapshot[6][8] , \sa_snapshot[6].f.lower[8] );
tran (\sa_snapshot[6][7] , \sa_snapshot[6].r.part0[7] );
tran (\sa_snapshot[6][7] , \sa_snapshot[6].f.lower[7] );
tran (\sa_snapshot[6][6] , \sa_snapshot[6].r.part0[6] );
tran (\sa_snapshot[6][6] , \sa_snapshot[6].f.lower[6] );
tran (\sa_snapshot[6][5] , \sa_snapshot[6].r.part0[5] );
tran (\sa_snapshot[6][5] , \sa_snapshot[6].f.lower[5] );
tran (\sa_snapshot[6][4] , \sa_snapshot[6].r.part0[4] );
tran (\sa_snapshot[6][4] , \sa_snapshot[6].f.lower[4] );
tran (\sa_snapshot[6][3] , \sa_snapshot[6].r.part0[3] );
tran (\sa_snapshot[6][3] , \sa_snapshot[6].f.lower[3] );
tran (\sa_snapshot[6][2] , \sa_snapshot[6].r.part0[2] );
tran (\sa_snapshot[6][2] , \sa_snapshot[6].f.lower[2] );
tran (\sa_snapshot[6][1] , \sa_snapshot[6].r.part0[1] );
tran (\sa_snapshot[6][1] , \sa_snapshot[6].f.lower[1] );
tran (\sa_snapshot[6][0] , \sa_snapshot[6].r.part0[0] );
tran (\sa_snapshot[6][0] , \sa_snapshot[6].f.lower[0] );
tran (\sa_snapshot[5][63] , \sa_snapshot[5].r.part1[31] );
tran (\sa_snapshot[5][63] , \sa_snapshot[5].f.unused[13] );
tran (\sa_snapshot[5][62] , \sa_snapshot[5].r.part1[30] );
tran (\sa_snapshot[5][62] , \sa_snapshot[5].f.unused[12] );
tran (\sa_snapshot[5][61] , \sa_snapshot[5].r.part1[29] );
tran (\sa_snapshot[5][61] , \sa_snapshot[5].f.unused[11] );
tran (\sa_snapshot[5][60] , \sa_snapshot[5].r.part1[28] );
tran (\sa_snapshot[5][60] , \sa_snapshot[5].f.unused[10] );
tran (\sa_snapshot[5][59] , \sa_snapshot[5].r.part1[27] );
tran (\sa_snapshot[5][59] , \sa_snapshot[5].f.unused[9] );
tran (\sa_snapshot[5][58] , \sa_snapshot[5].r.part1[26] );
tran (\sa_snapshot[5][58] , \sa_snapshot[5].f.unused[8] );
tran (\sa_snapshot[5][57] , \sa_snapshot[5].r.part1[25] );
tran (\sa_snapshot[5][57] , \sa_snapshot[5].f.unused[7] );
tran (\sa_snapshot[5][56] , \sa_snapshot[5].r.part1[24] );
tran (\sa_snapshot[5][56] , \sa_snapshot[5].f.unused[6] );
tran (\sa_snapshot[5][55] , \sa_snapshot[5].r.part1[23] );
tran (\sa_snapshot[5][55] , \sa_snapshot[5].f.unused[5] );
tran (\sa_snapshot[5][54] , \sa_snapshot[5].r.part1[22] );
tran (\sa_snapshot[5][54] , \sa_snapshot[5].f.unused[4] );
tran (\sa_snapshot[5][53] , \sa_snapshot[5].r.part1[21] );
tran (\sa_snapshot[5][53] , \sa_snapshot[5].f.unused[3] );
tran (\sa_snapshot[5][52] , \sa_snapshot[5].r.part1[20] );
tran (\sa_snapshot[5][52] , \sa_snapshot[5].f.unused[2] );
tran (\sa_snapshot[5][51] , \sa_snapshot[5].r.part1[19] );
tran (\sa_snapshot[5][51] , \sa_snapshot[5].f.unused[1] );
tran (\sa_snapshot[5][50] , \sa_snapshot[5].r.part1[18] );
tran (\sa_snapshot[5][50] , \sa_snapshot[5].f.unused[0] );
tran (\sa_snapshot[5][49] , \sa_snapshot[5].r.part1[17] );
tran (\sa_snapshot[5][49] , \sa_snapshot[5].f.upper[17] );
tran (\sa_snapshot[5][48] , \sa_snapshot[5].r.part1[16] );
tran (\sa_snapshot[5][48] , \sa_snapshot[5].f.upper[16] );
tran (\sa_snapshot[5][47] , \sa_snapshot[5].r.part1[15] );
tran (\sa_snapshot[5][47] , \sa_snapshot[5].f.upper[15] );
tran (\sa_snapshot[5][46] , \sa_snapshot[5].r.part1[14] );
tran (\sa_snapshot[5][46] , \sa_snapshot[5].f.upper[14] );
tran (\sa_snapshot[5][45] , \sa_snapshot[5].r.part1[13] );
tran (\sa_snapshot[5][45] , \sa_snapshot[5].f.upper[13] );
tran (\sa_snapshot[5][44] , \sa_snapshot[5].r.part1[12] );
tran (\sa_snapshot[5][44] , \sa_snapshot[5].f.upper[12] );
tran (\sa_snapshot[5][43] , \sa_snapshot[5].r.part1[11] );
tran (\sa_snapshot[5][43] , \sa_snapshot[5].f.upper[11] );
tran (\sa_snapshot[5][42] , \sa_snapshot[5].r.part1[10] );
tran (\sa_snapshot[5][42] , \sa_snapshot[5].f.upper[10] );
tran (\sa_snapshot[5][41] , \sa_snapshot[5].r.part1[9] );
tran (\sa_snapshot[5][41] , \sa_snapshot[5].f.upper[9] );
tran (\sa_snapshot[5][40] , \sa_snapshot[5].r.part1[8] );
tran (\sa_snapshot[5][40] , \sa_snapshot[5].f.upper[8] );
tran (\sa_snapshot[5][39] , \sa_snapshot[5].r.part1[7] );
tran (\sa_snapshot[5][39] , \sa_snapshot[5].f.upper[7] );
tran (\sa_snapshot[5][38] , \sa_snapshot[5].r.part1[6] );
tran (\sa_snapshot[5][38] , \sa_snapshot[5].f.upper[6] );
tran (\sa_snapshot[5][37] , \sa_snapshot[5].r.part1[5] );
tran (\sa_snapshot[5][37] , \sa_snapshot[5].f.upper[5] );
tran (\sa_snapshot[5][36] , \sa_snapshot[5].r.part1[4] );
tran (\sa_snapshot[5][36] , \sa_snapshot[5].f.upper[4] );
tran (\sa_snapshot[5][35] , \sa_snapshot[5].r.part1[3] );
tran (\sa_snapshot[5][35] , \sa_snapshot[5].f.upper[3] );
tran (\sa_snapshot[5][34] , \sa_snapshot[5].r.part1[2] );
tran (\sa_snapshot[5][34] , \sa_snapshot[5].f.upper[2] );
tran (\sa_snapshot[5][33] , \sa_snapshot[5].r.part1[1] );
tran (\sa_snapshot[5][33] , \sa_snapshot[5].f.upper[1] );
tran (\sa_snapshot[5][32] , \sa_snapshot[5].r.part1[0] );
tran (\sa_snapshot[5][32] , \sa_snapshot[5].f.upper[0] );
tran (\sa_snapshot[5][31] , \sa_snapshot[5].r.part0[31] );
tran (\sa_snapshot[5][31] , \sa_snapshot[5].f.lower[31] );
tran (\sa_snapshot[5][30] , \sa_snapshot[5].r.part0[30] );
tran (\sa_snapshot[5][30] , \sa_snapshot[5].f.lower[30] );
tran (\sa_snapshot[5][29] , \sa_snapshot[5].r.part0[29] );
tran (\sa_snapshot[5][29] , \sa_snapshot[5].f.lower[29] );
tran (\sa_snapshot[5][28] , \sa_snapshot[5].r.part0[28] );
tran (\sa_snapshot[5][28] , \sa_snapshot[5].f.lower[28] );
tran (\sa_snapshot[5][27] , \sa_snapshot[5].r.part0[27] );
tran (\sa_snapshot[5][27] , \sa_snapshot[5].f.lower[27] );
tran (\sa_snapshot[5][26] , \sa_snapshot[5].r.part0[26] );
tran (\sa_snapshot[5][26] , \sa_snapshot[5].f.lower[26] );
tran (\sa_snapshot[5][25] , \sa_snapshot[5].r.part0[25] );
tran (\sa_snapshot[5][25] , \sa_snapshot[5].f.lower[25] );
tran (\sa_snapshot[5][24] , \sa_snapshot[5].r.part0[24] );
tran (\sa_snapshot[5][24] , \sa_snapshot[5].f.lower[24] );
tran (\sa_snapshot[5][23] , \sa_snapshot[5].r.part0[23] );
tran (\sa_snapshot[5][23] , \sa_snapshot[5].f.lower[23] );
tran (\sa_snapshot[5][22] , \sa_snapshot[5].r.part0[22] );
tran (\sa_snapshot[5][22] , \sa_snapshot[5].f.lower[22] );
tran (\sa_snapshot[5][21] , \sa_snapshot[5].r.part0[21] );
tran (\sa_snapshot[5][21] , \sa_snapshot[5].f.lower[21] );
tran (\sa_snapshot[5][20] , \sa_snapshot[5].r.part0[20] );
tran (\sa_snapshot[5][20] , \sa_snapshot[5].f.lower[20] );
tran (\sa_snapshot[5][19] , \sa_snapshot[5].r.part0[19] );
tran (\sa_snapshot[5][19] , \sa_snapshot[5].f.lower[19] );
tran (\sa_snapshot[5][18] , \sa_snapshot[5].r.part0[18] );
tran (\sa_snapshot[5][18] , \sa_snapshot[5].f.lower[18] );
tran (\sa_snapshot[5][17] , \sa_snapshot[5].r.part0[17] );
tran (\sa_snapshot[5][17] , \sa_snapshot[5].f.lower[17] );
tran (\sa_snapshot[5][16] , \sa_snapshot[5].r.part0[16] );
tran (\sa_snapshot[5][16] , \sa_snapshot[5].f.lower[16] );
tran (\sa_snapshot[5][15] , \sa_snapshot[5].r.part0[15] );
tran (\sa_snapshot[5][15] , \sa_snapshot[5].f.lower[15] );
tran (\sa_snapshot[5][14] , \sa_snapshot[5].r.part0[14] );
tran (\sa_snapshot[5][14] , \sa_snapshot[5].f.lower[14] );
tran (\sa_snapshot[5][13] , \sa_snapshot[5].r.part0[13] );
tran (\sa_snapshot[5][13] , \sa_snapshot[5].f.lower[13] );
tran (\sa_snapshot[5][12] , \sa_snapshot[5].r.part0[12] );
tran (\sa_snapshot[5][12] , \sa_snapshot[5].f.lower[12] );
tran (\sa_snapshot[5][11] , \sa_snapshot[5].r.part0[11] );
tran (\sa_snapshot[5][11] , \sa_snapshot[5].f.lower[11] );
tran (\sa_snapshot[5][10] , \sa_snapshot[5].r.part0[10] );
tran (\sa_snapshot[5][10] , \sa_snapshot[5].f.lower[10] );
tran (\sa_snapshot[5][9] , \sa_snapshot[5].r.part0[9] );
tran (\sa_snapshot[5][9] , \sa_snapshot[5].f.lower[9] );
tran (\sa_snapshot[5][8] , \sa_snapshot[5].r.part0[8] );
tran (\sa_snapshot[5][8] , \sa_snapshot[5].f.lower[8] );
tran (\sa_snapshot[5][7] , \sa_snapshot[5].r.part0[7] );
tran (\sa_snapshot[5][7] , \sa_snapshot[5].f.lower[7] );
tran (\sa_snapshot[5][6] , \sa_snapshot[5].r.part0[6] );
tran (\sa_snapshot[5][6] , \sa_snapshot[5].f.lower[6] );
tran (\sa_snapshot[5][5] , \sa_snapshot[5].r.part0[5] );
tran (\sa_snapshot[5][5] , \sa_snapshot[5].f.lower[5] );
tran (\sa_snapshot[5][4] , \sa_snapshot[5].r.part0[4] );
tran (\sa_snapshot[5][4] , \sa_snapshot[5].f.lower[4] );
tran (\sa_snapshot[5][3] , \sa_snapshot[5].r.part0[3] );
tran (\sa_snapshot[5][3] , \sa_snapshot[5].f.lower[3] );
tran (\sa_snapshot[5][2] , \sa_snapshot[5].r.part0[2] );
tran (\sa_snapshot[5][2] , \sa_snapshot[5].f.lower[2] );
tran (\sa_snapshot[5][1] , \sa_snapshot[5].r.part0[1] );
tran (\sa_snapshot[5][1] , \sa_snapshot[5].f.lower[1] );
tran (\sa_snapshot[5][0] , \sa_snapshot[5].r.part0[0] );
tran (\sa_snapshot[5][0] , \sa_snapshot[5].f.lower[0] );
tran (\sa_snapshot[4][63] , \sa_snapshot[4].r.part1[31] );
tran (\sa_snapshot[4][63] , \sa_snapshot[4].f.unused[13] );
tran (\sa_snapshot[4][62] , \sa_snapshot[4].r.part1[30] );
tran (\sa_snapshot[4][62] , \sa_snapshot[4].f.unused[12] );
tran (\sa_snapshot[4][61] , \sa_snapshot[4].r.part1[29] );
tran (\sa_snapshot[4][61] , \sa_snapshot[4].f.unused[11] );
tran (\sa_snapshot[4][60] , \sa_snapshot[4].r.part1[28] );
tran (\sa_snapshot[4][60] , \sa_snapshot[4].f.unused[10] );
tran (\sa_snapshot[4][59] , \sa_snapshot[4].r.part1[27] );
tran (\sa_snapshot[4][59] , \sa_snapshot[4].f.unused[9] );
tran (\sa_snapshot[4][58] , \sa_snapshot[4].r.part1[26] );
tran (\sa_snapshot[4][58] , \sa_snapshot[4].f.unused[8] );
tran (\sa_snapshot[4][57] , \sa_snapshot[4].r.part1[25] );
tran (\sa_snapshot[4][57] , \sa_snapshot[4].f.unused[7] );
tran (\sa_snapshot[4][56] , \sa_snapshot[4].r.part1[24] );
tran (\sa_snapshot[4][56] , \sa_snapshot[4].f.unused[6] );
tran (\sa_snapshot[4][55] , \sa_snapshot[4].r.part1[23] );
tran (\sa_snapshot[4][55] , \sa_snapshot[4].f.unused[5] );
tran (\sa_snapshot[4][54] , \sa_snapshot[4].r.part1[22] );
tran (\sa_snapshot[4][54] , \sa_snapshot[4].f.unused[4] );
tran (\sa_snapshot[4][53] , \sa_snapshot[4].r.part1[21] );
tran (\sa_snapshot[4][53] , \sa_snapshot[4].f.unused[3] );
tran (\sa_snapshot[4][52] , \sa_snapshot[4].r.part1[20] );
tran (\sa_snapshot[4][52] , \sa_snapshot[4].f.unused[2] );
tran (\sa_snapshot[4][51] , \sa_snapshot[4].r.part1[19] );
tran (\sa_snapshot[4][51] , \sa_snapshot[4].f.unused[1] );
tran (\sa_snapshot[4][50] , \sa_snapshot[4].r.part1[18] );
tran (\sa_snapshot[4][50] , \sa_snapshot[4].f.unused[0] );
tran (\sa_snapshot[4][49] , \sa_snapshot[4].r.part1[17] );
tran (\sa_snapshot[4][49] , \sa_snapshot[4].f.upper[17] );
tran (\sa_snapshot[4][48] , \sa_snapshot[4].r.part1[16] );
tran (\sa_snapshot[4][48] , \sa_snapshot[4].f.upper[16] );
tran (\sa_snapshot[4][47] , \sa_snapshot[4].r.part1[15] );
tran (\sa_snapshot[4][47] , \sa_snapshot[4].f.upper[15] );
tran (\sa_snapshot[4][46] , \sa_snapshot[4].r.part1[14] );
tran (\sa_snapshot[4][46] , \sa_snapshot[4].f.upper[14] );
tran (\sa_snapshot[4][45] , \sa_snapshot[4].r.part1[13] );
tran (\sa_snapshot[4][45] , \sa_snapshot[4].f.upper[13] );
tran (\sa_snapshot[4][44] , \sa_snapshot[4].r.part1[12] );
tran (\sa_snapshot[4][44] , \sa_snapshot[4].f.upper[12] );
tran (\sa_snapshot[4][43] , \sa_snapshot[4].r.part1[11] );
tran (\sa_snapshot[4][43] , \sa_snapshot[4].f.upper[11] );
tran (\sa_snapshot[4][42] , \sa_snapshot[4].r.part1[10] );
tran (\sa_snapshot[4][42] , \sa_snapshot[4].f.upper[10] );
tran (\sa_snapshot[4][41] , \sa_snapshot[4].r.part1[9] );
tran (\sa_snapshot[4][41] , \sa_snapshot[4].f.upper[9] );
tran (\sa_snapshot[4][40] , \sa_snapshot[4].r.part1[8] );
tran (\sa_snapshot[4][40] , \sa_snapshot[4].f.upper[8] );
tran (\sa_snapshot[4][39] , \sa_snapshot[4].r.part1[7] );
tran (\sa_snapshot[4][39] , \sa_snapshot[4].f.upper[7] );
tran (\sa_snapshot[4][38] , \sa_snapshot[4].r.part1[6] );
tran (\sa_snapshot[4][38] , \sa_snapshot[4].f.upper[6] );
tran (\sa_snapshot[4][37] , \sa_snapshot[4].r.part1[5] );
tran (\sa_snapshot[4][37] , \sa_snapshot[4].f.upper[5] );
tran (\sa_snapshot[4][36] , \sa_snapshot[4].r.part1[4] );
tran (\sa_snapshot[4][36] , \sa_snapshot[4].f.upper[4] );
tran (\sa_snapshot[4][35] , \sa_snapshot[4].r.part1[3] );
tran (\sa_snapshot[4][35] , \sa_snapshot[4].f.upper[3] );
tran (\sa_snapshot[4][34] , \sa_snapshot[4].r.part1[2] );
tran (\sa_snapshot[4][34] , \sa_snapshot[4].f.upper[2] );
tran (\sa_snapshot[4][33] , \sa_snapshot[4].r.part1[1] );
tran (\sa_snapshot[4][33] , \sa_snapshot[4].f.upper[1] );
tran (\sa_snapshot[4][32] , \sa_snapshot[4].r.part1[0] );
tran (\sa_snapshot[4][32] , \sa_snapshot[4].f.upper[0] );
tran (\sa_snapshot[4][31] , \sa_snapshot[4].r.part0[31] );
tran (\sa_snapshot[4][31] , \sa_snapshot[4].f.lower[31] );
tran (\sa_snapshot[4][30] , \sa_snapshot[4].r.part0[30] );
tran (\sa_snapshot[4][30] , \sa_snapshot[4].f.lower[30] );
tran (\sa_snapshot[4][29] , \sa_snapshot[4].r.part0[29] );
tran (\sa_snapshot[4][29] , \sa_snapshot[4].f.lower[29] );
tran (\sa_snapshot[4][28] , \sa_snapshot[4].r.part0[28] );
tran (\sa_snapshot[4][28] , \sa_snapshot[4].f.lower[28] );
tran (\sa_snapshot[4][27] , \sa_snapshot[4].r.part0[27] );
tran (\sa_snapshot[4][27] , \sa_snapshot[4].f.lower[27] );
tran (\sa_snapshot[4][26] , \sa_snapshot[4].r.part0[26] );
tran (\sa_snapshot[4][26] , \sa_snapshot[4].f.lower[26] );
tran (\sa_snapshot[4][25] , \sa_snapshot[4].r.part0[25] );
tran (\sa_snapshot[4][25] , \sa_snapshot[4].f.lower[25] );
tran (\sa_snapshot[4][24] , \sa_snapshot[4].r.part0[24] );
tran (\sa_snapshot[4][24] , \sa_snapshot[4].f.lower[24] );
tran (\sa_snapshot[4][23] , \sa_snapshot[4].r.part0[23] );
tran (\sa_snapshot[4][23] , \sa_snapshot[4].f.lower[23] );
tran (\sa_snapshot[4][22] , \sa_snapshot[4].r.part0[22] );
tran (\sa_snapshot[4][22] , \sa_snapshot[4].f.lower[22] );
tran (\sa_snapshot[4][21] , \sa_snapshot[4].r.part0[21] );
tran (\sa_snapshot[4][21] , \sa_snapshot[4].f.lower[21] );
tran (\sa_snapshot[4][20] , \sa_snapshot[4].r.part0[20] );
tran (\sa_snapshot[4][20] , \sa_snapshot[4].f.lower[20] );
tran (\sa_snapshot[4][19] , \sa_snapshot[4].r.part0[19] );
tran (\sa_snapshot[4][19] , \sa_snapshot[4].f.lower[19] );
tran (\sa_snapshot[4][18] , \sa_snapshot[4].r.part0[18] );
tran (\sa_snapshot[4][18] , \sa_snapshot[4].f.lower[18] );
tran (\sa_snapshot[4][17] , \sa_snapshot[4].r.part0[17] );
tran (\sa_snapshot[4][17] , \sa_snapshot[4].f.lower[17] );
tran (\sa_snapshot[4][16] , \sa_snapshot[4].r.part0[16] );
tran (\sa_snapshot[4][16] , \sa_snapshot[4].f.lower[16] );
tran (\sa_snapshot[4][15] , \sa_snapshot[4].r.part0[15] );
tran (\sa_snapshot[4][15] , \sa_snapshot[4].f.lower[15] );
tran (\sa_snapshot[4][14] , \sa_snapshot[4].r.part0[14] );
tran (\sa_snapshot[4][14] , \sa_snapshot[4].f.lower[14] );
tran (\sa_snapshot[4][13] , \sa_snapshot[4].r.part0[13] );
tran (\sa_snapshot[4][13] , \sa_snapshot[4].f.lower[13] );
tran (\sa_snapshot[4][12] , \sa_snapshot[4].r.part0[12] );
tran (\sa_snapshot[4][12] , \sa_snapshot[4].f.lower[12] );
tran (\sa_snapshot[4][11] , \sa_snapshot[4].r.part0[11] );
tran (\sa_snapshot[4][11] , \sa_snapshot[4].f.lower[11] );
tran (\sa_snapshot[4][10] , \sa_snapshot[4].r.part0[10] );
tran (\sa_snapshot[4][10] , \sa_snapshot[4].f.lower[10] );
tran (\sa_snapshot[4][9] , \sa_snapshot[4].r.part0[9] );
tran (\sa_snapshot[4][9] , \sa_snapshot[4].f.lower[9] );
tran (\sa_snapshot[4][8] , \sa_snapshot[4].r.part0[8] );
tran (\sa_snapshot[4][8] , \sa_snapshot[4].f.lower[8] );
tran (\sa_snapshot[4][7] , \sa_snapshot[4].r.part0[7] );
tran (\sa_snapshot[4][7] , \sa_snapshot[4].f.lower[7] );
tran (\sa_snapshot[4][6] , \sa_snapshot[4].r.part0[6] );
tran (\sa_snapshot[4][6] , \sa_snapshot[4].f.lower[6] );
tran (\sa_snapshot[4][5] , \sa_snapshot[4].r.part0[5] );
tran (\sa_snapshot[4][5] , \sa_snapshot[4].f.lower[5] );
tran (\sa_snapshot[4][4] , \sa_snapshot[4].r.part0[4] );
tran (\sa_snapshot[4][4] , \sa_snapshot[4].f.lower[4] );
tran (\sa_snapshot[4][3] , \sa_snapshot[4].r.part0[3] );
tran (\sa_snapshot[4][3] , \sa_snapshot[4].f.lower[3] );
tran (\sa_snapshot[4][2] , \sa_snapshot[4].r.part0[2] );
tran (\sa_snapshot[4][2] , \sa_snapshot[4].f.lower[2] );
tran (\sa_snapshot[4][1] , \sa_snapshot[4].r.part0[1] );
tran (\sa_snapshot[4][1] , \sa_snapshot[4].f.lower[1] );
tran (\sa_snapshot[4][0] , \sa_snapshot[4].r.part0[0] );
tran (\sa_snapshot[4][0] , \sa_snapshot[4].f.lower[0] );
tran (\sa_snapshot[3][63] , \sa_snapshot[3].r.part1[31] );
tran (\sa_snapshot[3][63] , \sa_snapshot[3].f.unused[13] );
tran (\sa_snapshot[3][62] , \sa_snapshot[3].r.part1[30] );
tran (\sa_snapshot[3][62] , \sa_snapshot[3].f.unused[12] );
tran (\sa_snapshot[3][61] , \sa_snapshot[3].r.part1[29] );
tran (\sa_snapshot[3][61] , \sa_snapshot[3].f.unused[11] );
tran (\sa_snapshot[3][60] , \sa_snapshot[3].r.part1[28] );
tran (\sa_snapshot[3][60] , \sa_snapshot[3].f.unused[10] );
tran (\sa_snapshot[3][59] , \sa_snapshot[3].r.part1[27] );
tran (\sa_snapshot[3][59] , \sa_snapshot[3].f.unused[9] );
tran (\sa_snapshot[3][58] , \sa_snapshot[3].r.part1[26] );
tran (\sa_snapshot[3][58] , \sa_snapshot[3].f.unused[8] );
tran (\sa_snapshot[3][57] , \sa_snapshot[3].r.part1[25] );
tran (\sa_snapshot[3][57] , \sa_snapshot[3].f.unused[7] );
tran (\sa_snapshot[3][56] , \sa_snapshot[3].r.part1[24] );
tran (\sa_snapshot[3][56] , \sa_snapshot[3].f.unused[6] );
tran (\sa_snapshot[3][55] , \sa_snapshot[3].r.part1[23] );
tran (\sa_snapshot[3][55] , \sa_snapshot[3].f.unused[5] );
tran (\sa_snapshot[3][54] , \sa_snapshot[3].r.part1[22] );
tran (\sa_snapshot[3][54] , \sa_snapshot[3].f.unused[4] );
tran (\sa_snapshot[3][53] , \sa_snapshot[3].r.part1[21] );
tran (\sa_snapshot[3][53] , \sa_snapshot[3].f.unused[3] );
tran (\sa_snapshot[3][52] , \sa_snapshot[3].r.part1[20] );
tran (\sa_snapshot[3][52] , \sa_snapshot[3].f.unused[2] );
tran (\sa_snapshot[3][51] , \sa_snapshot[3].r.part1[19] );
tran (\sa_snapshot[3][51] , \sa_snapshot[3].f.unused[1] );
tran (\sa_snapshot[3][50] , \sa_snapshot[3].r.part1[18] );
tran (\sa_snapshot[3][50] , \sa_snapshot[3].f.unused[0] );
tran (\sa_snapshot[3][49] , \sa_snapshot[3].r.part1[17] );
tran (\sa_snapshot[3][49] , \sa_snapshot[3].f.upper[17] );
tran (\sa_snapshot[3][48] , \sa_snapshot[3].r.part1[16] );
tran (\sa_snapshot[3][48] , \sa_snapshot[3].f.upper[16] );
tran (\sa_snapshot[3][47] , \sa_snapshot[3].r.part1[15] );
tran (\sa_snapshot[3][47] , \sa_snapshot[3].f.upper[15] );
tran (\sa_snapshot[3][46] , \sa_snapshot[3].r.part1[14] );
tran (\sa_snapshot[3][46] , \sa_snapshot[3].f.upper[14] );
tran (\sa_snapshot[3][45] , \sa_snapshot[3].r.part1[13] );
tran (\sa_snapshot[3][45] , \sa_snapshot[3].f.upper[13] );
tran (\sa_snapshot[3][44] , \sa_snapshot[3].r.part1[12] );
tran (\sa_snapshot[3][44] , \sa_snapshot[3].f.upper[12] );
tran (\sa_snapshot[3][43] , \sa_snapshot[3].r.part1[11] );
tran (\sa_snapshot[3][43] , \sa_snapshot[3].f.upper[11] );
tran (\sa_snapshot[3][42] , \sa_snapshot[3].r.part1[10] );
tran (\sa_snapshot[3][42] , \sa_snapshot[3].f.upper[10] );
tran (\sa_snapshot[3][41] , \sa_snapshot[3].r.part1[9] );
tran (\sa_snapshot[3][41] , \sa_snapshot[3].f.upper[9] );
tran (\sa_snapshot[3][40] , \sa_snapshot[3].r.part1[8] );
tran (\sa_snapshot[3][40] , \sa_snapshot[3].f.upper[8] );
tran (\sa_snapshot[3][39] , \sa_snapshot[3].r.part1[7] );
tran (\sa_snapshot[3][39] , \sa_snapshot[3].f.upper[7] );
tran (\sa_snapshot[3][38] , \sa_snapshot[3].r.part1[6] );
tran (\sa_snapshot[3][38] , \sa_snapshot[3].f.upper[6] );
tran (\sa_snapshot[3][37] , \sa_snapshot[3].r.part1[5] );
tran (\sa_snapshot[3][37] , \sa_snapshot[3].f.upper[5] );
tran (\sa_snapshot[3][36] , \sa_snapshot[3].r.part1[4] );
tran (\sa_snapshot[3][36] , \sa_snapshot[3].f.upper[4] );
tran (\sa_snapshot[3][35] , \sa_snapshot[3].r.part1[3] );
tran (\sa_snapshot[3][35] , \sa_snapshot[3].f.upper[3] );
tran (\sa_snapshot[3][34] , \sa_snapshot[3].r.part1[2] );
tran (\sa_snapshot[3][34] , \sa_snapshot[3].f.upper[2] );
tran (\sa_snapshot[3][33] , \sa_snapshot[3].r.part1[1] );
tran (\sa_snapshot[3][33] , \sa_snapshot[3].f.upper[1] );
tran (\sa_snapshot[3][32] , \sa_snapshot[3].r.part1[0] );
tran (\sa_snapshot[3][32] , \sa_snapshot[3].f.upper[0] );
tran (\sa_snapshot[3][31] , \sa_snapshot[3].r.part0[31] );
tran (\sa_snapshot[3][31] , \sa_snapshot[3].f.lower[31] );
tran (\sa_snapshot[3][30] , \sa_snapshot[3].r.part0[30] );
tran (\sa_snapshot[3][30] , \sa_snapshot[3].f.lower[30] );
tran (\sa_snapshot[3][29] , \sa_snapshot[3].r.part0[29] );
tran (\sa_snapshot[3][29] , \sa_snapshot[3].f.lower[29] );
tran (\sa_snapshot[3][28] , \sa_snapshot[3].r.part0[28] );
tran (\sa_snapshot[3][28] , \sa_snapshot[3].f.lower[28] );
tran (\sa_snapshot[3][27] , \sa_snapshot[3].r.part0[27] );
tran (\sa_snapshot[3][27] , \sa_snapshot[3].f.lower[27] );
tran (\sa_snapshot[3][26] , \sa_snapshot[3].r.part0[26] );
tran (\sa_snapshot[3][26] , \sa_snapshot[3].f.lower[26] );
tran (\sa_snapshot[3][25] , \sa_snapshot[3].r.part0[25] );
tran (\sa_snapshot[3][25] , \sa_snapshot[3].f.lower[25] );
tran (\sa_snapshot[3][24] , \sa_snapshot[3].r.part0[24] );
tran (\sa_snapshot[3][24] , \sa_snapshot[3].f.lower[24] );
tran (\sa_snapshot[3][23] , \sa_snapshot[3].r.part0[23] );
tran (\sa_snapshot[3][23] , \sa_snapshot[3].f.lower[23] );
tran (\sa_snapshot[3][22] , \sa_snapshot[3].r.part0[22] );
tran (\sa_snapshot[3][22] , \sa_snapshot[3].f.lower[22] );
tran (\sa_snapshot[3][21] , \sa_snapshot[3].r.part0[21] );
tran (\sa_snapshot[3][21] , \sa_snapshot[3].f.lower[21] );
tran (\sa_snapshot[3][20] , \sa_snapshot[3].r.part0[20] );
tran (\sa_snapshot[3][20] , \sa_snapshot[3].f.lower[20] );
tran (\sa_snapshot[3][19] , \sa_snapshot[3].r.part0[19] );
tran (\sa_snapshot[3][19] , \sa_snapshot[3].f.lower[19] );
tran (\sa_snapshot[3][18] , \sa_snapshot[3].r.part0[18] );
tran (\sa_snapshot[3][18] , \sa_snapshot[3].f.lower[18] );
tran (\sa_snapshot[3][17] , \sa_snapshot[3].r.part0[17] );
tran (\sa_snapshot[3][17] , \sa_snapshot[3].f.lower[17] );
tran (\sa_snapshot[3][16] , \sa_snapshot[3].r.part0[16] );
tran (\sa_snapshot[3][16] , \sa_snapshot[3].f.lower[16] );
tran (\sa_snapshot[3][15] , \sa_snapshot[3].r.part0[15] );
tran (\sa_snapshot[3][15] , \sa_snapshot[3].f.lower[15] );
tran (\sa_snapshot[3][14] , \sa_snapshot[3].r.part0[14] );
tran (\sa_snapshot[3][14] , \sa_snapshot[3].f.lower[14] );
tran (\sa_snapshot[3][13] , \sa_snapshot[3].r.part0[13] );
tran (\sa_snapshot[3][13] , \sa_snapshot[3].f.lower[13] );
tran (\sa_snapshot[3][12] , \sa_snapshot[3].r.part0[12] );
tran (\sa_snapshot[3][12] , \sa_snapshot[3].f.lower[12] );
tran (\sa_snapshot[3][11] , \sa_snapshot[3].r.part0[11] );
tran (\sa_snapshot[3][11] , \sa_snapshot[3].f.lower[11] );
tran (\sa_snapshot[3][10] , \sa_snapshot[3].r.part0[10] );
tran (\sa_snapshot[3][10] , \sa_snapshot[3].f.lower[10] );
tran (\sa_snapshot[3][9] , \sa_snapshot[3].r.part0[9] );
tran (\sa_snapshot[3][9] , \sa_snapshot[3].f.lower[9] );
tran (\sa_snapshot[3][8] , \sa_snapshot[3].r.part0[8] );
tran (\sa_snapshot[3][8] , \sa_snapshot[3].f.lower[8] );
tran (\sa_snapshot[3][7] , \sa_snapshot[3].r.part0[7] );
tran (\sa_snapshot[3][7] , \sa_snapshot[3].f.lower[7] );
tran (\sa_snapshot[3][6] , \sa_snapshot[3].r.part0[6] );
tran (\sa_snapshot[3][6] , \sa_snapshot[3].f.lower[6] );
tran (\sa_snapshot[3][5] , \sa_snapshot[3].r.part0[5] );
tran (\sa_snapshot[3][5] , \sa_snapshot[3].f.lower[5] );
tran (\sa_snapshot[3][4] , \sa_snapshot[3].r.part0[4] );
tran (\sa_snapshot[3][4] , \sa_snapshot[3].f.lower[4] );
tran (\sa_snapshot[3][3] , \sa_snapshot[3].r.part0[3] );
tran (\sa_snapshot[3][3] , \sa_snapshot[3].f.lower[3] );
tran (\sa_snapshot[3][2] , \sa_snapshot[3].r.part0[2] );
tran (\sa_snapshot[3][2] , \sa_snapshot[3].f.lower[2] );
tran (\sa_snapshot[3][1] , \sa_snapshot[3].r.part0[1] );
tran (\sa_snapshot[3][1] , \sa_snapshot[3].f.lower[1] );
tran (\sa_snapshot[3][0] , \sa_snapshot[3].r.part0[0] );
tran (\sa_snapshot[3][0] , \sa_snapshot[3].f.lower[0] );
tran (\sa_snapshot[2][63] , \sa_snapshot[2].r.part1[31] );
tran (\sa_snapshot[2][63] , \sa_snapshot[2].f.unused[13] );
tran (\sa_snapshot[2][62] , \sa_snapshot[2].r.part1[30] );
tran (\sa_snapshot[2][62] , \sa_snapshot[2].f.unused[12] );
tran (\sa_snapshot[2][61] , \sa_snapshot[2].r.part1[29] );
tran (\sa_snapshot[2][61] , \sa_snapshot[2].f.unused[11] );
tran (\sa_snapshot[2][60] , \sa_snapshot[2].r.part1[28] );
tran (\sa_snapshot[2][60] , \sa_snapshot[2].f.unused[10] );
tran (\sa_snapshot[2][59] , \sa_snapshot[2].r.part1[27] );
tran (\sa_snapshot[2][59] , \sa_snapshot[2].f.unused[9] );
tran (\sa_snapshot[2][58] , \sa_snapshot[2].r.part1[26] );
tran (\sa_snapshot[2][58] , \sa_snapshot[2].f.unused[8] );
tran (\sa_snapshot[2][57] , \sa_snapshot[2].r.part1[25] );
tran (\sa_snapshot[2][57] , \sa_snapshot[2].f.unused[7] );
tran (\sa_snapshot[2][56] , \sa_snapshot[2].r.part1[24] );
tran (\sa_snapshot[2][56] , \sa_snapshot[2].f.unused[6] );
tran (\sa_snapshot[2][55] , \sa_snapshot[2].r.part1[23] );
tran (\sa_snapshot[2][55] , \sa_snapshot[2].f.unused[5] );
tran (\sa_snapshot[2][54] , \sa_snapshot[2].r.part1[22] );
tran (\sa_snapshot[2][54] , \sa_snapshot[2].f.unused[4] );
tran (\sa_snapshot[2][53] , \sa_snapshot[2].r.part1[21] );
tran (\sa_snapshot[2][53] , \sa_snapshot[2].f.unused[3] );
tran (\sa_snapshot[2][52] , \sa_snapshot[2].r.part1[20] );
tran (\sa_snapshot[2][52] , \sa_snapshot[2].f.unused[2] );
tran (\sa_snapshot[2][51] , \sa_snapshot[2].r.part1[19] );
tran (\sa_snapshot[2][51] , \sa_snapshot[2].f.unused[1] );
tran (\sa_snapshot[2][50] , \sa_snapshot[2].r.part1[18] );
tran (\sa_snapshot[2][50] , \sa_snapshot[2].f.unused[0] );
tran (\sa_snapshot[2][49] , \sa_snapshot[2].r.part1[17] );
tran (\sa_snapshot[2][49] , \sa_snapshot[2].f.upper[17] );
tran (\sa_snapshot[2][48] , \sa_snapshot[2].r.part1[16] );
tran (\sa_snapshot[2][48] , \sa_snapshot[2].f.upper[16] );
tran (\sa_snapshot[2][47] , \sa_snapshot[2].r.part1[15] );
tran (\sa_snapshot[2][47] , \sa_snapshot[2].f.upper[15] );
tran (\sa_snapshot[2][46] , \sa_snapshot[2].r.part1[14] );
tran (\sa_snapshot[2][46] , \sa_snapshot[2].f.upper[14] );
tran (\sa_snapshot[2][45] , \sa_snapshot[2].r.part1[13] );
tran (\sa_snapshot[2][45] , \sa_snapshot[2].f.upper[13] );
tran (\sa_snapshot[2][44] , \sa_snapshot[2].r.part1[12] );
tran (\sa_snapshot[2][44] , \sa_snapshot[2].f.upper[12] );
tran (\sa_snapshot[2][43] , \sa_snapshot[2].r.part1[11] );
tran (\sa_snapshot[2][43] , \sa_snapshot[2].f.upper[11] );
tran (\sa_snapshot[2][42] , \sa_snapshot[2].r.part1[10] );
tran (\sa_snapshot[2][42] , \sa_snapshot[2].f.upper[10] );
tran (\sa_snapshot[2][41] , \sa_snapshot[2].r.part1[9] );
tran (\sa_snapshot[2][41] , \sa_snapshot[2].f.upper[9] );
tran (\sa_snapshot[2][40] , \sa_snapshot[2].r.part1[8] );
tran (\sa_snapshot[2][40] , \sa_snapshot[2].f.upper[8] );
tran (\sa_snapshot[2][39] , \sa_snapshot[2].r.part1[7] );
tran (\sa_snapshot[2][39] , \sa_snapshot[2].f.upper[7] );
tran (\sa_snapshot[2][38] , \sa_snapshot[2].r.part1[6] );
tran (\sa_snapshot[2][38] , \sa_snapshot[2].f.upper[6] );
tran (\sa_snapshot[2][37] , \sa_snapshot[2].r.part1[5] );
tran (\sa_snapshot[2][37] , \sa_snapshot[2].f.upper[5] );
tran (\sa_snapshot[2][36] , \sa_snapshot[2].r.part1[4] );
tran (\sa_snapshot[2][36] , \sa_snapshot[2].f.upper[4] );
tran (\sa_snapshot[2][35] , \sa_snapshot[2].r.part1[3] );
tran (\sa_snapshot[2][35] , \sa_snapshot[2].f.upper[3] );
tran (\sa_snapshot[2][34] , \sa_snapshot[2].r.part1[2] );
tran (\sa_snapshot[2][34] , \sa_snapshot[2].f.upper[2] );
tran (\sa_snapshot[2][33] , \sa_snapshot[2].r.part1[1] );
tran (\sa_snapshot[2][33] , \sa_snapshot[2].f.upper[1] );
tran (\sa_snapshot[2][32] , \sa_snapshot[2].r.part1[0] );
tran (\sa_snapshot[2][32] , \sa_snapshot[2].f.upper[0] );
tran (\sa_snapshot[2][31] , \sa_snapshot[2].r.part0[31] );
tran (\sa_snapshot[2][31] , \sa_snapshot[2].f.lower[31] );
tran (\sa_snapshot[2][30] , \sa_snapshot[2].r.part0[30] );
tran (\sa_snapshot[2][30] , \sa_snapshot[2].f.lower[30] );
tran (\sa_snapshot[2][29] , \sa_snapshot[2].r.part0[29] );
tran (\sa_snapshot[2][29] , \sa_snapshot[2].f.lower[29] );
tran (\sa_snapshot[2][28] , \sa_snapshot[2].r.part0[28] );
tran (\sa_snapshot[2][28] , \sa_snapshot[2].f.lower[28] );
tran (\sa_snapshot[2][27] , \sa_snapshot[2].r.part0[27] );
tran (\sa_snapshot[2][27] , \sa_snapshot[2].f.lower[27] );
tran (\sa_snapshot[2][26] , \sa_snapshot[2].r.part0[26] );
tran (\sa_snapshot[2][26] , \sa_snapshot[2].f.lower[26] );
tran (\sa_snapshot[2][25] , \sa_snapshot[2].r.part0[25] );
tran (\sa_snapshot[2][25] , \sa_snapshot[2].f.lower[25] );
tran (\sa_snapshot[2][24] , \sa_snapshot[2].r.part0[24] );
tran (\sa_snapshot[2][24] , \sa_snapshot[2].f.lower[24] );
tran (\sa_snapshot[2][23] , \sa_snapshot[2].r.part0[23] );
tran (\sa_snapshot[2][23] , \sa_snapshot[2].f.lower[23] );
tran (\sa_snapshot[2][22] , \sa_snapshot[2].r.part0[22] );
tran (\sa_snapshot[2][22] , \sa_snapshot[2].f.lower[22] );
tran (\sa_snapshot[2][21] , \sa_snapshot[2].r.part0[21] );
tran (\sa_snapshot[2][21] , \sa_snapshot[2].f.lower[21] );
tran (\sa_snapshot[2][20] , \sa_snapshot[2].r.part0[20] );
tran (\sa_snapshot[2][20] , \sa_snapshot[2].f.lower[20] );
tran (\sa_snapshot[2][19] , \sa_snapshot[2].r.part0[19] );
tran (\sa_snapshot[2][19] , \sa_snapshot[2].f.lower[19] );
tran (\sa_snapshot[2][18] , \sa_snapshot[2].r.part0[18] );
tran (\sa_snapshot[2][18] , \sa_snapshot[2].f.lower[18] );
tran (\sa_snapshot[2][17] , \sa_snapshot[2].r.part0[17] );
tran (\sa_snapshot[2][17] , \sa_snapshot[2].f.lower[17] );
tran (\sa_snapshot[2][16] , \sa_snapshot[2].r.part0[16] );
tran (\sa_snapshot[2][16] , \sa_snapshot[2].f.lower[16] );
tran (\sa_snapshot[2][15] , \sa_snapshot[2].r.part0[15] );
tran (\sa_snapshot[2][15] , \sa_snapshot[2].f.lower[15] );
tran (\sa_snapshot[2][14] , \sa_snapshot[2].r.part0[14] );
tran (\sa_snapshot[2][14] , \sa_snapshot[2].f.lower[14] );
tran (\sa_snapshot[2][13] , \sa_snapshot[2].r.part0[13] );
tran (\sa_snapshot[2][13] , \sa_snapshot[2].f.lower[13] );
tran (\sa_snapshot[2][12] , \sa_snapshot[2].r.part0[12] );
tran (\sa_snapshot[2][12] , \sa_snapshot[2].f.lower[12] );
tran (\sa_snapshot[2][11] , \sa_snapshot[2].r.part0[11] );
tran (\sa_snapshot[2][11] , \sa_snapshot[2].f.lower[11] );
tran (\sa_snapshot[2][10] , \sa_snapshot[2].r.part0[10] );
tran (\sa_snapshot[2][10] , \sa_snapshot[2].f.lower[10] );
tran (\sa_snapshot[2][9] , \sa_snapshot[2].r.part0[9] );
tran (\sa_snapshot[2][9] , \sa_snapshot[2].f.lower[9] );
tran (\sa_snapshot[2][8] , \sa_snapshot[2].r.part0[8] );
tran (\sa_snapshot[2][8] , \sa_snapshot[2].f.lower[8] );
tran (\sa_snapshot[2][7] , \sa_snapshot[2].r.part0[7] );
tran (\sa_snapshot[2][7] , \sa_snapshot[2].f.lower[7] );
tran (\sa_snapshot[2][6] , \sa_snapshot[2].r.part0[6] );
tran (\sa_snapshot[2][6] , \sa_snapshot[2].f.lower[6] );
tran (\sa_snapshot[2][5] , \sa_snapshot[2].r.part0[5] );
tran (\sa_snapshot[2][5] , \sa_snapshot[2].f.lower[5] );
tran (\sa_snapshot[2][4] , \sa_snapshot[2].r.part0[4] );
tran (\sa_snapshot[2][4] , \sa_snapshot[2].f.lower[4] );
tran (\sa_snapshot[2][3] , \sa_snapshot[2].r.part0[3] );
tran (\sa_snapshot[2][3] , \sa_snapshot[2].f.lower[3] );
tran (\sa_snapshot[2][2] , \sa_snapshot[2].r.part0[2] );
tran (\sa_snapshot[2][2] , \sa_snapshot[2].f.lower[2] );
tran (\sa_snapshot[2][1] , \sa_snapshot[2].r.part0[1] );
tran (\sa_snapshot[2][1] , \sa_snapshot[2].f.lower[1] );
tran (\sa_snapshot[2][0] , \sa_snapshot[2].r.part0[0] );
tran (\sa_snapshot[2][0] , \sa_snapshot[2].f.lower[0] );
tran (\sa_snapshot[1][63] , \sa_snapshot[1].r.part1[31] );
tran (\sa_snapshot[1][63] , \sa_snapshot[1].f.unused[13] );
tran (\sa_snapshot[1][62] , \sa_snapshot[1].r.part1[30] );
tran (\sa_snapshot[1][62] , \sa_snapshot[1].f.unused[12] );
tran (\sa_snapshot[1][61] , \sa_snapshot[1].r.part1[29] );
tran (\sa_snapshot[1][61] , \sa_snapshot[1].f.unused[11] );
tran (\sa_snapshot[1][60] , \sa_snapshot[1].r.part1[28] );
tran (\sa_snapshot[1][60] , \sa_snapshot[1].f.unused[10] );
tran (\sa_snapshot[1][59] , \sa_snapshot[1].r.part1[27] );
tran (\sa_snapshot[1][59] , \sa_snapshot[1].f.unused[9] );
tran (\sa_snapshot[1][58] , \sa_snapshot[1].r.part1[26] );
tran (\sa_snapshot[1][58] , \sa_snapshot[1].f.unused[8] );
tran (\sa_snapshot[1][57] , \sa_snapshot[1].r.part1[25] );
tran (\sa_snapshot[1][57] , \sa_snapshot[1].f.unused[7] );
tran (\sa_snapshot[1][56] , \sa_snapshot[1].r.part1[24] );
tran (\sa_snapshot[1][56] , \sa_snapshot[1].f.unused[6] );
tran (\sa_snapshot[1][55] , \sa_snapshot[1].r.part1[23] );
tran (\sa_snapshot[1][55] , \sa_snapshot[1].f.unused[5] );
tran (\sa_snapshot[1][54] , \sa_snapshot[1].r.part1[22] );
tran (\sa_snapshot[1][54] , \sa_snapshot[1].f.unused[4] );
tran (\sa_snapshot[1][53] , \sa_snapshot[1].r.part1[21] );
tran (\sa_snapshot[1][53] , \sa_snapshot[1].f.unused[3] );
tran (\sa_snapshot[1][52] , \sa_snapshot[1].r.part1[20] );
tran (\sa_snapshot[1][52] , \sa_snapshot[1].f.unused[2] );
tran (\sa_snapshot[1][51] , \sa_snapshot[1].r.part1[19] );
tran (\sa_snapshot[1][51] , \sa_snapshot[1].f.unused[1] );
tran (\sa_snapshot[1][50] , \sa_snapshot[1].r.part1[18] );
tran (\sa_snapshot[1][50] , \sa_snapshot[1].f.unused[0] );
tran (\sa_snapshot[1][49] , \sa_snapshot[1].r.part1[17] );
tran (\sa_snapshot[1][49] , \sa_snapshot[1].f.upper[17] );
tran (\sa_snapshot[1][48] , \sa_snapshot[1].r.part1[16] );
tran (\sa_snapshot[1][48] , \sa_snapshot[1].f.upper[16] );
tran (\sa_snapshot[1][47] , \sa_snapshot[1].r.part1[15] );
tran (\sa_snapshot[1][47] , \sa_snapshot[1].f.upper[15] );
tran (\sa_snapshot[1][46] , \sa_snapshot[1].r.part1[14] );
tran (\sa_snapshot[1][46] , \sa_snapshot[1].f.upper[14] );
tran (\sa_snapshot[1][45] , \sa_snapshot[1].r.part1[13] );
tran (\sa_snapshot[1][45] , \sa_snapshot[1].f.upper[13] );
tran (\sa_snapshot[1][44] , \sa_snapshot[1].r.part1[12] );
tran (\sa_snapshot[1][44] , \sa_snapshot[1].f.upper[12] );
tran (\sa_snapshot[1][43] , \sa_snapshot[1].r.part1[11] );
tran (\sa_snapshot[1][43] , \sa_snapshot[1].f.upper[11] );
tran (\sa_snapshot[1][42] , \sa_snapshot[1].r.part1[10] );
tran (\sa_snapshot[1][42] , \sa_snapshot[1].f.upper[10] );
tran (\sa_snapshot[1][41] , \sa_snapshot[1].r.part1[9] );
tran (\sa_snapshot[1][41] , \sa_snapshot[1].f.upper[9] );
tran (\sa_snapshot[1][40] , \sa_snapshot[1].r.part1[8] );
tran (\sa_snapshot[1][40] , \sa_snapshot[1].f.upper[8] );
tran (\sa_snapshot[1][39] , \sa_snapshot[1].r.part1[7] );
tran (\sa_snapshot[1][39] , \sa_snapshot[1].f.upper[7] );
tran (\sa_snapshot[1][38] , \sa_snapshot[1].r.part1[6] );
tran (\sa_snapshot[1][38] , \sa_snapshot[1].f.upper[6] );
tran (\sa_snapshot[1][37] , \sa_snapshot[1].r.part1[5] );
tran (\sa_snapshot[1][37] , \sa_snapshot[1].f.upper[5] );
tran (\sa_snapshot[1][36] , \sa_snapshot[1].r.part1[4] );
tran (\sa_snapshot[1][36] , \sa_snapshot[1].f.upper[4] );
tran (\sa_snapshot[1][35] , \sa_snapshot[1].r.part1[3] );
tran (\sa_snapshot[1][35] , \sa_snapshot[1].f.upper[3] );
tran (\sa_snapshot[1][34] , \sa_snapshot[1].r.part1[2] );
tran (\sa_snapshot[1][34] , \sa_snapshot[1].f.upper[2] );
tran (\sa_snapshot[1][33] , \sa_snapshot[1].r.part1[1] );
tran (\sa_snapshot[1][33] , \sa_snapshot[1].f.upper[1] );
tran (\sa_snapshot[1][32] , \sa_snapshot[1].r.part1[0] );
tran (\sa_snapshot[1][32] , \sa_snapshot[1].f.upper[0] );
tran (\sa_snapshot[1][31] , \sa_snapshot[1].r.part0[31] );
tran (\sa_snapshot[1][31] , \sa_snapshot[1].f.lower[31] );
tran (\sa_snapshot[1][30] , \sa_snapshot[1].r.part0[30] );
tran (\sa_snapshot[1][30] , \sa_snapshot[1].f.lower[30] );
tran (\sa_snapshot[1][29] , \sa_snapshot[1].r.part0[29] );
tran (\sa_snapshot[1][29] , \sa_snapshot[1].f.lower[29] );
tran (\sa_snapshot[1][28] , \sa_snapshot[1].r.part0[28] );
tran (\sa_snapshot[1][28] , \sa_snapshot[1].f.lower[28] );
tran (\sa_snapshot[1][27] , \sa_snapshot[1].r.part0[27] );
tran (\sa_snapshot[1][27] , \sa_snapshot[1].f.lower[27] );
tran (\sa_snapshot[1][26] , \sa_snapshot[1].r.part0[26] );
tran (\sa_snapshot[1][26] , \sa_snapshot[1].f.lower[26] );
tran (\sa_snapshot[1][25] , \sa_snapshot[1].r.part0[25] );
tran (\sa_snapshot[1][25] , \sa_snapshot[1].f.lower[25] );
tran (\sa_snapshot[1][24] , \sa_snapshot[1].r.part0[24] );
tran (\sa_snapshot[1][24] , \sa_snapshot[1].f.lower[24] );
tran (\sa_snapshot[1][23] , \sa_snapshot[1].r.part0[23] );
tran (\sa_snapshot[1][23] , \sa_snapshot[1].f.lower[23] );
tran (\sa_snapshot[1][22] , \sa_snapshot[1].r.part0[22] );
tran (\sa_snapshot[1][22] , \sa_snapshot[1].f.lower[22] );
tran (\sa_snapshot[1][21] , \sa_snapshot[1].r.part0[21] );
tran (\sa_snapshot[1][21] , \sa_snapshot[1].f.lower[21] );
tran (\sa_snapshot[1][20] , \sa_snapshot[1].r.part0[20] );
tran (\sa_snapshot[1][20] , \sa_snapshot[1].f.lower[20] );
tran (\sa_snapshot[1][19] , \sa_snapshot[1].r.part0[19] );
tran (\sa_snapshot[1][19] , \sa_snapshot[1].f.lower[19] );
tran (\sa_snapshot[1][18] , \sa_snapshot[1].r.part0[18] );
tran (\sa_snapshot[1][18] , \sa_snapshot[1].f.lower[18] );
tran (\sa_snapshot[1][17] , \sa_snapshot[1].r.part0[17] );
tran (\sa_snapshot[1][17] , \sa_snapshot[1].f.lower[17] );
tran (\sa_snapshot[1][16] , \sa_snapshot[1].r.part0[16] );
tran (\sa_snapshot[1][16] , \sa_snapshot[1].f.lower[16] );
tran (\sa_snapshot[1][15] , \sa_snapshot[1].r.part0[15] );
tran (\sa_snapshot[1][15] , \sa_snapshot[1].f.lower[15] );
tran (\sa_snapshot[1][14] , \sa_snapshot[1].r.part0[14] );
tran (\sa_snapshot[1][14] , \sa_snapshot[1].f.lower[14] );
tran (\sa_snapshot[1][13] , \sa_snapshot[1].r.part0[13] );
tran (\sa_snapshot[1][13] , \sa_snapshot[1].f.lower[13] );
tran (\sa_snapshot[1][12] , \sa_snapshot[1].r.part0[12] );
tran (\sa_snapshot[1][12] , \sa_snapshot[1].f.lower[12] );
tran (\sa_snapshot[1][11] , \sa_snapshot[1].r.part0[11] );
tran (\sa_snapshot[1][11] , \sa_snapshot[1].f.lower[11] );
tran (\sa_snapshot[1][10] , \sa_snapshot[1].r.part0[10] );
tran (\sa_snapshot[1][10] , \sa_snapshot[1].f.lower[10] );
tran (\sa_snapshot[1][9] , \sa_snapshot[1].r.part0[9] );
tran (\sa_snapshot[1][9] , \sa_snapshot[1].f.lower[9] );
tran (\sa_snapshot[1][8] , \sa_snapshot[1].r.part0[8] );
tran (\sa_snapshot[1][8] , \sa_snapshot[1].f.lower[8] );
tran (\sa_snapshot[1][7] , \sa_snapshot[1].r.part0[7] );
tran (\sa_snapshot[1][7] , \sa_snapshot[1].f.lower[7] );
tran (\sa_snapshot[1][6] , \sa_snapshot[1].r.part0[6] );
tran (\sa_snapshot[1][6] , \sa_snapshot[1].f.lower[6] );
tran (\sa_snapshot[1][5] , \sa_snapshot[1].r.part0[5] );
tran (\sa_snapshot[1][5] , \sa_snapshot[1].f.lower[5] );
tran (\sa_snapshot[1][4] , \sa_snapshot[1].r.part0[4] );
tran (\sa_snapshot[1][4] , \sa_snapshot[1].f.lower[4] );
tran (\sa_snapshot[1][3] , \sa_snapshot[1].r.part0[3] );
tran (\sa_snapshot[1][3] , \sa_snapshot[1].f.lower[3] );
tran (\sa_snapshot[1][2] , \sa_snapshot[1].r.part0[2] );
tran (\sa_snapshot[1][2] , \sa_snapshot[1].f.lower[2] );
tran (\sa_snapshot[1][1] , \sa_snapshot[1].r.part0[1] );
tran (\sa_snapshot[1][1] , \sa_snapshot[1].f.lower[1] );
tran (\sa_snapshot[1][0] , \sa_snapshot[1].r.part0[0] );
tran (\sa_snapshot[1][0] , \sa_snapshot[1].f.lower[0] );
tran (\sa_snapshot[0][63] , \sa_snapshot[0].r.part1[31] );
tran (\sa_snapshot[0][63] , \sa_snapshot[0].f.unused[13] );
tran (\sa_snapshot[0][62] , \sa_snapshot[0].r.part1[30] );
tran (\sa_snapshot[0][62] , \sa_snapshot[0].f.unused[12] );
tran (\sa_snapshot[0][61] , \sa_snapshot[0].r.part1[29] );
tran (\sa_snapshot[0][61] , \sa_snapshot[0].f.unused[11] );
tran (\sa_snapshot[0][60] , \sa_snapshot[0].r.part1[28] );
tran (\sa_snapshot[0][60] , \sa_snapshot[0].f.unused[10] );
tran (\sa_snapshot[0][59] , \sa_snapshot[0].r.part1[27] );
tran (\sa_snapshot[0][59] , \sa_snapshot[0].f.unused[9] );
tran (\sa_snapshot[0][58] , \sa_snapshot[0].r.part1[26] );
tran (\sa_snapshot[0][58] , \sa_snapshot[0].f.unused[8] );
tran (\sa_snapshot[0][57] , \sa_snapshot[0].r.part1[25] );
tran (\sa_snapshot[0][57] , \sa_snapshot[0].f.unused[7] );
tran (\sa_snapshot[0][56] , \sa_snapshot[0].r.part1[24] );
tran (\sa_snapshot[0][56] , \sa_snapshot[0].f.unused[6] );
tran (\sa_snapshot[0][55] , \sa_snapshot[0].r.part1[23] );
tran (\sa_snapshot[0][55] , \sa_snapshot[0].f.unused[5] );
tran (\sa_snapshot[0][54] , \sa_snapshot[0].r.part1[22] );
tran (\sa_snapshot[0][54] , \sa_snapshot[0].f.unused[4] );
tran (\sa_snapshot[0][53] , \sa_snapshot[0].r.part1[21] );
tran (\sa_snapshot[0][53] , \sa_snapshot[0].f.unused[3] );
tran (\sa_snapshot[0][52] , \sa_snapshot[0].r.part1[20] );
tran (\sa_snapshot[0][52] , \sa_snapshot[0].f.unused[2] );
tran (\sa_snapshot[0][51] , \sa_snapshot[0].r.part1[19] );
tran (\sa_snapshot[0][51] , \sa_snapshot[0].f.unused[1] );
tran (\sa_snapshot[0][50] , \sa_snapshot[0].r.part1[18] );
tran (\sa_snapshot[0][50] , \sa_snapshot[0].f.unused[0] );
tran (\sa_snapshot[0][49] , \sa_snapshot[0].r.part1[17] );
tran (\sa_snapshot[0][49] , \sa_snapshot[0].f.upper[17] );
tran (\sa_snapshot[0][48] , \sa_snapshot[0].r.part1[16] );
tran (\sa_snapshot[0][48] , \sa_snapshot[0].f.upper[16] );
tran (\sa_snapshot[0][47] , \sa_snapshot[0].r.part1[15] );
tran (\sa_snapshot[0][47] , \sa_snapshot[0].f.upper[15] );
tran (\sa_snapshot[0][46] , \sa_snapshot[0].r.part1[14] );
tran (\sa_snapshot[0][46] , \sa_snapshot[0].f.upper[14] );
tran (\sa_snapshot[0][45] , \sa_snapshot[0].r.part1[13] );
tran (\sa_snapshot[0][45] , \sa_snapshot[0].f.upper[13] );
tran (\sa_snapshot[0][44] , \sa_snapshot[0].r.part1[12] );
tran (\sa_snapshot[0][44] , \sa_snapshot[0].f.upper[12] );
tran (\sa_snapshot[0][43] , \sa_snapshot[0].r.part1[11] );
tran (\sa_snapshot[0][43] , \sa_snapshot[0].f.upper[11] );
tran (\sa_snapshot[0][42] , \sa_snapshot[0].r.part1[10] );
tran (\sa_snapshot[0][42] , \sa_snapshot[0].f.upper[10] );
tran (\sa_snapshot[0][41] , \sa_snapshot[0].r.part1[9] );
tran (\sa_snapshot[0][41] , \sa_snapshot[0].f.upper[9] );
tran (\sa_snapshot[0][40] , \sa_snapshot[0].r.part1[8] );
tran (\sa_snapshot[0][40] , \sa_snapshot[0].f.upper[8] );
tran (\sa_snapshot[0][39] , \sa_snapshot[0].r.part1[7] );
tran (\sa_snapshot[0][39] , \sa_snapshot[0].f.upper[7] );
tran (\sa_snapshot[0][38] , \sa_snapshot[0].r.part1[6] );
tran (\sa_snapshot[0][38] , \sa_snapshot[0].f.upper[6] );
tran (\sa_snapshot[0][37] , \sa_snapshot[0].r.part1[5] );
tran (\sa_snapshot[0][37] , \sa_snapshot[0].f.upper[5] );
tran (\sa_snapshot[0][36] , \sa_snapshot[0].r.part1[4] );
tran (\sa_snapshot[0][36] , \sa_snapshot[0].f.upper[4] );
tran (\sa_snapshot[0][35] , \sa_snapshot[0].r.part1[3] );
tran (\sa_snapshot[0][35] , \sa_snapshot[0].f.upper[3] );
tran (\sa_snapshot[0][34] , \sa_snapshot[0].r.part1[2] );
tran (\sa_snapshot[0][34] , \sa_snapshot[0].f.upper[2] );
tran (\sa_snapshot[0][33] , \sa_snapshot[0].r.part1[1] );
tran (\sa_snapshot[0][33] , \sa_snapshot[0].f.upper[1] );
tran (\sa_snapshot[0][32] , \sa_snapshot[0].r.part1[0] );
tran (\sa_snapshot[0][32] , \sa_snapshot[0].f.upper[0] );
tran (\sa_snapshot[0][31] , \sa_snapshot[0].r.part0[31] );
tran (\sa_snapshot[0][31] , \sa_snapshot[0].f.lower[31] );
tran (\sa_snapshot[0][30] , \sa_snapshot[0].r.part0[30] );
tran (\sa_snapshot[0][30] , \sa_snapshot[0].f.lower[30] );
tran (\sa_snapshot[0][29] , \sa_snapshot[0].r.part0[29] );
tran (\sa_snapshot[0][29] , \sa_snapshot[0].f.lower[29] );
tran (\sa_snapshot[0][28] , \sa_snapshot[0].r.part0[28] );
tran (\sa_snapshot[0][28] , \sa_snapshot[0].f.lower[28] );
tran (\sa_snapshot[0][27] , \sa_snapshot[0].r.part0[27] );
tran (\sa_snapshot[0][27] , \sa_snapshot[0].f.lower[27] );
tran (\sa_snapshot[0][26] , \sa_snapshot[0].r.part0[26] );
tran (\sa_snapshot[0][26] , \sa_snapshot[0].f.lower[26] );
tran (\sa_snapshot[0][25] , \sa_snapshot[0].r.part0[25] );
tran (\sa_snapshot[0][25] , \sa_snapshot[0].f.lower[25] );
tran (\sa_snapshot[0][24] , \sa_snapshot[0].r.part0[24] );
tran (\sa_snapshot[0][24] , \sa_snapshot[0].f.lower[24] );
tran (\sa_snapshot[0][23] , \sa_snapshot[0].r.part0[23] );
tran (\sa_snapshot[0][23] , \sa_snapshot[0].f.lower[23] );
tran (\sa_snapshot[0][22] , \sa_snapshot[0].r.part0[22] );
tran (\sa_snapshot[0][22] , \sa_snapshot[0].f.lower[22] );
tran (\sa_snapshot[0][21] , \sa_snapshot[0].r.part0[21] );
tran (\sa_snapshot[0][21] , \sa_snapshot[0].f.lower[21] );
tran (\sa_snapshot[0][20] , \sa_snapshot[0].r.part0[20] );
tran (\sa_snapshot[0][20] , \sa_snapshot[0].f.lower[20] );
tran (\sa_snapshot[0][19] , \sa_snapshot[0].r.part0[19] );
tran (\sa_snapshot[0][19] , \sa_snapshot[0].f.lower[19] );
tran (\sa_snapshot[0][18] , \sa_snapshot[0].r.part0[18] );
tran (\sa_snapshot[0][18] , \sa_snapshot[0].f.lower[18] );
tran (\sa_snapshot[0][17] , \sa_snapshot[0].r.part0[17] );
tran (\sa_snapshot[0][17] , \sa_snapshot[0].f.lower[17] );
tran (\sa_snapshot[0][16] , \sa_snapshot[0].r.part0[16] );
tran (\sa_snapshot[0][16] , \sa_snapshot[0].f.lower[16] );
tran (\sa_snapshot[0][15] , \sa_snapshot[0].r.part0[15] );
tran (\sa_snapshot[0][15] , \sa_snapshot[0].f.lower[15] );
tran (\sa_snapshot[0][14] , \sa_snapshot[0].r.part0[14] );
tran (\sa_snapshot[0][14] , \sa_snapshot[0].f.lower[14] );
tran (\sa_snapshot[0][13] , \sa_snapshot[0].r.part0[13] );
tran (\sa_snapshot[0][13] , \sa_snapshot[0].f.lower[13] );
tran (\sa_snapshot[0][12] , \sa_snapshot[0].r.part0[12] );
tran (\sa_snapshot[0][12] , \sa_snapshot[0].f.lower[12] );
tran (\sa_snapshot[0][11] , \sa_snapshot[0].r.part0[11] );
tran (\sa_snapshot[0][11] , \sa_snapshot[0].f.lower[11] );
tran (\sa_snapshot[0][10] , \sa_snapshot[0].r.part0[10] );
tran (\sa_snapshot[0][10] , \sa_snapshot[0].f.lower[10] );
tran (\sa_snapshot[0][9] , \sa_snapshot[0].r.part0[9] );
tran (\sa_snapshot[0][9] , \sa_snapshot[0].f.lower[9] );
tran (\sa_snapshot[0][8] , \sa_snapshot[0].r.part0[8] );
tran (\sa_snapshot[0][8] , \sa_snapshot[0].f.lower[8] );
tran (\sa_snapshot[0][7] , \sa_snapshot[0].r.part0[7] );
tran (\sa_snapshot[0][7] , \sa_snapshot[0].f.lower[7] );
tran (\sa_snapshot[0][6] , \sa_snapshot[0].r.part0[6] );
tran (\sa_snapshot[0][6] , \sa_snapshot[0].f.lower[6] );
tran (\sa_snapshot[0][5] , \sa_snapshot[0].r.part0[5] );
tran (\sa_snapshot[0][5] , \sa_snapshot[0].f.lower[5] );
tran (\sa_snapshot[0][4] , \sa_snapshot[0].r.part0[4] );
tran (\sa_snapshot[0][4] , \sa_snapshot[0].f.lower[4] );
tran (\sa_snapshot[0][3] , \sa_snapshot[0].r.part0[3] );
tran (\sa_snapshot[0][3] , \sa_snapshot[0].f.lower[3] );
tran (\sa_snapshot[0][2] , \sa_snapshot[0].r.part0[2] );
tran (\sa_snapshot[0][2] , \sa_snapshot[0].f.lower[2] );
tran (\sa_snapshot[0][1] , \sa_snapshot[0].r.part0[1] );
tran (\sa_snapshot[0][1] , \sa_snapshot[0].f.lower[1] );
tran (\sa_snapshot[0][0] , \sa_snapshot[0].r.part0[0] );
tran (\sa_snapshot[0][0] , \sa_snapshot[0].f.lower[0] );
tran (\sa_count[31][63] , \sa_count[31].r.part1[31] );
tran (\sa_count[31][63] , \sa_count[31].f.unused[13] );
tran (\sa_count[31][62] , \sa_count[31].r.part1[30] );
tran (\sa_count[31][62] , \sa_count[31].f.unused[12] );
tran (\sa_count[31][61] , \sa_count[31].r.part1[29] );
tran (\sa_count[31][61] , \sa_count[31].f.unused[11] );
tran (\sa_count[31][60] , \sa_count[31].r.part1[28] );
tran (\sa_count[31][60] , \sa_count[31].f.unused[10] );
tran (\sa_count[31][59] , \sa_count[31].r.part1[27] );
tran (\sa_count[31][59] , \sa_count[31].f.unused[9] );
tran (\sa_count[31][58] , \sa_count[31].r.part1[26] );
tran (\sa_count[31][58] , \sa_count[31].f.unused[8] );
tran (\sa_count[31][57] , \sa_count[31].r.part1[25] );
tran (\sa_count[31][57] , \sa_count[31].f.unused[7] );
tran (\sa_count[31][56] , \sa_count[31].r.part1[24] );
tran (\sa_count[31][56] , \sa_count[31].f.unused[6] );
tran (\sa_count[31][55] , \sa_count[31].r.part1[23] );
tran (\sa_count[31][55] , \sa_count[31].f.unused[5] );
tran (\sa_count[31][54] , \sa_count[31].r.part1[22] );
tran (\sa_count[31][54] , \sa_count[31].f.unused[4] );
tran (\sa_count[31][53] , \sa_count[31].r.part1[21] );
tran (\sa_count[31][53] , \sa_count[31].f.unused[3] );
tran (\sa_count[31][52] , \sa_count[31].r.part1[20] );
tran (\sa_count[31][52] , \sa_count[31].f.unused[2] );
tran (\sa_count[31][51] , \sa_count[31].r.part1[19] );
tran (\sa_count[31][51] , \sa_count[31].f.unused[1] );
tran (\sa_count[31][50] , \sa_count[31].r.part1[18] );
tran (\sa_count[31][50] , \sa_count[31].f.unused[0] );
tran (\sa_count[31][49] , \sa_count[31].r.part1[17] );
tran (\sa_count[31][49] , \sa_count[31].f.upper[17] );
tran (\sa_count[31][48] , \sa_count[31].r.part1[16] );
tran (\sa_count[31][48] , \sa_count[31].f.upper[16] );
tran (\sa_count[31][47] , \sa_count[31].r.part1[15] );
tran (\sa_count[31][47] , \sa_count[31].f.upper[15] );
tran (\sa_count[31][46] , \sa_count[31].r.part1[14] );
tran (\sa_count[31][46] , \sa_count[31].f.upper[14] );
tran (\sa_count[31][45] , \sa_count[31].r.part1[13] );
tran (\sa_count[31][45] , \sa_count[31].f.upper[13] );
tran (\sa_count[31][44] , \sa_count[31].r.part1[12] );
tran (\sa_count[31][44] , \sa_count[31].f.upper[12] );
tran (\sa_count[31][43] , \sa_count[31].r.part1[11] );
tran (\sa_count[31][43] , \sa_count[31].f.upper[11] );
tran (\sa_count[31][42] , \sa_count[31].r.part1[10] );
tran (\sa_count[31][42] , \sa_count[31].f.upper[10] );
tran (\sa_count[31][41] , \sa_count[31].r.part1[9] );
tran (\sa_count[31][41] , \sa_count[31].f.upper[9] );
tran (\sa_count[31][40] , \sa_count[31].r.part1[8] );
tran (\sa_count[31][40] , \sa_count[31].f.upper[8] );
tran (\sa_count[31][39] , \sa_count[31].r.part1[7] );
tran (\sa_count[31][39] , \sa_count[31].f.upper[7] );
tran (\sa_count[31][38] , \sa_count[31].r.part1[6] );
tran (\sa_count[31][38] , \sa_count[31].f.upper[6] );
tran (\sa_count[31][37] , \sa_count[31].r.part1[5] );
tran (\sa_count[31][37] , \sa_count[31].f.upper[5] );
tran (\sa_count[31][36] , \sa_count[31].r.part1[4] );
tran (\sa_count[31][36] , \sa_count[31].f.upper[4] );
tran (\sa_count[31][35] , \sa_count[31].r.part1[3] );
tran (\sa_count[31][35] , \sa_count[31].f.upper[3] );
tran (\sa_count[31][34] , \sa_count[31].r.part1[2] );
tran (\sa_count[31][34] , \sa_count[31].f.upper[2] );
tran (\sa_count[31][33] , \sa_count[31].r.part1[1] );
tran (\sa_count[31][33] , \sa_count[31].f.upper[1] );
tran (\sa_count[31][32] , \sa_count[31].r.part1[0] );
tran (\sa_count[31][32] , \sa_count[31].f.upper[0] );
tran (\sa_count[31][31] , \sa_count[31].r.part0[31] );
tran (\sa_count[31][31] , \sa_count[31].f.lower[31] );
tran (\sa_count[31][30] , \sa_count[31].r.part0[30] );
tran (\sa_count[31][30] , \sa_count[31].f.lower[30] );
tran (\sa_count[31][29] , \sa_count[31].r.part0[29] );
tran (\sa_count[31][29] , \sa_count[31].f.lower[29] );
tran (\sa_count[31][28] , \sa_count[31].r.part0[28] );
tran (\sa_count[31][28] , \sa_count[31].f.lower[28] );
tran (\sa_count[31][27] , \sa_count[31].r.part0[27] );
tran (\sa_count[31][27] , \sa_count[31].f.lower[27] );
tran (\sa_count[31][26] , \sa_count[31].r.part0[26] );
tran (\sa_count[31][26] , \sa_count[31].f.lower[26] );
tran (\sa_count[31][25] , \sa_count[31].r.part0[25] );
tran (\sa_count[31][25] , \sa_count[31].f.lower[25] );
tran (\sa_count[31][24] , \sa_count[31].r.part0[24] );
tran (\sa_count[31][24] , \sa_count[31].f.lower[24] );
tran (\sa_count[31][23] , \sa_count[31].r.part0[23] );
tran (\sa_count[31][23] , \sa_count[31].f.lower[23] );
tran (\sa_count[31][22] , \sa_count[31].r.part0[22] );
tran (\sa_count[31][22] , \sa_count[31].f.lower[22] );
tran (\sa_count[31][21] , \sa_count[31].r.part0[21] );
tran (\sa_count[31][21] , \sa_count[31].f.lower[21] );
tran (\sa_count[31][20] , \sa_count[31].r.part0[20] );
tran (\sa_count[31][20] , \sa_count[31].f.lower[20] );
tran (\sa_count[31][19] , \sa_count[31].r.part0[19] );
tran (\sa_count[31][19] , \sa_count[31].f.lower[19] );
tran (\sa_count[31][18] , \sa_count[31].r.part0[18] );
tran (\sa_count[31][18] , \sa_count[31].f.lower[18] );
tran (\sa_count[31][17] , \sa_count[31].r.part0[17] );
tran (\sa_count[31][17] , \sa_count[31].f.lower[17] );
tran (\sa_count[31][16] , \sa_count[31].r.part0[16] );
tran (\sa_count[31][16] , \sa_count[31].f.lower[16] );
tran (\sa_count[31][15] , \sa_count[31].r.part0[15] );
tran (\sa_count[31][15] , \sa_count[31].f.lower[15] );
tran (\sa_count[31][14] , \sa_count[31].r.part0[14] );
tran (\sa_count[31][14] , \sa_count[31].f.lower[14] );
tran (\sa_count[31][13] , \sa_count[31].r.part0[13] );
tran (\sa_count[31][13] , \sa_count[31].f.lower[13] );
tran (\sa_count[31][12] , \sa_count[31].r.part0[12] );
tran (\sa_count[31][12] , \sa_count[31].f.lower[12] );
tran (\sa_count[31][11] , \sa_count[31].r.part0[11] );
tran (\sa_count[31][11] , \sa_count[31].f.lower[11] );
tran (\sa_count[31][10] , \sa_count[31].r.part0[10] );
tran (\sa_count[31][10] , \sa_count[31].f.lower[10] );
tran (\sa_count[31][9] , \sa_count[31].r.part0[9] );
tran (\sa_count[31][9] , \sa_count[31].f.lower[9] );
tran (\sa_count[31][8] , \sa_count[31].r.part0[8] );
tran (\sa_count[31][8] , \sa_count[31].f.lower[8] );
tran (\sa_count[31][7] , \sa_count[31].r.part0[7] );
tran (\sa_count[31][7] , \sa_count[31].f.lower[7] );
tran (\sa_count[31][6] , \sa_count[31].r.part0[6] );
tran (\sa_count[31][6] , \sa_count[31].f.lower[6] );
tran (\sa_count[31][5] , \sa_count[31].r.part0[5] );
tran (\sa_count[31][5] , \sa_count[31].f.lower[5] );
tran (\sa_count[31][4] , \sa_count[31].r.part0[4] );
tran (\sa_count[31][4] , \sa_count[31].f.lower[4] );
tran (\sa_count[31][3] , \sa_count[31].r.part0[3] );
tran (\sa_count[31][3] , \sa_count[31].f.lower[3] );
tran (\sa_count[31][2] , \sa_count[31].r.part0[2] );
tran (\sa_count[31][2] , \sa_count[31].f.lower[2] );
tran (\sa_count[31][1] , \sa_count[31].r.part0[1] );
tran (\sa_count[31][1] , \sa_count[31].f.lower[1] );
tran (\sa_count[31][0] , \sa_count[31].r.part0[0] );
tran (\sa_count[31][0] , \sa_count[31].f.lower[0] );
tran (\sa_count[30][63] , \sa_count[30].r.part1[31] );
tran (\sa_count[30][63] , \sa_count[30].f.unused[13] );
tran (\sa_count[30][62] , \sa_count[30].r.part1[30] );
tran (\sa_count[30][62] , \sa_count[30].f.unused[12] );
tran (\sa_count[30][61] , \sa_count[30].r.part1[29] );
tran (\sa_count[30][61] , \sa_count[30].f.unused[11] );
tran (\sa_count[30][60] , \sa_count[30].r.part1[28] );
tran (\sa_count[30][60] , \sa_count[30].f.unused[10] );
tran (\sa_count[30][59] , \sa_count[30].r.part1[27] );
tran (\sa_count[30][59] , \sa_count[30].f.unused[9] );
tran (\sa_count[30][58] , \sa_count[30].r.part1[26] );
tran (\sa_count[30][58] , \sa_count[30].f.unused[8] );
tran (\sa_count[30][57] , \sa_count[30].r.part1[25] );
tran (\sa_count[30][57] , \sa_count[30].f.unused[7] );
tran (\sa_count[30][56] , \sa_count[30].r.part1[24] );
tran (\sa_count[30][56] , \sa_count[30].f.unused[6] );
tran (\sa_count[30][55] , \sa_count[30].r.part1[23] );
tran (\sa_count[30][55] , \sa_count[30].f.unused[5] );
tran (\sa_count[30][54] , \sa_count[30].r.part1[22] );
tran (\sa_count[30][54] , \sa_count[30].f.unused[4] );
tran (\sa_count[30][53] , \sa_count[30].r.part1[21] );
tran (\sa_count[30][53] , \sa_count[30].f.unused[3] );
tran (\sa_count[30][52] , \sa_count[30].r.part1[20] );
tran (\sa_count[30][52] , \sa_count[30].f.unused[2] );
tran (\sa_count[30][51] , \sa_count[30].r.part1[19] );
tran (\sa_count[30][51] , \sa_count[30].f.unused[1] );
tran (\sa_count[30][50] , \sa_count[30].r.part1[18] );
tran (\sa_count[30][50] , \sa_count[30].f.unused[0] );
tran (\sa_count[30][49] , \sa_count[30].r.part1[17] );
tran (\sa_count[30][49] , \sa_count[30].f.upper[17] );
tran (\sa_count[30][48] , \sa_count[30].r.part1[16] );
tran (\sa_count[30][48] , \sa_count[30].f.upper[16] );
tran (\sa_count[30][47] , \sa_count[30].r.part1[15] );
tran (\sa_count[30][47] , \sa_count[30].f.upper[15] );
tran (\sa_count[30][46] , \sa_count[30].r.part1[14] );
tran (\sa_count[30][46] , \sa_count[30].f.upper[14] );
tran (\sa_count[30][45] , \sa_count[30].r.part1[13] );
tran (\sa_count[30][45] , \sa_count[30].f.upper[13] );
tran (\sa_count[30][44] , \sa_count[30].r.part1[12] );
tran (\sa_count[30][44] , \sa_count[30].f.upper[12] );
tran (\sa_count[30][43] , \sa_count[30].r.part1[11] );
tran (\sa_count[30][43] , \sa_count[30].f.upper[11] );
tran (\sa_count[30][42] , \sa_count[30].r.part1[10] );
tran (\sa_count[30][42] , \sa_count[30].f.upper[10] );
tran (\sa_count[30][41] , \sa_count[30].r.part1[9] );
tran (\sa_count[30][41] , \sa_count[30].f.upper[9] );
tran (\sa_count[30][40] , \sa_count[30].r.part1[8] );
tran (\sa_count[30][40] , \sa_count[30].f.upper[8] );
tran (\sa_count[30][39] , \sa_count[30].r.part1[7] );
tran (\sa_count[30][39] , \sa_count[30].f.upper[7] );
tran (\sa_count[30][38] , \sa_count[30].r.part1[6] );
tran (\sa_count[30][38] , \sa_count[30].f.upper[6] );
tran (\sa_count[30][37] , \sa_count[30].r.part1[5] );
tran (\sa_count[30][37] , \sa_count[30].f.upper[5] );
tran (\sa_count[30][36] , \sa_count[30].r.part1[4] );
tran (\sa_count[30][36] , \sa_count[30].f.upper[4] );
tran (\sa_count[30][35] , \sa_count[30].r.part1[3] );
tran (\sa_count[30][35] , \sa_count[30].f.upper[3] );
tran (\sa_count[30][34] , \sa_count[30].r.part1[2] );
tran (\sa_count[30][34] , \sa_count[30].f.upper[2] );
tran (\sa_count[30][33] , \sa_count[30].r.part1[1] );
tran (\sa_count[30][33] , \sa_count[30].f.upper[1] );
tran (\sa_count[30][32] , \sa_count[30].r.part1[0] );
tran (\sa_count[30][32] , \sa_count[30].f.upper[0] );
tran (\sa_count[30][31] , \sa_count[30].r.part0[31] );
tran (\sa_count[30][31] , \sa_count[30].f.lower[31] );
tran (\sa_count[30][30] , \sa_count[30].r.part0[30] );
tran (\sa_count[30][30] , \sa_count[30].f.lower[30] );
tran (\sa_count[30][29] , \sa_count[30].r.part0[29] );
tran (\sa_count[30][29] , \sa_count[30].f.lower[29] );
tran (\sa_count[30][28] , \sa_count[30].r.part0[28] );
tran (\sa_count[30][28] , \sa_count[30].f.lower[28] );
tran (\sa_count[30][27] , \sa_count[30].r.part0[27] );
tran (\sa_count[30][27] , \sa_count[30].f.lower[27] );
tran (\sa_count[30][26] , \sa_count[30].r.part0[26] );
tran (\sa_count[30][26] , \sa_count[30].f.lower[26] );
tran (\sa_count[30][25] , \sa_count[30].r.part0[25] );
tran (\sa_count[30][25] , \sa_count[30].f.lower[25] );
tran (\sa_count[30][24] , \sa_count[30].r.part0[24] );
tran (\sa_count[30][24] , \sa_count[30].f.lower[24] );
tran (\sa_count[30][23] , \sa_count[30].r.part0[23] );
tran (\sa_count[30][23] , \sa_count[30].f.lower[23] );
tran (\sa_count[30][22] , \sa_count[30].r.part0[22] );
tran (\sa_count[30][22] , \sa_count[30].f.lower[22] );
tran (\sa_count[30][21] , \sa_count[30].r.part0[21] );
tran (\sa_count[30][21] , \sa_count[30].f.lower[21] );
tran (\sa_count[30][20] , \sa_count[30].r.part0[20] );
tran (\sa_count[30][20] , \sa_count[30].f.lower[20] );
tran (\sa_count[30][19] , \sa_count[30].r.part0[19] );
tran (\sa_count[30][19] , \sa_count[30].f.lower[19] );
tran (\sa_count[30][18] , \sa_count[30].r.part0[18] );
tran (\sa_count[30][18] , \sa_count[30].f.lower[18] );
tran (\sa_count[30][17] , \sa_count[30].r.part0[17] );
tran (\sa_count[30][17] , \sa_count[30].f.lower[17] );
tran (\sa_count[30][16] , \sa_count[30].r.part0[16] );
tran (\sa_count[30][16] , \sa_count[30].f.lower[16] );
tran (\sa_count[30][15] , \sa_count[30].r.part0[15] );
tran (\sa_count[30][15] , \sa_count[30].f.lower[15] );
tran (\sa_count[30][14] , \sa_count[30].r.part0[14] );
tran (\sa_count[30][14] , \sa_count[30].f.lower[14] );
tran (\sa_count[30][13] , \sa_count[30].r.part0[13] );
tran (\sa_count[30][13] , \sa_count[30].f.lower[13] );
tran (\sa_count[30][12] , \sa_count[30].r.part0[12] );
tran (\sa_count[30][12] , \sa_count[30].f.lower[12] );
tran (\sa_count[30][11] , \sa_count[30].r.part0[11] );
tran (\sa_count[30][11] , \sa_count[30].f.lower[11] );
tran (\sa_count[30][10] , \sa_count[30].r.part0[10] );
tran (\sa_count[30][10] , \sa_count[30].f.lower[10] );
tran (\sa_count[30][9] , \sa_count[30].r.part0[9] );
tran (\sa_count[30][9] , \sa_count[30].f.lower[9] );
tran (\sa_count[30][8] , \sa_count[30].r.part0[8] );
tran (\sa_count[30][8] , \sa_count[30].f.lower[8] );
tran (\sa_count[30][7] , \sa_count[30].r.part0[7] );
tran (\sa_count[30][7] , \sa_count[30].f.lower[7] );
tran (\sa_count[30][6] , \sa_count[30].r.part0[6] );
tran (\sa_count[30][6] , \sa_count[30].f.lower[6] );
tran (\sa_count[30][5] , \sa_count[30].r.part0[5] );
tran (\sa_count[30][5] , \sa_count[30].f.lower[5] );
tran (\sa_count[30][4] , \sa_count[30].r.part0[4] );
tran (\sa_count[30][4] , \sa_count[30].f.lower[4] );
tran (\sa_count[30][3] , \sa_count[30].r.part0[3] );
tran (\sa_count[30][3] , \sa_count[30].f.lower[3] );
tran (\sa_count[30][2] , \sa_count[30].r.part0[2] );
tran (\sa_count[30][2] , \sa_count[30].f.lower[2] );
tran (\sa_count[30][1] , \sa_count[30].r.part0[1] );
tran (\sa_count[30][1] , \sa_count[30].f.lower[1] );
tran (\sa_count[30][0] , \sa_count[30].r.part0[0] );
tran (\sa_count[30][0] , \sa_count[30].f.lower[0] );
tran (\sa_count[29][63] , \sa_count[29].r.part1[31] );
tran (\sa_count[29][63] , \sa_count[29].f.unused[13] );
tran (\sa_count[29][62] , \sa_count[29].r.part1[30] );
tran (\sa_count[29][62] , \sa_count[29].f.unused[12] );
tran (\sa_count[29][61] , \sa_count[29].r.part1[29] );
tran (\sa_count[29][61] , \sa_count[29].f.unused[11] );
tran (\sa_count[29][60] , \sa_count[29].r.part1[28] );
tran (\sa_count[29][60] , \sa_count[29].f.unused[10] );
tran (\sa_count[29][59] , \sa_count[29].r.part1[27] );
tran (\sa_count[29][59] , \sa_count[29].f.unused[9] );
tran (\sa_count[29][58] , \sa_count[29].r.part1[26] );
tran (\sa_count[29][58] , \sa_count[29].f.unused[8] );
tran (\sa_count[29][57] , \sa_count[29].r.part1[25] );
tran (\sa_count[29][57] , \sa_count[29].f.unused[7] );
tran (\sa_count[29][56] , \sa_count[29].r.part1[24] );
tran (\sa_count[29][56] , \sa_count[29].f.unused[6] );
tran (\sa_count[29][55] , \sa_count[29].r.part1[23] );
tran (\sa_count[29][55] , \sa_count[29].f.unused[5] );
tran (\sa_count[29][54] , \sa_count[29].r.part1[22] );
tran (\sa_count[29][54] , \sa_count[29].f.unused[4] );
tran (\sa_count[29][53] , \sa_count[29].r.part1[21] );
tran (\sa_count[29][53] , \sa_count[29].f.unused[3] );
tran (\sa_count[29][52] , \sa_count[29].r.part1[20] );
tran (\sa_count[29][52] , \sa_count[29].f.unused[2] );
tran (\sa_count[29][51] , \sa_count[29].r.part1[19] );
tran (\sa_count[29][51] , \sa_count[29].f.unused[1] );
tran (\sa_count[29][50] , \sa_count[29].r.part1[18] );
tran (\sa_count[29][50] , \sa_count[29].f.unused[0] );
tran (\sa_count[29][49] , \sa_count[29].r.part1[17] );
tran (\sa_count[29][49] , \sa_count[29].f.upper[17] );
tran (\sa_count[29][48] , \sa_count[29].r.part1[16] );
tran (\sa_count[29][48] , \sa_count[29].f.upper[16] );
tran (\sa_count[29][47] , \sa_count[29].r.part1[15] );
tran (\sa_count[29][47] , \sa_count[29].f.upper[15] );
tran (\sa_count[29][46] , \sa_count[29].r.part1[14] );
tran (\sa_count[29][46] , \sa_count[29].f.upper[14] );
tran (\sa_count[29][45] , \sa_count[29].r.part1[13] );
tran (\sa_count[29][45] , \sa_count[29].f.upper[13] );
tran (\sa_count[29][44] , \sa_count[29].r.part1[12] );
tran (\sa_count[29][44] , \sa_count[29].f.upper[12] );
tran (\sa_count[29][43] , \sa_count[29].r.part1[11] );
tran (\sa_count[29][43] , \sa_count[29].f.upper[11] );
tran (\sa_count[29][42] , \sa_count[29].r.part1[10] );
tran (\sa_count[29][42] , \sa_count[29].f.upper[10] );
tran (\sa_count[29][41] , \sa_count[29].r.part1[9] );
tran (\sa_count[29][41] , \sa_count[29].f.upper[9] );
tran (\sa_count[29][40] , \sa_count[29].r.part1[8] );
tran (\sa_count[29][40] , \sa_count[29].f.upper[8] );
tran (\sa_count[29][39] , \sa_count[29].r.part1[7] );
tran (\sa_count[29][39] , \sa_count[29].f.upper[7] );
tran (\sa_count[29][38] , \sa_count[29].r.part1[6] );
tran (\sa_count[29][38] , \sa_count[29].f.upper[6] );
tran (\sa_count[29][37] , \sa_count[29].r.part1[5] );
tran (\sa_count[29][37] , \sa_count[29].f.upper[5] );
tran (\sa_count[29][36] , \sa_count[29].r.part1[4] );
tran (\sa_count[29][36] , \sa_count[29].f.upper[4] );
tran (\sa_count[29][35] , \sa_count[29].r.part1[3] );
tran (\sa_count[29][35] , \sa_count[29].f.upper[3] );
tran (\sa_count[29][34] , \sa_count[29].r.part1[2] );
tran (\sa_count[29][34] , \sa_count[29].f.upper[2] );
tran (\sa_count[29][33] , \sa_count[29].r.part1[1] );
tran (\sa_count[29][33] , \sa_count[29].f.upper[1] );
tran (\sa_count[29][32] , \sa_count[29].r.part1[0] );
tran (\sa_count[29][32] , \sa_count[29].f.upper[0] );
tran (\sa_count[29][31] , \sa_count[29].r.part0[31] );
tran (\sa_count[29][31] , \sa_count[29].f.lower[31] );
tran (\sa_count[29][30] , \sa_count[29].r.part0[30] );
tran (\sa_count[29][30] , \sa_count[29].f.lower[30] );
tran (\sa_count[29][29] , \sa_count[29].r.part0[29] );
tran (\sa_count[29][29] , \sa_count[29].f.lower[29] );
tran (\sa_count[29][28] , \sa_count[29].r.part0[28] );
tran (\sa_count[29][28] , \sa_count[29].f.lower[28] );
tran (\sa_count[29][27] , \sa_count[29].r.part0[27] );
tran (\sa_count[29][27] , \sa_count[29].f.lower[27] );
tran (\sa_count[29][26] , \sa_count[29].r.part0[26] );
tran (\sa_count[29][26] , \sa_count[29].f.lower[26] );
tran (\sa_count[29][25] , \sa_count[29].r.part0[25] );
tran (\sa_count[29][25] , \sa_count[29].f.lower[25] );
tran (\sa_count[29][24] , \sa_count[29].r.part0[24] );
tran (\sa_count[29][24] , \sa_count[29].f.lower[24] );
tran (\sa_count[29][23] , \sa_count[29].r.part0[23] );
tran (\sa_count[29][23] , \sa_count[29].f.lower[23] );
tran (\sa_count[29][22] , \sa_count[29].r.part0[22] );
tran (\sa_count[29][22] , \sa_count[29].f.lower[22] );
tran (\sa_count[29][21] , \sa_count[29].r.part0[21] );
tran (\sa_count[29][21] , \sa_count[29].f.lower[21] );
tran (\sa_count[29][20] , \sa_count[29].r.part0[20] );
tran (\sa_count[29][20] , \sa_count[29].f.lower[20] );
tran (\sa_count[29][19] , \sa_count[29].r.part0[19] );
tran (\sa_count[29][19] , \sa_count[29].f.lower[19] );
tran (\sa_count[29][18] , \sa_count[29].r.part0[18] );
tran (\sa_count[29][18] , \sa_count[29].f.lower[18] );
tran (\sa_count[29][17] , \sa_count[29].r.part0[17] );
tran (\sa_count[29][17] , \sa_count[29].f.lower[17] );
tran (\sa_count[29][16] , \sa_count[29].r.part0[16] );
tran (\sa_count[29][16] , \sa_count[29].f.lower[16] );
tran (\sa_count[29][15] , \sa_count[29].r.part0[15] );
tran (\sa_count[29][15] , \sa_count[29].f.lower[15] );
tran (\sa_count[29][14] , \sa_count[29].r.part0[14] );
tran (\sa_count[29][14] , \sa_count[29].f.lower[14] );
tran (\sa_count[29][13] , \sa_count[29].r.part0[13] );
tran (\sa_count[29][13] , \sa_count[29].f.lower[13] );
tran (\sa_count[29][12] , \sa_count[29].r.part0[12] );
tran (\sa_count[29][12] , \sa_count[29].f.lower[12] );
tran (\sa_count[29][11] , \sa_count[29].r.part0[11] );
tran (\sa_count[29][11] , \sa_count[29].f.lower[11] );
tran (\sa_count[29][10] , \sa_count[29].r.part0[10] );
tran (\sa_count[29][10] , \sa_count[29].f.lower[10] );
tran (\sa_count[29][9] , \sa_count[29].r.part0[9] );
tran (\sa_count[29][9] , \sa_count[29].f.lower[9] );
tran (\sa_count[29][8] , \sa_count[29].r.part0[8] );
tran (\sa_count[29][8] , \sa_count[29].f.lower[8] );
tran (\sa_count[29][7] , \sa_count[29].r.part0[7] );
tran (\sa_count[29][7] , \sa_count[29].f.lower[7] );
tran (\sa_count[29][6] , \sa_count[29].r.part0[6] );
tran (\sa_count[29][6] , \sa_count[29].f.lower[6] );
tran (\sa_count[29][5] , \sa_count[29].r.part0[5] );
tran (\sa_count[29][5] , \sa_count[29].f.lower[5] );
tran (\sa_count[29][4] , \sa_count[29].r.part0[4] );
tran (\sa_count[29][4] , \sa_count[29].f.lower[4] );
tran (\sa_count[29][3] , \sa_count[29].r.part0[3] );
tran (\sa_count[29][3] , \sa_count[29].f.lower[3] );
tran (\sa_count[29][2] , \sa_count[29].r.part0[2] );
tran (\sa_count[29][2] , \sa_count[29].f.lower[2] );
tran (\sa_count[29][1] , \sa_count[29].r.part0[1] );
tran (\sa_count[29][1] , \sa_count[29].f.lower[1] );
tran (\sa_count[29][0] , \sa_count[29].r.part0[0] );
tran (\sa_count[29][0] , \sa_count[29].f.lower[0] );
tran (\sa_count[28][63] , \sa_count[28].r.part1[31] );
tran (\sa_count[28][63] , \sa_count[28].f.unused[13] );
tran (\sa_count[28][62] , \sa_count[28].r.part1[30] );
tran (\sa_count[28][62] , \sa_count[28].f.unused[12] );
tran (\sa_count[28][61] , \sa_count[28].r.part1[29] );
tran (\sa_count[28][61] , \sa_count[28].f.unused[11] );
tran (\sa_count[28][60] , \sa_count[28].r.part1[28] );
tran (\sa_count[28][60] , \sa_count[28].f.unused[10] );
tran (\sa_count[28][59] , \sa_count[28].r.part1[27] );
tran (\sa_count[28][59] , \sa_count[28].f.unused[9] );
tran (\sa_count[28][58] , \sa_count[28].r.part1[26] );
tran (\sa_count[28][58] , \sa_count[28].f.unused[8] );
tran (\sa_count[28][57] , \sa_count[28].r.part1[25] );
tran (\sa_count[28][57] , \sa_count[28].f.unused[7] );
tran (\sa_count[28][56] , \sa_count[28].r.part1[24] );
tran (\sa_count[28][56] , \sa_count[28].f.unused[6] );
tran (\sa_count[28][55] , \sa_count[28].r.part1[23] );
tran (\sa_count[28][55] , \sa_count[28].f.unused[5] );
tran (\sa_count[28][54] , \sa_count[28].r.part1[22] );
tran (\sa_count[28][54] , \sa_count[28].f.unused[4] );
tran (\sa_count[28][53] , \sa_count[28].r.part1[21] );
tran (\sa_count[28][53] , \sa_count[28].f.unused[3] );
tran (\sa_count[28][52] , \sa_count[28].r.part1[20] );
tran (\sa_count[28][52] , \sa_count[28].f.unused[2] );
tran (\sa_count[28][51] , \sa_count[28].r.part1[19] );
tran (\sa_count[28][51] , \sa_count[28].f.unused[1] );
tran (\sa_count[28][50] , \sa_count[28].r.part1[18] );
tran (\sa_count[28][50] , \sa_count[28].f.unused[0] );
tran (\sa_count[28][49] , \sa_count[28].r.part1[17] );
tran (\sa_count[28][49] , \sa_count[28].f.upper[17] );
tran (\sa_count[28][48] , \sa_count[28].r.part1[16] );
tran (\sa_count[28][48] , \sa_count[28].f.upper[16] );
tran (\sa_count[28][47] , \sa_count[28].r.part1[15] );
tran (\sa_count[28][47] , \sa_count[28].f.upper[15] );
tran (\sa_count[28][46] , \sa_count[28].r.part1[14] );
tran (\sa_count[28][46] , \sa_count[28].f.upper[14] );
tran (\sa_count[28][45] , \sa_count[28].r.part1[13] );
tran (\sa_count[28][45] , \sa_count[28].f.upper[13] );
tran (\sa_count[28][44] , \sa_count[28].r.part1[12] );
tran (\sa_count[28][44] , \sa_count[28].f.upper[12] );
tran (\sa_count[28][43] , \sa_count[28].r.part1[11] );
tran (\sa_count[28][43] , \sa_count[28].f.upper[11] );
tran (\sa_count[28][42] , \sa_count[28].r.part1[10] );
tran (\sa_count[28][42] , \sa_count[28].f.upper[10] );
tran (\sa_count[28][41] , \sa_count[28].r.part1[9] );
tran (\sa_count[28][41] , \sa_count[28].f.upper[9] );
tran (\sa_count[28][40] , \sa_count[28].r.part1[8] );
tran (\sa_count[28][40] , \sa_count[28].f.upper[8] );
tran (\sa_count[28][39] , \sa_count[28].r.part1[7] );
tran (\sa_count[28][39] , \sa_count[28].f.upper[7] );
tran (\sa_count[28][38] , \sa_count[28].r.part1[6] );
tran (\sa_count[28][38] , \sa_count[28].f.upper[6] );
tran (\sa_count[28][37] , \sa_count[28].r.part1[5] );
tran (\sa_count[28][37] , \sa_count[28].f.upper[5] );
tran (\sa_count[28][36] , \sa_count[28].r.part1[4] );
tran (\sa_count[28][36] , \sa_count[28].f.upper[4] );
tran (\sa_count[28][35] , \sa_count[28].r.part1[3] );
tran (\sa_count[28][35] , \sa_count[28].f.upper[3] );
tran (\sa_count[28][34] , \sa_count[28].r.part1[2] );
tran (\sa_count[28][34] , \sa_count[28].f.upper[2] );
tran (\sa_count[28][33] , \sa_count[28].r.part1[1] );
tran (\sa_count[28][33] , \sa_count[28].f.upper[1] );
tran (\sa_count[28][32] , \sa_count[28].r.part1[0] );
tran (\sa_count[28][32] , \sa_count[28].f.upper[0] );
tran (\sa_count[28][31] , \sa_count[28].r.part0[31] );
tran (\sa_count[28][31] , \sa_count[28].f.lower[31] );
tran (\sa_count[28][30] , \sa_count[28].r.part0[30] );
tran (\sa_count[28][30] , \sa_count[28].f.lower[30] );
tran (\sa_count[28][29] , \sa_count[28].r.part0[29] );
tran (\sa_count[28][29] , \sa_count[28].f.lower[29] );
tran (\sa_count[28][28] , \sa_count[28].r.part0[28] );
tran (\sa_count[28][28] , \sa_count[28].f.lower[28] );
tran (\sa_count[28][27] , \sa_count[28].r.part0[27] );
tran (\sa_count[28][27] , \sa_count[28].f.lower[27] );
tran (\sa_count[28][26] , \sa_count[28].r.part0[26] );
tran (\sa_count[28][26] , \sa_count[28].f.lower[26] );
tran (\sa_count[28][25] , \sa_count[28].r.part0[25] );
tran (\sa_count[28][25] , \sa_count[28].f.lower[25] );
tran (\sa_count[28][24] , \sa_count[28].r.part0[24] );
tran (\sa_count[28][24] , \sa_count[28].f.lower[24] );
tran (\sa_count[28][23] , \sa_count[28].r.part0[23] );
tran (\sa_count[28][23] , \sa_count[28].f.lower[23] );
tran (\sa_count[28][22] , \sa_count[28].r.part0[22] );
tran (\sa_count[28][22] , \sa_count[28].f.lower[22] );
tran (\sa_count[28][21] , \sa_count[28].r.part0[21] );
tran (\sa_count[28][21] , \sa_count[28].f.lower[21] );
tran (\sa_count[28][20] , \sa_count[28].r.part0[20] );
tran (\sa_count[28][20] , \sa_count[28].f.lower[20] );
tran (\sa_count[28][19] , \sa_count[28].r.part0[19] );
tran (\sa_count[28][19] , \sa_count[28].f.lower[19] );
tran (\sa_count[28][18] , \sa_count[28].r.part0[18] );
tran (\sa_count[28][18] , \sa_count[28].f.lower[18] );
tran (\sa_count[28][17] , \sa_count[28].r.part0[17] );
tran (\sa_count[28][17] , \sa_count[28].f.lower[17] );
tran (\sa_count[28][16] , \sa_count[28].r.part0[16] );
tran (\sa_count[28][16] , \sa_count[28].f.lower[16] );
tran (\sa_count[28][15] , \sa_count[28].r.part0[15] );
tran (\sa_count[28][15] , \sa_count[28].f.lower[15] );
tran (\sa_count[28][14] , \sa_count[28].r.part0[14] );
tran (\sa_count[28][14] , \sa_count[28].f.lower[14] );
tran (\sa_count[28][13] , \sa_count[28].r.part0[13] );
tran (\sa_count[28][13] , \sa_count[28].f.lower[13] );
tran (\sa_count[28][12] , \sa_count[28].r.part0[12] );
tran (\sa_count[28][12] , \sa_count[28].f.lower[12] );
tran (\sa_count[28][11] , \sa_count[28].r.part0[11] );
tran (\sa_count[28][11] , \sa_count[28].f.lower[11] );
tran (\sa_count[28][10] , \sa_count[28].r.part0[10] );
tran (\sa_count[28][10] , \sa_count[28].f.lower[10] );
tran (\sa_count[28][9] , \sa_count[28].r.part0[9] );
tran (\sa_count[28][9] , \sa_count[28].f.lower[9] );
tran (\sa_count[28][8] , \sa_count[28].r.part0[8] );
tran (\sa_count[28][8] , \sa_count[28].f.lower[8] );
tran (\sa_count[28][7] , \sa_count[28].r.part0[7] );
tran (\sa_count[28][7] , \sa_count[28].f.lower[7] );
tran (\sa_count[28][6] , \sa_count[28].r.part0[6] );
tran (\sa_count[28][6] , \sa_count[28].f.lower[6] );
tran (\sa_count[28][5] , \sa_count[28].r.part0[5] );
tran (\sa_count[28][5] , \sa_count[28].f.lower[5] );
tran (\sa_count[28][4] , \sa_count[28].r.part0[4] );
tran (\sa_count[28][4] , \sa_count[28].f.lower[4] );
tran (\sa_count[28][3] , \sa_count[28].r.part0[3] );
tran (\sa_count[28][3] , \sa_count[28].f.lower[3] );
tran (\sa_count[28][2] , \sa_count[28].r.part0[2] );
tran (\sa_count[28][2] , \sa_count[28].f.lower[2] );
tran (\sa_count[28][1] , \sa_count[28].r.part0[1] );
tran (\sa_count[28][1] , \sa_count[28].f.lower[1] );
tran (\sa_count[28][0] , \sa_count[28].r.part0[0] );
tran (\sa_count[28][0] , \sa_count[28].f.lower[0] );
tran (\sa_count[27][63] , \sa_count[27].r.part1[31] );
tran (\sa_count[27][63] , \sa_count[27].f.unused[13] );
tran (\sa_count[27][62] , \sa_count[27].r.part1[30] );
tran (\sa_count[27][62] , \sa_count[27].f.unused[12] );
tran (\sa_count[27][61] , \sa_count[27].r.part1[29] );
tran (\sa_count[27][61] , \sa_count[27].f.unused[11] );
tran (\sa_count[27][60] , \sa_count[27].r.part1[28] );
tran (\sa_count[27][60] , \sa_count[27].f.unused[10] );
tran (\sa_count[27][59] , \sa_count[27].r.part1[27] );
tran (\sa_count[27][59] , \sa_count[27].f.unused[9] );
tran (\sa_count[27][58] , \sa_count[27].r.part1[26] );
tran (\sa_count[27][58] , \sa_count[27].f.unused[8] );
tran (\sa_count[27][57] , \sa_count[27].r.part1[25] );
tran (\sa_count[27][57] , \sa_count[27].f.unused[7] );
tran (\sa_count[27][56] , \sa_count[27].r.part1[24] );
tran (\sa_count[27][56] , \sa_count[27].f.unused[6] );
tran (\sa_count[27][55] , \sa_count[27].r.part1[23] );
tran (\sa_count[27][55] , \sa_count[27].f.unused[5] );
tran (\sa_count[27][54] , \sa_count[27].r.part1[22] );
tran (\sa_count[27][54] , \sa_count[27].f.unused[4] );
tran (\sa_count[27][53] , \sa_count[27].r.part1[21] );
tran (\sa_count[27][53] , \sa_count[27].f.unused[3] );
tran (\sa_count[27][52] , \sa_count[27].r.part1[20] );
tran (\sa_count[27][52] , \sa_count[27].f.unused[2] );
tran (\sa_count[27][51] , \sa_count[27].r.part1[19] );
tran (\sa_count[27][51] , \sa_count[27].f.unused[1] );
tran (\sa_count[27][50] , \sa_count[27].r.part1[18] );
tran (\sa_count[27][50] , \sa_count[27].f.unused[0] );
tran (\sa_count[27][49] , \sa_count[27].r.part1[17] );
tran (\sa_count[27][49] , \sa_count[27].f.upper[17] );
tran (\sa_count[27][48] , \sa_count[27].r.part1[16] );
tran (\sa_count[27][48] , \sa_count[27].f.upper[16] );
tran (\sa_count[27][47] , \sa_count[27].r.part1[15] );
tran (\sa_count[27][47] , \sa_count[27].f.upper[15] );
tran (\sa_count[27][46] , \sa_count[27].r.part1[14] );
tran (\sa_count[27][46] , \sa_count[27].f.upper[14] );
tran (\sa_count[27][45] , \sa_count[27].r.part1[13] );
tran (\sa_count[27][45] , \sa_count[27].f.upper[13] );
tran (\sa_count[27][44] , \sa_count[27].r.part1[12] );
tran (\sa_count[27][44] , \sa_count[27].f.upper[12] );
tran (\sa_count[27][43] , \sa_count[27].r.part1[11] );
tran (\sa_count[27][43] , \sa_count[27].f.upper[11] );
tran (\sa_count[27][42] , \sa_count[27].r.part1[10] );
tran (\sa_count[27][42] , \sa_count[27].f.upper[10] );
tran (\sa_count[27][41] , \sa_count[27].r.part1[9] );
tran (\sa_count[27][41] , \sa_count[27].f.upper[9] );
tran (\sa_count[27][40] , \sa_count[27].r.part1[8] );
tran (\sa_count[27][40] , \sa_count[27].f.upper[8] );
tran (\sa_count[27][39] , \sa_count[27].r.part1[7] );
tran (\sa_count[27][39] , \sa_count[27].f.upper[7] );
tran (\sa_count[27][38] , \sa_count[27].r.part1[6] );
tran (\sa_count[27][38] , \sa_count[27].f.upper[6] );
tran (\sa_count[27][37] , \sa_count[27].r.part1[5] );
tran (\sa_count[27][37] , \sa_count[27].f.upper[5] );
tran (\sa_count[27][36] , \sa_count[27].r.part1[4] );
tran (\sa_count[27][36] , \sa_count[27].f.upper[4] );
tran (\sa_count[27][35] , \sa_count[27].r.part1[3] );
tran (\sa_count[27][35] , \sa_count[27].f.upper[3] );
tran (\sa_count[27][34] , \sa_count[27].r.part1[2] );
tran (\sa_count[27][34] , \sa_count[27].f.upper[2] );
tran (\sa_count[27][33] , \sa_count[27].r.part1[1] );
tran (\sa_count[27][33] , \sa_count[27].f.upper[1] );
tran (\sa_count[27][32] , \sa_count[27].r.part1[0] );
tran (\sa_count[27][32] , \sa_count[27].f.upper[0] );
tran (\sa_count[27][31] , \sa_count[27].r.part0[31] );
tran (\sa_count[27][31] , \sa_count[27].f.lower[31] );
tran (\sa_count[27][30] , \sa_count[27].r.part0[30] );
tran (\sa_count[27][30] , \sa_count[27].f.lower[30] );
tran (\sa_count[27][29] , \sa_count[27].r.part0[29] );
tran (\sa_count[27][29] , \sa_count[27].f.lower[29] );
tran (\sa_count[27][28] , \sa_count[27].r.part0[28] );
tran (\sa_count[27][28] , \sa_count[27].f.lower[28] );
tran (\sa_count[27][27] , \sa_count[27].r.part0[27] );
tran (\sa_count[27][27] , \sa_count[27].f.lower[27] );
tran (\sa_count[27][26] , \sa_count[27].r.part0[26] );
tran (\sa_count[27][26] , \sa_count[27].f.lower[26] );
tran (\sa_count[27][25] , \sa_count[27].r.part0[25] );
tran (\sa_count[27][25] , \sa_count[27].f.lower[25] );
tran (\sa_count[27][24] , \sa_count[27].r.part0[24] );
tran (\sa_count[27][24] , \sa_count[27].f.lower[24] );
tran (\sa_count[27][23] , \sa_count[27].r.part0[23] );
tran (\sa_count[27][23] , \sa_count[27].f.lower[23] );
tran (\sa_count[27][22] , \sa_count[27].r.part0[22] );
tran (\sa_count[27][22] , \sa_count[27].f.lower[22] );
tran (\sa_count[27][21] , \sa_count[27].r.part0[21] );
tran (\sa_count[27][21] , \sa_count[27].f.lower[21] );
tran (\sa_count[27][20] , \sa_count[27].r.part0[20] );
tran (\sa_count[27][20] , \sa_count[27].f.lower[20] );
tran (\sa_count[27][19] , \sa_count[27].r.part0[19] );
tran (\sa_count[27][19] , \sa_count[27].f.lower[19] );
tran (\sa_count[27][18] , \sa_count[27].r.part0[18] );
tran (\sa_count[27][18] , \sa_count[27].f.lower[18] );
tran (\sa_count[27][17] , \sa_count[27].r.part0[17] );
tran (\sa_count[27][17] , \sa_count[27].f.lower[17] );
tran (\sa_count[27][16] , \sa_count[27].r.part0[16] );
tran (\sa_count[27][16] , \sa_count[27].f.lower[16] );
tran (\sa_count[27][15] , \sa_count[27].r.part0[15] );
tran (\sa_count[27][15] , \sa_count[27].f.lower[15] );
tran (\sa_count[27][14] , \sa_count[27].r.part0[14] );
tran (\sa_count[27][14] , \sa_count[27].f.lower[14] );
tran (\sa_count[27][13] , \sa_count[27].r.part0[13] );
tran (\sa_count[27][13] , \sa_count[27].f.lower[13] );
tran (\sa_count[27][12] , \sa_count[27].r.part0[12] );
tran (\sa_count[27][12] , \sa_count[27].f.lower[12] );
tran (\sa_count[27][11] , \sa_count[27].r.part0[11] );
tran (\sa_count[27][11] , \sa_count[27].f.lower[11] );
tran (\sa_count[27][10] , \sa_count[27].r.part0[10] );
tran (\sa_count[27][10] , \sa_count[27].f.lower[10] );
tran (\sa_count[27][9] , \sa_count[27].r.part0[9] );
tran (\sa_count[27][9] , \sa_count[27].f.lower[9] );
tran (\sa_count[27][8] , \sa_count[27].r.part0[8] );
tran (\sa_count[27][8] , \sa_count[27].f.lower[8] );
tran (\sa_count[27][7] , \sa_count[27].r.part0[7] );
tran (\sa_count[27][7] , \sa_count[27].f.lower[7] );
tran (\sa_count[27][6] , \sa_count[27].r.part0[6] );
tran (\sa_count[27][6] , \sa_count[27].f.lower[6] );
tran (\sa_count[27][5] , \sa_count[27].r.part0[5] );
tran (\sa_count[27][5] , \sa_count[27].f.lower[5] );
tran (\sa_count[27][4] , \sa_count[27].r.part0[4] );
tran (\sa_count[27][4] , \sa_count[27].f.lower[4] );
tran (\sa_count[27][3] , \sa_count[27].r.part0[3] );
tran (\sa_count[27][3] , \sa_count[27].f.lower[3] );
tran (\sa_count[27][2] , \sa_count[27].r.part0[2] );
tran (\sa_count[27][2] , \sa_count[27].f.lower[2] );
tran (\sa_count[27][1] , \sa_count[27].r.part0[1] );
tran (\sa_count[27][1] , \sa_count[27].f.lower[1] );
tran (\sa_count[27][0] , \sa_count[27].r.part0[0] );
tran (\sa_count[27][0] , \sa_count[27].f.lower[0] );
tran (\sa_count[26][63] , \sa_count[26].r.part1[31] );
tran (\sa_count[26][63] , \sa_count[26].f.unused[13] );
tran (\sa_count[26][62] , \sa_count[26].r.part1[30] );
tran (\sa_count[26][62] , \sa_count[26].f.unused[12] );
tran (\sa_count[26][61] , \sa_count[26].r.part1[29] );
tran (\sa_count[26][61] , \sa_count[26].f.unused[11] );
tran (\sa_count[26][60] , \sa_count[26].r.part1[28] );
tran (\sa_count[26][60] , \sa_count[26].f.unused[10] );
tran (\sa_count[26][59] , \sa_count[26].r.part1[27] );
tran (\sa_count[26][59] , \sa_count[26].f.unused[9] );
tran (\sa_count[26][58] , \sa_count[26].r.part1[26] );
tran (\sa_count[26][58] , \sa_count[26].f.unused[8] );
tran (\sa_count[26][57] , \sa_count[26].r.part1[25] );
tran (\sa_count[26][57] , \sa_count[26].f.unused[7] );
tran (\sa_count[26][56] , \sa_count[26].r.part1[24] );
tran (\sa_count[26][56] , \sa_count[26].f.unused[6] );
tran (\sa_count[26][55] , \sa_count[26].r.part1[23] );
tran (\sa_count[26][55] , \sa_count[26].f.unused[5] );
tran (\sa_count[26][54] , \sa_count[26].r.part1[22] );
tran (\sa_count[26][54] , \sa_count[26].f.unused[4] );
tran (\sa_count[26][53] , \sa_count[26].r.part1[21] );
tran (\sa_count[26][53] , \sa_count[26].f.unused[3] );
tran (\sa_count[26][52] , \sa_count[26].r.part1[20] );
tran (\sa_count[26][52] , \sa_count[26].f.unused[2] );
tran (\sa_count[26][51] , \sa_count[26].r.part1[19] );
tran (\sa_count[26][51] , \sa_count[26].f.unused[1] );
tran (\sa_count[26][50] , \sa_count[26].r.part1[18] );
tran (\sa_count[26][50] , \sa_count[26].f.unused[0] );
tran (\sa_count[26][49] , \sa_count[26].r.part1[17] );
tran (\sa_count[26][49] , \sa_count[26].f.upper[17] );
tran (\sa_count[26][48] , \sa_count[26].r.part1[16] );
tran (\sa_count[26][48] , \sa_count[26].f.upper[16] );
tran (\sa_count[26][47] , \sa_count[26].r.part1[15] );
tran (\sa_count[26][47] , \sa_count[26].f.upper[15] );
tran (\sa_count[26][46] , \sa_count[26].r.part1[14] );
tran (\sa_count[26][46] , \sa_count[26].f.upper[14] );
tran (\sa_count[26][45] , \sa_count[26].r.part1[13] );
tran (\sa_count[26][45] , \sa_count[26].f.upper[13] );
tran (\sa_count[26][44] , \sa_count[26].r.part1[12] );
tran (\sa_count[26][44] , \sa_count[26].f.upper[12] );
tran (\sa_count[26][43] , \sa_count[26].r.part1[11] );
tran (\sa_count[26][43] , \sa_count[26].f.upper[11] );
tran (\sa_count[26][42] , \sa_count[26].r.part1[10] );
tran (\sa_count[26][42] , \sa_count[26].f.upper[10] );
tran (\sa_count[26][41] , \sa_count[26].r.part1[9] );
tran (\sa_count[26][41] , \sa_count[26].f.upper[9] );
tran (\sa_count[26][40] , \sa_count[26].r.part1[8] );
tran (\sa_count[26][40] , \sa_count[26].f.upper[8] );
tran (\sa_count[26][39] , \sa_count[26].r.part1[7] );
tran (\sa_count[26][39] , \sa_count[26].f.upper[7] );
tran (\sa_count[26][38] , \sa_count[26].r.part1[6] );
tran (\sa_count[26][38] , \sa_count[26].f.upper[6] );
tran (\sa_count[26][37] , \sa_count[26].r.part1[5] );
tran (\sa_count[26][37] , \sa_count[26].f.upper[5] );
tran (\sa_count[26][36] , \sa_count[26].r.part1[4] );
tran (\sa_count[26][36] , \sa_count[26].f.upper[4] );
tran (\sa_count[26][35] , \sa_count[26].r.part1[3] );
tran (\sa_count[26][35] , \sa_count[26].f.upper[3] );
tran (\sa_count[26][34] , \sa_count[26].r.part1[2] );
tran (\sa_count[26][34] , \sa_count[26].f.upper[2] );
tran (\sa_count[26][33] , \sa_count[26].r.part1[1] );
tran (\sa_count[26][33] , \sa_count[26].f.upper[1] );
tran (\sa_count[26][32] , \sa_count[26].r.part1[0] );
tran (\sa_count[26][32] , \sa_count[26].f.upper[0] );
tran (\sa_count[26][31] , \sa_count[26].r.part0[31] );
tran (\sa_count[26][31] , \sa_count[26].f.lower[31] );
tran (\sa_count[26][30] , \sa_count[26].r.part0[30] );
tran (\sa_count[26][30] , \sa_count[26].f.lower[30] );
tran (\sa_count[26][29] , \sa_count[26].r.part0[29] );
tran (\sa_count[26][29] , \sa_count[26].f.lower[29] );
tran (\sa_count[26][28] , \sa_count[26].r.part0[28] );
tran (\sa_count[26][28] , \sa_count[26].f.lower[28] );
tran (\sa_count[26][27] , \sa_count[26].r.part0[27] );
tran (\sa_count[26][27] , \sa_count[26].f.lower[27] );
tran (\sa_count[26][26] , \sa_count[26].r.part0[26] );
tran (\sa_count[26][26] , \sa_count[26].f.lower[26] );
tran (\sa_count[26][25] , \sa_count[26].r.part0[25] );
tran (\sa_count[26][25] , \sa_count[26].f.lower[25] );
tran (\sa_count[26][24] , \sa_count[26].r.part0[24] );
tran (\sa_count[26][24] , \sa_count[26].f.lower[24] );
tran (\sa_count[26][23] , \sa_count[26].r.part0[23] );
tran (\sa_count[26][23] , \sa_count[26].f.lower[23] );
tran (\sa_count[26][22] , \sa_count[26].r.part0[22] );
tran (\sa_count[26][22] , \sa_count[26].f.lower[22] );
tran (\sa_count[26][21] , \sa_count[26].r.part0[21] );
tran (\sa_count[26][21] , \sa_count[26].f.lower[21] );
tran (\sa_count[26][20] , \sa_count[26].r.part0[20] );
tran (\sa_count[26][20] , \sa_count[26].f.lower[20] );
tran (\sa_count[26][19] , \sa_count[26].r.part0[19] );
tran (\sa_count[26][19] , \sa_count[26].f.lower[19] );
tran (\sa_count[26][18] , \sa_count[26].r.part0[18] );
tran (\sa_count[26][18] , \sa_count[26].f.lower[18] );
tran (\sa_count[26][17] , \sa_count[26].r.part0[17] );
tran (\sa_count[26][17] , \sa_count[26].f.lower[17] );
tran (\sa_count[26][16] , \sa_count[26].r.part0[16] );
tran (\sa_count[26][16] , \sa_count[26].f.lower[16] );
tran (\sa_count[26][15] , \sa_count[26].r.part0[15] );
tran (\sa_count[26][15] , \sa_count[26].f.lower[15] );
tran (\sa_count[26][14] , \sa_count[26].r.part0[14] );
tran (\sa_count[26][14] , \sa_count[26].f.lower[14] );
tran (\sa_count[26][13] , \sa_count[26].r.part0[13] );
tran (\sa_count[26][13] , \sa_count[26].f.lower[13] );
tran (\sa_count[26][12] , \sa_count[26].r.part0[12] );
tran (\sa_count[26][12] , \sa_count[26].f.lower[12] );
tran (\sa_count[26][11] , \sa_count[26].r.part0[11] );
tran (\sa_count[26][11] , \sa_count[26].f.lower[11] );
tran (\sa_count[26][10] , \sa_count[26].r.part0[10] );
tran (\sa_count[26][10] , \sa_count[26].f.lower[10] );
tran (\sa_count[26][9] , \sa_count[26].r.part0[9] );
tran (\sa_count[26][9] , \sa_count[26].f.lower[9] );
tran (\sa_count[26][8] , \sa_count[26].r.part0[8] );
tran (\sa_count[26][8] , \sa_count[26].f.lower[8] );
tran (\sa_count[26][7] , \sa_count[26].r.part0[7] );
tran (\sa_count[26][7] , \sa_count[26].f.lower[7] );
tran (\sa_count[26][6] , \sa_count[26].r.part0[6] );
tran (\sa_count[26][6] , \sa_count[26].f.lower[6] );
tran (\sa_count[26][5] , \sa_count[26].r.part0[5] );
tran (\sa_count[26][5] , \sa_count[26].f.lower[5] );
tran (\sa_count[26][4] , \sa_count[26].r.part0[4] );
tran (\sa_count[26][4] , \sa_count[26].f.lower[4] );
tran (\sa_count[26][3] , \sa_count[26].r.part0[3] );
tran (\sa_count[26][3] , \sa_count[26].f.lower[3] );
tran (\sa_count[26][2] , \sa_count[26].r.part0[2] );
tran (\sa_count[26][2] , \sa_count[26].f.lower[2] );
tran (\sa_count[26][1] , \sa_count[26].r.part0[1] );
tran (\sa_count[26][1] , \sa_count[26].f.lower[1] );
tran (\sa_count[26][0] , \sa_count[26].r.part0[0] );
tran (\sa_count[26][0] , \sa_count[26].f.lower[0] );
tran (\sa_count[25][63] , \sa_count[25].r.part1[31] );
tran (\sa_count[25][63] , \sa_count[25].f.unused[13] );
tran (\sa_count[25][62] , \sa_count[25].r.part1[30] );
tran (\sa_count[25][62] , \sa_count[25].f.unused[12] );
tran (\sa_count[25][61] , \sa_count[25].r.part1[29] );
tran (\sa_count[25][61] , \sa_count[25].f.unused[11] );
tran (\sa_count[25][60] , \sa_count[25].r.part1[28] );
tran (\sa_count[25][60] , \sa_count[25].f.unused[10] );
tran (\sa_count[25][59] , \sa_count[25].r.part1[27] );
tran (\sa_count[25][59] , \sa_count[25].f.unused[9] );
tran (\sa_count[25][58] , \sa_count[25].r.part1[26] );
tran (\sa_count[25][58] , \sa_count[25].f.unused[8] );
tran (\sa_count[25][57] , \sa_count[25].r.part1[25] );
tran (\sa_count[25][57] , \sa_count[25].f.unused[7] );
tran (\sa_count[25][56] , \sa_count[25].r.part1[24] );
tran (\sa_count[25][56] , \sa_count[25].f.unused[6] );
tran (\sa_count[25][55] , \sa_count[25].r.part1[23] );
tran (\sa_count[25][55] , \sa_count[25].f.unused[5] );
tran (\sa_count[25][54] , \sa_count[25].r.part1[22] );
tran (\sa_count[25][54] , \sa_count[25].f.unused[4] );
tran (\sa_count[25][53] , \sa_count[25].r.part1[21] );
tran (\sa_count[25][53] , \sa_count[25].f.unused[3] );
tran (\sa_count[25][52] , \sa_count[25].r.part1[20] );
tran (\sa_count[25][52] , \sa_count[25].f.unused[2] );
tran (\sa_count[25][51] , \sa_count[25].r.part1[19] );
tran (\sa_count[25][51] , \sa_count[25].f.unused[1] );
tran (\sa_count[25][50] , \sa_count[25].r.part1[18] );
tran (\sa_count[25][50] , \sa_count[25].f.unused[0] );
tran (\sa_count[25][49] , \sa_count[25].r.part1[17] );
tran (\sa_count[25][49] , \sa_count[25].f.upper[17] );
tran (\sa_count[25][48] , \sa_count[25].r.part1[16] );
tran (\sa_count[25][48] , \sa_count[25].f.upper[16] );
tran (\sa_count[25][47] , \sa_count[25].r.part1[15] );
tran (\sa_count[25][47] , \sa_count[25].f.upper[15] );
tran (\sa_count[25][46] , \sa_count[25].r.part1[14] );
tran (\sa_count[25][46] , \sa_count[25].f.upper[14] );
tran (\sa_count[25][45] , \sa_count[25].r.part1[13] );
tran (\sa_count[25][45] , \sa_count[25].f.upper[13] );
tran (\sa_count[25][44] , \sa_count[25].r.part1[12] );
tran (\sa_count[25][44] , \sa_count[25].f.upper[12] );
tran (\sa_count[25][43] , \sa_count[25].r.part1[11] );
tran (\sa_count[25][43] , \sa_count[25].f.upper[11] );
tran (\sa_count[25][42] , \sa_count[25].r.part1[10] );
tran (\sa_count[25][42] , \sa_count[25].f.upper[10] );
tran (\sa_count[25][41] , \sa_count[25].r.part1[9] );
tran (\sa_count[25][41] , \sa_count[25].f.upper[9] );
tran (\sa_count[25][40] , \sa_count[25].r.part1[8] );
tran (\sa_count[25][40] , \sa_count[25].f.upper[8] );
tran (\sa_count[25][39] , \sa_count[25].r.part1[7] );
tran (\sa_count[25][39] , \sa_count[25].f.upper[7] );
tran (\sa_count[25][38] , \sa_count[25].r.part1[6] );
tran (\sa_count[25][38] , \sa_count[25].f.upper[6] );
tran (\sa_count[25][37] , \sa_count[25].r.part1[5] );
tran (\sa_count[25][37] , \sa_count[25].f.upper[5] );
tran (\sa_count[25][36] , \sa_count[25].r.part1[4] );
tran (\sa_count[25][36] , \sa_count[25].f.upper[4] );
tran (\sa_count[25][35] , \sa_count[25].r.part1[3] );
tran (\sa_count[25][35] , \sa_count[25].f.upper[3] );
tran (\sa_count[25][34] , \sa_count[25].r.part1[2] );
tran (\sa_count[25][34] , \sa_count[25].f.upper[2] );
tran (\sa_count[25][33] , \sa_count[25].r.part1[1] );
tran (\sa_count[25][33] , \sa_count[25].f.upper[1] );
tran (\sa_count[25][32] , \sa_count[25].r.part1[0] );
tran (\sa_count[25][32] , \sa_count[25].f.upper[0] );
tran (\sa_count[25][31] , \sa_count[25].r.part0[31] );
tran (\sa_count[25][31] , \sa_count[25].f.lower[31] );
tran (\sa_count[25][30] , \sa_count[25].r.part0[30] );
tran (\sa_count[25][30] , \sa_count[25].f.lower[30] );
tran (\sa_count[25][29] , \sa_count[25].r.part0[29] );
tran (\sa_count[25][29] , \sa_count[25].f.lower[29] );
tran (\sa_count[25][28] , \sa_count[25].r.part0[28] );
tran (\sa_count[25][28] , \sa_count[25].f.lower[28] );
tran (\sa_count[25][27] , \sa_count[25].r.part0[27] );
tran (\sa_count[25][27] , \sa_count[25].f.lower[27] );
tran (\sa_count[25][26] , \sa_count[25].r.part0[26] );
tran (\sa_count[25][26] , \sa_count[25].f.lower[26] );
tran (\sa_count[25][25] , \sa_count[25].r.part0[25] );
tran (\sa_count[25][25] , \sa_count[25].f.lower[25] );
tran (\sa_count[25][24] , \sa_count[25].r.part0[24] );
tran (\sa_count[25][24] , \sa_count[25].f.lower[24] );
tran (\sa_count[25][23] , \sa_count[25].r.part0[23] );
tran (\sa_count[25][23] , \sa_count[25].f.lower[23] );
tran (\sa_count[25][22] , \sa_count[25].r.part0[22] );
tran (\sa_count[25][22] , \sa_count[25].f.lower[22] );
tran (\sa_count[25][21] , \sa_count[25].r.part0[21] );
tran (\sa_count[25][21] , \sa_count[25].f.lower[21] );
tran (\sa_count[25][20] , \sa_count[25].r.part0[20] );
tran (\sa_count[25][20] , \sa_count[25].f.lower[20] );
tran (\sa_count[25][19] , \sa_count[25].r.part0[19] );
tran (\sa_count[25][19] , \sa_count[25].f.lower[19] );
tran (\sa_count[25][18] , \sa_count[25].r.part0[18] );
tran (\sa_count[25][18] , \sa_count[25].f.lower[18] );
tran (\sa_count[25][17] , \sa_count[25].r.part0[17] );
tran (\sa_count[25][17] , \sa_count[25].f.lower[17] );
tran (\sa_count[25][16] , \sa_count[25].r.part0[16] );
tran (\sa_count[25][16] , \sa_count[25].f.lower[16] );
tran (\sa_count[25][15] , \sa_count[25].r.part0[15] );
tran (\sa_count[25][15] , \sa_count[25].f.lower[15] );
tran (\sa_count[25][14] , \sa_count[25].r.part0[14] );
tran (\sa_count[25][14] , \sa_count[25].f.lower[14] );
tran (\sa_count[25][13] , \sa_count[25].r.part0[13] );
tran (\sa_count[25][13] , \sa_count[25].f.lower[13] );
tran (\sa_count[25][12] , \sa_count[25].r.part0[12] );
tran (\sa_count[25][12] , \sa_count[25].f.lower[12] );
tran (\sa_count[25][11] , \sa_count[25].r.part0[11] );
tran (\sa_count[25][11] , \sa_count[25].f.lower[11] );
tran (\sa_count[25][10] , \sa_count[25].r.part0[10] );
tran (\sa_count[25][10] , \sa_count[25].f.lower[10] );
tran (\sa_count[25][9] , \sa_count[25].r.part0[9] );
tran (\sa_count[25][9] , \sa_count[25].f.lower[9] );
tran (\sa_count[25][8] , \sa_count[25].r.part0[8] );
tran (\sa_count[25][8] , \sa_count[25].f.lower[8] );
tran (\sa_count[25][7] , \sa_count[25].r.part0[7] );
tran (\sa_count[25][7] , \sa_count[25].f.lower[7] );
tran (\sa_count[25][6] , \sa_count[25].r.part0[6] );
tran (\sa_count[25][6] , \sa_count[25].f.lower[6] );
tran (\sa_count[25][5] , \sa_count[25].r.part0[5] );
tran (\sa_count[25][5] , \sa_count[25].f.lower[5] );
tran (\sa_count[25][4] , \sa_count[25].r.part0[4] );
tran (\sa_count[25][4] , \sa_count[25].f.lower[4] );
tran (\sa_count[25][3] , \sa_count[25].r.part0[3] );
tran (\sa_count[25][3] , \sa_count[25].f.lower[3] );
tran (\sa_count[25][2] , \sa_count[25].r.part0[2] );
tran (\sa_count[25][2] , \sa_count[25].f.lower[2] );
tran (\sa_count[25][1] , \sa_count[25].r.part0[1] );
tran (\sa_count[25][1] , \sa_count[25].f.lower[1] );
tran (\sa_count[25][0] , \sa_count[25].r.part0[0] );
tran (\sa_count[25][0] , \sa_count[25].f.lower[0] );
tran (\sa_count[24][63] , \sa_count[24].r.part1[31] );
tran (\sa_count[24][63] , \sa_count[24].f.unused[13] );
tran (\sa_count[24][62] , \sa_count[24].r.part1[30] );
tran (\sa_count[24][62] , \sa_count[24].f.unused[12] );
tran (\sa_count[24][61] , \sa_count[24].r.part1[29] );
tran (\sa_count[24][61] , \sa_count[24].f.unused[11] );
tran (\sa_count[24][60] , \sa_count[24].r.part1[28] );
tran (\sa_count[24][60] , \sa_count[24].f.unused[10] );
tran (\sa_count[24][59] , \sa_count[24].r.part1[27] );
tran (\sa_count[24][59] , \sa_count[24].f.unused[9] );
tran (\sa_count[24][58] , \sa_count[24].r.part1[26] );
tran (\sa_count[24][58] , \sa_count[24].f.unused[8] );
tran (\sa_count[24][57] , \sa_count[24].r.part1[25] );
tran (\sa_count[24][57] , \sa_count[24].f.unused[7] );
tran (\sa_count[24][56] , \sa_count[24].r.part1[24] );
tran (\sa_count[24][56] , \sa_count[24].f.unused[6] );
tran (\sa_count[24][55] , \sa_count[24].r.part1[23] );
tran (\sa_count[24][55] , \sa_count[24].f.unused[5] );
tran (\sa_count[24][54] , \sa_count[24].r.part1[22] );
tran (\sa_count[24][54] , \sa_count[24].f.unused[4] );
tran (\sa_count[24][53] , \sa_count[24].r.part1[21] );
tran (\sa_count[24][53] , \sa_count[24].f.unused[3] );
tran (\sa_count[24][52] , \sa_count[24].r.part1[20] );
tran (\sa_count[24][52] , \sa_count[24].f.unused[2] );
tran (\sa_count[24][51] , \sa_count[24].r.part1[19] );
tran (\sa_count[24][51] , \sa_count[24].f.unused[1] );
tran (\sa_count[24][50] , \sa_count[24].r.part1[18] );
tran (\sa_count[24][50] , \sa_count[24].f.unused[0] );
tran (\sa_count[24][49] , \sa_count[24].r.part1[17] );
tran (\sa_count[24][49] , \sa_count[24].f.upper[17] );
tran (\sa_count[24][48] , \sa_count[24].r.part1[16] );
tran (\sa_count[24][48] , \sa_count[24].f.upper[16] );
tran (\sa_count[24][47] , \sa_count[24].r.part1[15] );
tran (\sa_count[24][47] , \sa_count[24].f.upper[15] );
tran (\sa_count[24][46] , \sa_count[24].r.part1[14] );
tran (\sa_count[24][46] , \sa_count[24].f.upper[14] );
tran (\sa_count[24][45] , \sa_count[24].r.part1[13] );
tran (\sa_count[24][45] , \sa_count[24].f.upper[13] );
tran (\sa_count[24][44] , \sa_count[24].r.part1[12] );
tran (\sa_count[24][44] , \sa_count[24].f.upper[12] );
tran (\sa_count[24][43] , \sa_count[24].r.part1[11] );
tran (\sa_count[24][43] , \sa_count[24].f.upper[11] );
tran (\sa_count[24][42] , \sa_count[24].r.part1[10] );
tran (\sa_count[24][42] , \sa_count[24].f.upper[10] );
tran (\sa_count[24][41] , \sa_count[24].r.part1[9] );
tran (\sa_count[24][41] , \sa_count[24].f.upper[9] );
tran (\sa_count[24][40] , \sa_count[24].r.part1[8] );
tran (\sa_count[24][40] , \sa_count[24].f.upper[8] );
tran (\sa_count[24][39] , \sa_count[24].r.part1[7] );
tran (\sa_count[24][39] , \sa_count[24].f.upper[7] );
tran (\sa_count[24][38] , \sa_count[24].r.part1[6] );
tran (\sa_count[24][38] , \sa_count[24].f.upper[6] );
tran (\sa_count[24][37] , \sa_count[24].r.part1[5] );
tran (\sa_count[24][37] , \sa_count[24].f.upper[5] );
tran (\sa_count[24][36] , \sa_count[24].r.part1[4] );
tran (\sa_count[24][36] , \sa_count[24].f.upper[4] );
tran (\sa_count[24][35] , \sa_count[24].r.part1[3] );
tran (\sa_count[24][35] , \sa_count[24].f.upper[3] );
tran (\sa_count[24][34] , \sa_count[24].r.part1[2] );
tran (\sa_count[24][34] , \sa_count[24].f.upper[2] );
tran (\sa_count[24][33] , \sa_count[24].r.part1[1] );
tran (\sa_count[24][33] , \sa_count[24].f.upper[1] );
tran (\sa_count[24][32] , \sa_count[24].r.part1[0] );
tran (\sa_count[24][32] , \sa_count[24].f.upper[0] );
tran (\sa_count[24][31] , \sa_count[24].r.part0[31] );
tran (\sa_count[24][31] , \sa_count[24].f.lower[31] );
tran (\sa_count[24][30] , \sa_count[24].r.part0[30] );
tran (\sa_count[24][30] , \sa_count[24].f.lower[30] );
tran (\sa_count[24][29] , \sa_count[24].r.part0[29] );
tran (\sa_count[24][29] , \sa_count[24].f.lower[29] );
tran (\sa_count[24][28] , \sa_count[24].r.part0[28] );
tran (\sa_count[24][28] , \sa_count[24].f.lower[28] );
tran (\sa_count[24][27] , \sa_count[24].r.part0[27] );
tran (\sa_count[24][27] , \sa_count[24].f.lower[27] );
tran (\sa_count[24][26] , \sa_count[24].r.part0[26] );
tran (\sa_count[24][26] , \sa_count[24].f.lower[26] );
tran (\sa_count[24][25] , \sa_count[24].r.part0[25] );
tran (\sa_count[24][25] , \sa_count[24].f.lower[25] );
tran (\sa_count[24][24] , \sa_count[24].r.part0[24] );
tran (\sa_count[24][24] , \sa_count[24].f.lower[24] );
tran (\sa_count[24][23] , \sa_count[24].r.part0[23] );
tran (\sa_count[24][23] , \sa_count[24].f.lower[23] );
tran (\sa_count[24][22] , \sa_count[24].r.part0[22] );
tran (\sa_count[24][22] , \sa_count[24].f.lower[22] );
tran (\sa_count[24][21] , \sa_count[24].r.part0[21] );
tran (\sa_count[24][21] , \sa_count[24].f.lower[21] );
tran (\sa_count[24][20] , \sa_count[24].r.part0[20] );
tran (\sa_count[24][20] , \sa_count[24].f.lower[20] );
tran (\sa_count[24][19] , \sa_count[24].r.part0[19] );
tran (\sa_count[24][19] , \sa_count[24].f.lower[19] );
tran (\sa_count[24][18] , \sa_count[24].r.part0[18] );
tran (\sa_count[24][18] , \sa_count[24].f.lower[18] );
tran (\sa_count[24][17] , \sa_count[24].r.part0[17] );
tran (\sa_count[24][17] , \sa_count[24].f.lower[17] );
tran (\sa_count[24][16] , \sa_count[24].r.part0[16] );
tran (\sa_count[24][16] , \sa_count[24].f.lower[16] );
tran (\sa_count[24][15] , \sa_count[24].r.part0[15] );
tran (\sa_count[24][15] , \sa_count[24].f.lower[15] );
tran (\sa_count[24][14] , \sa_count[24].r.part0[14] );
tran (\sa_count[24][14] , \sa_count[24].f.lower[14] );
tran (\sa_count[24][13] , \sa_count[24].r.part0[13] );
tran (\sa_count[24][13] , \sa_count[24].f.lower[13] );
tran (\sa_count[24][12] , \sa_count[24].r.part0[12] );
tran (\sa_count[24][12] , \sa_count[24].f.lower[12] );
tran (\sa_count[24][11] , \sa_count[24].r.part0[11] );
tran (\sa_count[24][11] , \sa_count[24].f.lower[11] );
tran (\sa_count[24][10] , \sa_count[24].r.part0[10] );
tran (\sa_count[24][10] , \sa_count[24].f.lower[10] );
tran (\sa_count[24][9] , \sa_count[24].r.part0[9] );
tran (\sa_count[24][9] , \sa_count[24].f.lower[9] );
tran (\sa_count[24][8] , \sa_count[24].r.part0[8] );
tran (\sa_count[24][8] , \sa_count[24].f.lower[8] );
tran (\sa_count[24][7] , \sa_count[24].r.part0[7] );
tran (\sa_count[24][7] , \sa_count[24].f.lower[7] );
tran (\sa_count[24][6] , \sa_count[24].r.part0[6] );
tran (\sa_count[24][6] , \sa_count[24].f.lower[6] );
tran (\sa_count[24][5] , \sa_count[24].r.part0[5] );
tran (\sa_count[24][5] , \sa_count[24].f.lower[5] );
tran (\sa_count[24][4] , \sa_count[24].r.part0[4] );
tran (\sa_count[24][4] , \sa_count[24].f.lower[4] );
tran (\sa_count[24][3] , \sa_count[24].r.part0[3] );
tran (\sa_count[24][3] , \sa_count[24].f.lower[3] );
tran (\sa_count[24][2] , \sa_count[24].r.part0[2] );
tran (\sa_count[24][2] , \sa_count[24].f.lower[2] );
tran (\sa_count[24][1] , \sa_count[24].r.part0[1] );
tran (\sa_count[24][1] , \sa_count[24].f.lower[1] );
tran (\sa_count[24][0] , \sa_count[24].r.part0[0] );
tran (\sa_count[24][0] , \sa_count[24].f.lower[0] );
tran (\sa_count[23][63] , \sa_count[23].r.part1[31] );
tran (\sa_count[23][63] , \sa_count[23].f.unused[13] );
tran (\sa_count[23][62] , \sa_count[23].r.part1[30] );
tran (\sa_count[23][62] , \sa_count[23].f.unused[12] );
tran (\sa_count[23][61] , \sa_count[23].r.part1[29] );
tran (\sa_count[23][61] , \sa_count[23].f.unused[11] );
tran (\sa_count[23][60] , \sa_count[23].r.part1[28] );
tran (\sa_count[23][60] , \sa_count[23].f.unused[10] );
tran (\sa_count[23][59] , \sa_count[23].r.part1[27] );
tran (\sa_count[23][59] , \sa_count[23].f.unused[9] );
tran (\sa_count[23][58] , \sa_count[23].r.part1[26] );
tran (\sa_count[23][58] , \sa_count[23].f.unused[8] );
tran (\sa_count[23][57] , \sa_count[23].r.part1[25] );
tran (\sa_count[23][57] , \sa_count[23].f.unused[7] );
tran (\sa_count[23][56] , \sa_count[23].r.part1[24] );
tran (\sa_count[23][56] , \sa_count[23].f.unused[6] );
tran (\sa_count[23][55] , \sa_count[23].r.part1[23] );
tran (\sa_count[23][55] , \sa_count[23].f.unused[5] );
tran (\sa_count[23][54] , \sa_count[23].r.part1[22] );
tran (\sa_count[23][54] , \sa_count[23].f.unused[4] );
tran (\sa_count[23][53] , \sa_count[23].r.part1[21] );
tran (\sa_count[23][53] , \sa_count[23].f.unused[3] );
tran (\sa_count[23][52] , \sa_count[23].r.part1[20] );
tran (\sa_count[23][52] , \sa_count[23].f.unused[2] );
tran (\sa_count[23][51] , \sa_count[23].r.part1[19] );
tran (\sa_count[23][51] , \sa_count[23].f.unused[1] );
tran (\sa_count[23][50] , \sa_count[23].r.part1[18] );
tran (\sa_count[23][50] , \sa_count[23].f.unused[0] );
tran (\sa_count[23][49] , \sa_count[23].r.part1[17] );
tran (\sa_count[23][49] , \sa_count[23].f.upper[17] );
tran (\sa_count[23][48] , \sa_count[23].r.part1[16] );
tran (\sa_count[23][48] , \sa_count[23].f.upper[16] );
tran (\sa_count[23][47] , \sa_count[23].r.part1[15] );
tran (\sa_count[23][47] , \sa_count[23].f.upper[15] );
tran (\sa_count[23][46] , \sa_count[23].r.part1[14] );
tran (\sa_count[23][46] , \sa_count[23].f.upper[14] );
tran (\sa_count[23][45] , \sa_count[23].r.part1[13] );
tran (\sa_count[23][45] , \sa_count[23].f.upper[13] );
tran (\sa_count[23][44] , \sa_count[23].r.part1[12] );
tran (\sa_count[23][44] , \sa_count[23].f.upper[12] );
tran (\sa_count[23][43] , \sa_count[23].r.part1[11] );
tran (\sa_count[23][43] , \sa_count[23].f.upper[11] );
tran (\sa_count[23][42] , \sa_count[23].r.part1[10] );
tran (\sa_count[23][42] , \sa_count[23].f.upper[10] );
tran (\sa_count[23][41] , \sa_count[23].r.part1[9] );
tran (\sa_count[23][41] , \sa_count[23].f.upper[9] );
tran (\sa_count[23][40] , \sa_count[23].r.part1[8] );
tran (\sa_count[23][40] , \sa_count[23].f.upper[8] );
tran (\sa_count[23][39] , \sa_count[23].r.part1[7] );
tran (\sa_count[23][39] , \sa_count[23].f.upper[7] );
tran (\sa_count[23][38] , \sa_count[23].r.part1[6] );
tran (\sa_count[23][38] , \sa_count[23].f.upper[6] );
tran (\sa_count[23][37] , \sa_count[23].r.part1[5] );
tran (\sa_count[23][37] , \sa_count[23].f.upper[5] );
tran (\sa_count[23][36] , \sa_count[23].r.part1[4] );
tran (\sa_count[23][36] , \sa_count[23].f.upper[4] );
tran (\sa_count[23][35] , \sa_count[23].r.part1[3] );
tran (\sa_count[23][35] , \sa_count[23].f.upper[3] );
tran (\sa_count[23][34] , \sa_count[23].r.part1[2] );
tran (\sa_count[23][34] , \sa_count[23].f.upper[2] );
tran (\sa_count[23][33] , \sa_count[23].r.part1[1] );
tran (\sa_count[23][33] , \sa_count[23].f.upper[1] );
tran (\sa_count[23][32] , \sa_count[23].r.part1[0] );
tran (\sa_count[23][32] , \sa_count[23].f.upper[0] );
tran (\sa_count[23][31] , \sa_count[23].r.part0[31] );
tran (\sa_count[23][31] , \sa_count[23].f.lower[31] );
tran (\sa_count[23][30] , \sa_count[23].r.part0[30] );
tran (\sa_count[23][30] , \sa_count[23].f.lower[30] );
tran (\sa_count[23][29] , \sa_count[23].r.part0[29] );
tran (\sa_count[23][29] , \sa_count[23].f.lower[29] );
tran (\sa_count[23][28] , \sa_count[23].r.part0[28] );
tran (\sa_count[23][28] , \sa_count[23].f.lower[28] );
tran (\sa_count[23][27] , \sa_count[23].r.part0[27] );
tran (\sa_count[23][27] , \sa_count[23].f.lower[27] );
tran (\sa_count[23][26] , \sa_count[23].r.part0[26] );
tran (\sa_count[23][26] , \sa_count[23].f.lower[26] );
tran (\sa_count[23][25] , \sa_count[23].r.part0[25] );
tran (\sa_count[23][25] , \sa_count[23].f.lower[25] );
tran (\sa_count[23][24] , \sa_count[23].r.part0[24] );
tran (\sa_count[23][24] , \sa_count[23].f.lower[24] );
tran (\sa_count[23][23] , \sa_count[23].r.part0[23] );
tran (\sa_count[23][23] , \sa_count[23].f.lower[23] );
tran (\sa_count[23][22] , \sa_count[23].r.part0[22] );
tran (\sa_count[23][22] , \sa_count[23].f.lower[22] );
tran (\sa_count[23][21] , \sa_count[23].r.part0[21] );
tran (\sa_count[23][21] , \sa_count[23].f.lower[21] );
tran (\sa_count[23][20] , \sa_count[23].r.part0[20] );
tran (\sa_count[23][20] , \sa_count[23].f.lower[20] );
tran (\sa_count[23][19] , \sa_count[23].r.part0[19] );
tran (\sa_count[23][19] , \sa_count[23].f.lower[19] );
tran (\sa_count[23][18] , \sa_count[23].r.part0[18] );
tran (\sa_count[23][18] , \sa_count[23].f.lower[18] );
tran (\sa_count[23][17] , \sa_count[23].r.part0[17] );
tran (\sa_count[23][17] , \sa_count[23].f.lower[17] );
tran (\sa_count[23][16] , \sa_count[23].r.part0[16] );
tran (\sa_count[23][16] , \sa_count[23].f.lower[16] );
tran (\sa_count[23][15] , \sa_count[23].r.part0[15] );
tran (\sa_count[23][15] , \sa_count[23].f.lower[15] );
tran (\sa_count[23][14] , \sa_count[23].r.part0[14] );
tran (\sa_count[23][14] , \sa_count[23].f.lower[14] );
tran (\sa_count[23][13] , \sa_count[23].r.part0[13] );
tran (\sa_count[23][13] , \sa_count[23].f.lower[13] );
tran (\sa_count[23][12] , \sa_count[23].r.part0[12] );
tran (\sa_count[23][12] , \sa_count[23].f.lower[12] );
tran (\sa_count[23][11] , \sa_count[23].r.part0[11] );
tran (\sa_count[23][11] , \sa_count[23].f.lower[11] );
tran (\sa_count[23][10] , \sa_count[23].r.part0[10] );
tran (\sa_count[23][10] , \sa_count[23].f.lower[10] );
tran (\sa_count[23][9] , \sa_count[23].r.part0[9] );
tran (\sa_count[23][9] , \sa_count[23].f.lower[9] );
tran (\sa_count[23][8] , \sa_count[23].r.part0[8] );
tran (\sa_count[23][8] , \sa_count[23].f.lower[8] );
tran (\sa_count[23][7] , \sa_count[23].r.part0[7] );
tran (\sa_count[23][7] , \sa_count[23].f.lower[7] );
tran (\sa_count[23][6] , \sa_count[23].r.part0[6] );
tran (\sa_count[23][6] , \sa_count[23].f.lower[6] );
tran (\sa_count[23][5] , \sa_count[23].r.part0[5] );
tran (\sa_count[23][5] , \sa_count[23].f.lower[5] );
tran (\sa_count[23][4] , \sa_count[23].r.part0[4] );
tran (\sa_count[23][4] , \sa_count[23].f.lower[4] );
tran (\sa_count[23][3] , \sa_count[23].r.part0[3] );
tran (\sa_count[23][3] , \sa_count[23].f.lower[3] );
tran (\sa_count[23][2] , \sa_count[23].r.part0[2] );
tran (\sa_count[23][2] , \sa_count[23].f.lower[2] );
tran (\sa_count[23][1] , \sa_count[23].r.part0[1] );
tran (\sa_count[23][1] , \sa_count[23].f.lower[1] );
tran (\sa_count[23][0] , \sa_count[23].r.part0[0] );
tran (\sa_count[23][0] , \sa_count[23].f.lower[0] );
tran (\sa_count[22][63] , \sa_count[22].r.part1[31] );
tran (\sa_count[22][63] , \sa_count[22].f.unused[13] );
tran (\sa_count[22][62] , \sa_count[22].r.part1[30] );
tran (\sa_count[22][62] , \sa_count[22].f.unused[12] );
tran (\sa_count[22][61] , \sa_count[22].r.part1[29] );
tran (\sa_count[22][61] , \sa_count[22].f.unused[11] );
tran (\sa_count[22][60] , \sa_count[22].r.part1[28] );
tran (\sa_count[22][60] , \sa_count[22].f.unused[10] );
tran (\sa_count[22][59] , \sa_count[22].r.part1[27] );
tran (\sa_count[22][59] , \sa_count[22].f.unused[9] );
tran (\sa_count[22][58] , \sa_count[22].r.part1[26] );
tran (\sa_count[22][58] , \sa_count[22].f.unused[8] );
tran (\sa_count[22][57] , \sa_count[22].r.part1[25] );
tran (\sa_count[22][57] , \sa_count[22].f.unused[7] );
tran (\sa_count[22][56] , \sa_count[22].r.part1[24] );
tran (\sa_count[22][56] , \sa_count[22].f.unused[6] );
tran (\sa_count[22][55] , \sa_count[22].r.part1[23] );
tran (\sa_count[22][55] , \sa_count[22].f.unused[5] );
tran (\sa_count[22][54] , \sa_count[22].r.part1[22] );
tran (\sa_count[22][54] , \sa_count[22].f.unused[4] );
tran (\sa_count[22][53] , \sa_count[22].r.part1[21] );
tran (\sa_count[22][53] , \sa_count[22].f.unused[3] );
tran (\sa_count[22][52] , \sa_count[22].r.part1[20] );
tran (\sa_count[22][52] , \sa_count[22].f.unused[2] );
tran (\sa_count[22][51] , \sa_count[22].r.part1[19] );
tran (\sa_count[22][51] , \sa_count[22].f.unused[1] );
tran (\sa_count[22][50] , \sa_count[22].r.part1[18] );
tran (\sa_count[22][50] , \sa_count[22].f.unused[0] );
tran (\sa_count[22][49] , \sa_count[22].r.part1[17] );
tran (\sa_count[22][49] , \sa_count[22].f.upper[17] );
tran (\sa_count[22][48] , \sa_count[22].r.part1[16] );
tran (\sa_count[22][48] , \sa_count[22].f.upper[16] );
tran (\sa_count[22][47] , \sa_count[22].r.part1[15] );
tran (\sa_count[22][47] , \sa_count[22].f.upper[15] );
tran (\sa_count[22][46] , \sa_count[22].r.part1[14] );
tran (\sa_count[22][46] , \sa_count[22].f.upper[14] );
tran (\sa_count[22][45] , \sa_count[22].r.part1[13] );
tran (\sa_count[22][45] , \sa_count[22].f.upper[13] );
tran (\sa_count[22][44] , \sa_count[22].r.part1[12] );
tran (\sa_count[22][44] , \sa_count[22].f.upper[12] );
tran (\sa_count[22][43] , \sa_count[22].r.part1[11] );
tran (\sa_count[22][43] , \sa_count[22].f.upper[11] );
tran (\sa_count[22][42] , \sa_count[22].r.part1[10] );
tran (\sa_count[22][42] , \sa_count[22].f.upper[10] );
tran (\sa_count[22][41] , \sa_count[22].r.part1[9] );
tran (\sa_count[22][41] , \sa_count[22].f.upper[9] );
tran (\sa_count[22][40] , \sa_count[22].r.part1[8] );
tran (\sa_count[22][40] , \sa_count[22].f.upper[8] );
tran (\sa_count[22][39] , \sa_count[22].r.part1[7] );
tran (\sa_count[22][39] , \sa_count[22].f.upper[7] );
tran (\sa_count[22][38] , \sa_count[22].r.part1[6] );
tran (\sa_count[22][38] , \sa_count[22].f.upper[6] );
tran (\sa_count[22][37] , \sa_count[22].r.part1[5] );
tran (\sa_count[22][37] , \sa_count[22].f.upper[5] );
tran (\sa_count[22][36] , \sa_count[22].r.part1[4] );
tran (\sa_count[22][36] , \sa_count[22].f.upper[4] );
tran (\sa_count[22][35] , \sa_count[22].r.part1[3] );
tran (\sa_count[22][35] , \sa_count[22].f.upper[3] );
tran (\sa_count[22][34] , \sa_count[22].r.part1[2] );
tran (\sa_count[22][34] , \sa_count[22].f.upper[2] );
tran (\sa_count[22][33] , \sa_count[22].r.part1[1] );
tran (\sa_count[22][33] , \sa_count[22].f.upper[1] );
tran (\sa_count[22][32] , \sa_count[22].r.part1[0] );
tran (\sa_count[22][32] , \sa_count[22].f.upper[0] );
tran (\sa_count[22][31] , \sa_count[22].r.part0[31] );
tran (\sa_count[22][31] , \sa_count[22].f.lower[31] );
tran (\sa_count[22][30] , \sa_count[22].r.part0[30] );
tran (\sa_count[22][30] , \sa_count[22].f.lower[30] );
tran (\sa_count[22][29] , \sa_count[22].r.part0[29] );
tran (\sa_count[22][29] , \sa_count[22].f.lower[29] );
tran (\sa_count[22][28] , \sa_count[22].r.part0[28] );
tran (\sa_count[22][28] , \sa_count[22].f.lower[28] );
tran (\sa_count[22][27] , \sa_count[22].r.part0[27] );
tran (\sa_count[22][27] , \sa_count[22].f.lower[27] );
tran (\sa_count[22][26] , \sa_count[22].r.part0[26] );
tran (\sa_count[22][26] , \sa_count[22].f.lower[26] );
tran (\sa_count[22][25] , \sa_count[22].r.part0[25] );
tran (\sa_count[22][25] , \sa_count[22].f.lower[25] );
tran (\sa_count[22][24] , \sa_count[22].r.part0[24] );
tran (\sa_count[22][24] , \sa_count[22].f.lower[24] );
tran (\sa_count[22][23] , \sa_count[22].r.part0[23] );
tran (\sa_count[22][23] , \sa_count[22].f.lower[23] );
tran (\sa_count[22][22] , \sa_count[22].r.part0[22] );
tran (\sa_count[22][22] , \sa_count[22].f.lower[22] );
tran (\sa_count[22][21] , \sa_count[22].r.part0[21] );
tran (\sa_count[22][21] , \sa_count[22].f.lower[21] );
tran (\sa_count[22][20] , \sa_count[22].r.part0[20] );
tran (\sa_count[22][20] , \sa_count[22].f.lower[20] );
tran (\sa_count[22][19] , \sa_count[22].r.part0[19] );
tran (\sa_count[22][19] , \sa_count[22].f.lower[19] );
tran (\sa_count[22][18] , \sa_count[22].r.part0[18] );
tran (\sa_count[22][18] , \sa_count[22].f.lower[18] );
tran (\sa_count[22][17] , \sa_count[22].r.part0[17] );
tran (\sa_count[22][17] , \sa_count[22].f.lower[17] );
tran (\sa_count[22][16] , \sa_count[22].r.part0[16] );
tran (\sa_count[22][16] , \sa_count[22].f.lower[16] );
tran (\sa_count[22][15] , \sa_count[22].r.part0[15] );
tran (\sa_count[22][15] , \sa_count[22].f.lower[15] );
tran (\sa_count[22][14] , \sa_count[22].r.part0[14] );
tran (\sa_count[22][14] , \sa_count[22].f.lower[14] );
tran (\sa_count[22][13] , \sa_count[22].r.part0[13] );
tran (\sa_count[22][13] , \sa_count[22].f.lower[13] );
tran (\sa_count[22][12] , \sa_count[22].r.part0[12] );
tran (\sa_count[22][12] , \sa_count[22].f.lower[12] );
tran (\sa_count[22][11] , \sa_count[22].r.part0[11] );
tran (\sa_count[22][11] , \sa_count[22].f.lower[11] );
tran (\sa_count[22][10] , \sa_count[22].r.part0[10] );
tran (\sa_count[22][10] , \sa_count[22].f.lower[10] );
tran (\sa_count[22][9] , \sa_count[22].r.part0[9] );
tran (\sa_count[22][9] , \sa_count[22].f.lower[9] );
tran (\sa_count[22][8] , \sa_count[22].r.part0[8] );
tran (\sa_count[22][8] , \sa_count[22].f.lower[8] );
tran (\sa_count[22][7] , \sa_count[22].r.part0[7] );
tran (\sa_count[22][7] , \sa_count[22].f.lower[7] );
tran (\sa_count[22][6] , \sa_count[22].r.part0[6] );
tran (\sa_count[22][6] , \sa_count[22].f.lower[6] );
tran (\sa_count[22][5] , \sa_count[22].r.part0[5] );
tran (\sa_count[22][5] , \sa_count[22].f.lower[5] );
tran (\sa_count[22][4] , \sa_count[22].r.part0[4] );
tran (\sa_count[22][4] , \sa_count[22].f.lower[4] );
tran (\sa_count[22][3] , \sa_count[22].r.part0[3] );
tran (\sa_count[22][3] , \sa_count[22].f.lower[3] );
tran (\sa_count[22][2] , \sa_count[22].r.part0[2] );
tran (\sa_count[22][2] , \sa_count[22].f.lower[2] );
tran (\sa_count[22][1] , \sa_count[22].r.part0[1] );
tran (\sa_count[22][1] , \sa_count[22].f.lower[1] );
tran (\sa_count[22][0] , \sa_count[22].r.part0[0] );
tran (\sa_count[22][0] , \sa_count[22].f.lower[0] );
tran (\sa_count[21][63] , \sa_count[21].r.part1[31] );
tran (\sa_count[21][63] , \sa_count[21].f.unused[13] );
tran (\sa_count[21][62] , \sa_count[21].r.part1[30] );
tran (\sa_count[21][62] , \sa_count[21].f.unused[12] );
tran (\sa_count[21][61] , \sa_count[21].r.part1[29] );
tran (\sa_count[21][61] , \sa_count[21].f.unused[11] );
tran (\sa_count[21][60] , \sa_count[21].r.part1[28] );
tran (\sa_count[21][60] , \sa_count[21].f.unused[10] );
tran (\sa_count[21][59] , \sa_count[21].r.part1[27] );
tran (\sa_count[21][59] , \sa_count[21].f.unused[9] );
tran (\sa_count[21][58] , \sa_count[21].r.part1[26] );
tran (\sa_count[21][58] , \sa_count[21].f.unused[8] );
tran (\sa_count[21][57] , \sa_count[21].r.part1[25] );
tran (\sa_count[21][57] , \sa_count[21].f.unused[7] );
tran (\sa_count[21][56] , \sa_count[21].r.part1[24] );
tran (\sa_count[21][56] , \sa_count[21].f.unused[6] );
tran (\sa_count[21][55] , \sa_count[21].r.part1[23] );
tran (\sa_count[21][55] , \sa_count[21].f.unused[5] );
tran (\sa_count[21][54] , \sa_count[21].r.part1[22] );
tran (\sa_count[21][54] , \sa_count[21].f.unused[4] );
tran (\sa_count[21][53] , \sa_count[21].r.part1[21] );
tran (\sa_count[21][53] , \sa_count[21].f.unused[3] );
tran (\sa_count[21][52] , \sa_count[21].r.part1[20] );
tran (\sa_count[21][52] , \sa_count[21].f.unused[2] );
tran (\sa_count[21][51] , \sa_count[21].r.part1[19] );
tran (\sa_count[21][51] , \sa_count[21].f.unused[1] );
tran (\sa_count[21][50] , \sa_count[21].r.part1[18] );
tran (\sa_count[21][50] , \sa_count[21].f.unused[0] );
tran (\sa_count[21][49] , \sa_count[21].r.part1[17] );
tran (\sa_count[21][49] , \sa_count[21].f.upper[17] );
tran (\sa_count[21][48] , \sa_count[21].r.part1[16] );
tran (\sa_count[21][48] , \sa_count[21].f.upper[16] );
tran (\sa_count[21][47] , \sa_count[21].r.part1[15] );
tran (\sa_count[21][47] , \sa_count[21].f.upper[15] );
tran (\sa_count[21][46] , \sa_count[21].r.part1[14] );
tran (\sa_count[21][46] , \sa_count[21].f.upper[14] );
tran (\sa_count[21][45] , \sa_count[21].r.part1[13] );
tran (\sa_count[21][45] , \sa_count[21].f.upper[13] );
tran (\sa_count[21][44] , \sa_count[21].r.part1[12] );
tran (\sa_count[21][44] , \sa_count[21].f.upper[12] );
tran (\sa_count[21][43] , \sa_count[21].r.part1[11] );
tran (\sa_count[21][43] , \sa_count[21].f.upper[11] );
tran (\sa_count[21][42] , \sa_count[21].r.part1[10] );
tran (\sa_count[21][42] , \sa_count[21].f.upper[10] );
tran (\sa_count[21][41] , \sa_count[21].r.part1[9] );
tran (\sa_count[21][41] , \sa_count[21].f.upper[9] );
tran (\sa_count[21][40] , \sa_count[21].r.part1[8] );
tran (\sa_count[21][40] , \sa_count[21].f.upper[8] );
tran (\sa_count[21][39] , \sa_count[21].r.part1[7] );
tran (\sa_count[21][39] , \sa_count[21].f.upper[7] );
tran (\sa_count[21][38] , \sa_count[21].r.part1[6] );
tran (\sa_count[21][38] , \sa_count[21].f.upper[6] );
tran (\sa_count[21][37] , \sa_count[21].r.part1[5] );
tran (\sa_count[21][37] , \sa_count[21].f.upper[5] );
tran (\sa_count[21][36] , \sa_count[21].r.part1[4] );
tran (\sa_count[21][36] , \sa_count[21].f.upper[4] );
tran (\sa_count[21][35] , \sa_count[21].r.part1[3] );
tran (\sa_count[21][35] , \sa_count[21].f.upper[3] );
tran (\sa_count[21][34] , \sa_count[21].r.part1[2] );
tran (\sa_count[21][34] , \sa_count[21].f.upper[2] );
tran (\sa_count[21][33] , \sa_count[21].r.part1[1] );
tran (\sa_count[21][33] , \sa_count[21].f.upper[1] );
tran (\sa_count[21][32] , \sa_count[21].r.part1[0] );
tran (\sa_count[21][32] , \sa_count[21].f.upper[0] );
tran (\sa_count[21][31] , \sa_count[21].r.part0[31] );
tran (\sa_count[21][31] , \sa_count[21].f.lower[31] );
tran (\sa_count[21][30] , \sa_count[21].r.part0[30] );
tran (\sa_count[21][30] , \sa_count[21].f.lower[30] );
tran (\sa_count[21][29] , \sa_count[21].r.part0[29] );
tran (\sa_count[21][29] , \sa_count[21].f.lower[29] );
tran (\sa_count[21][28] , \sa_count[21].r.part0[28] );
tran (\sa_count[21][28] , \sa_count[21].f.lower[28] );
tran (\sa_count[21][27] , \sa_count[21].r.part0[27] );
tran (\sa_count[21][27] , \sa_count[21].f.lower[27] );
tran (\sa_count[21][26] , \sa_count[21].r.part0[26] );
tran (\sa_count[21][26] , \sa_count[21].f.lower[26] );
tran (\sa_count[21][25] , \sa_count[21].r.part0[25] );
tran (\sa_count[21][25] , \sa_count[21].f.lower[25] );
tran (\sa_count[21][24] , \sa_count[21].r.part0[24] );
tran (\sa_count[21][24] , \sa_count[21].f.lower[24] );
tran (\sa_count[21][23] , \sa_count[21].r.part0[23] );
tran (\sa_count[21][23] , \sa_count[21].f.lower[23] );
tran (\sa_count[21][22] , \sa_count[21].r.part0[22] );
tran (\sa_count[21][22] , \sa_count[21].f.lower[22] );
tran (\sa_count[21][21] , \sa_count[21].r.part0[21] );
tran (\sa_count[21][21] , \sa_count[21].f.lower[21] );
tran (\sa_count[21][20] , \sa_count[21].r.part0[20] );
tran (\sa_count[21][20] , \sa_count[21].f.lower[20] );
tran (\sa_count[21][19] , \sa_count[21].r.part0[19] );
tran (\sa_count[21][19] , \sa_count[21].f.lower[19] );
tran (\sa_count[21][18] , \sa_count[21].r.part0[18] );
tran (\sa_count[21][18] , \sa_count[21].f.lower[18] );
tran (\sa_count[21][17] , \sa_count[21].r.part0[17] );
tran (\sa_count[21][17] , \sa_count[21].f.lower[17] );
tran (\sa_count[21][16] , \sa_count[21].r.part0[16] );
tran (\sa_count[21][16] , \sa_count[21].f.lower[16] );
tran (\sa_count[21][15] , \sa_count[21].r.part0[15] );
tran (\sa_count[21][15] , \sa_count[21].f.lower[15] );
tran (\sa_count[21][14] , \sa_count[21].r.part0[14] );
tran (\sa_count[21][14] , \sa_count[21].f.lower[14] );
tran (\sa_count[21][13] , \sa_count[21].r.part0[13] );
tran (\sa_count[21][13] , \sa_count[21].f.lower[13] );
tran (\sa_count[21][12] , \sa_count[21].r.part0[12] );
tran (\sa_count[21][12] , \sa_count[21].f.lower[12] );
tran (\sa_count[21][11] , \sa_count[21].r.part0[11] );
tran (\sa_count[21][11] , \sa_count[21].f.lower[11] );
tran (\sa_count[21][10] , \sa_count[21].r.part0[10] );
tran (\sa_count[21][10] , \sa_count[21].f.lower[10] );
tran (\sa_count[21][9] , \sa_count[21].r.part0[9] );
tran (\sa_count[21][9] , \sa_count[21].f.lower[9] );
tran (\sa_count[21][8] , \sa_count[21].r.part0[8] );
tran (\sa_count[21][8] , \sa_count[21].f.lower[8] );
tran (\sa_count[21][7] , \sa_count[21].r.part0[7] );
tran (\sa_count[21][7] , \sa_count[21].f.lower[7] );
tran (\sa_count[21][6] , \sa_count[21].r.part0[6] );
tran (\sa_count[21][6] , \sa_count[21].f.lower[6] );
tran (\sa_count[21][5] , \sa_count[21].r.part0[5] );
tran (\sa_count[21][5] , \sa_count[21].f.lower[5] );
tran (\sa_count[21][4] , \sa_count[21].r.part0[4] );
tran (\sa_count[21][4] , \sa_count[21].f.lower[4] );
tran (\sa_count[21][3] , \sa_count[21].r.part0[3] );
tran (\sa_count[21][3] , \sa_count[21].f.lower[3] );
tran (\sa_count[21][2] , \sa_count[21].r.part0[2] );
tran (\sa_count[21][2] , \sa_count[21].f.lower[2] );
tran (\sa_count[21][1] , \sa_count[21].r.part0[1] );
tran (\sa_count[21][1] , \sa_count[21].f.lower[1] );
tran (\sa_count[21][0] , \sa_count[21].r.part0[0] );
tran (\sa_count[21][0] , \sa_count[21].f.lower[0] );
tran (\sa_count[20][63] , \sa_count[20].r.part1[31] );
tran (\sa_count[20][63] , \sa_count[20].f.unused[13] );
tran (\sa_count[20][62] , \sa_count[20].r.part1[30] );
tran (\sa_count[20][62] , \sa_count[20].f.unused[12] );
tran (\sa_count[20][61] , \sa_count[20].r.part1[29] );
tran (\sa_count[20][61] , \sa_count[20].f.unused[11] );
tran (\sa_count[20][60] , \sa_count[20].r.part1[28] );
tran (\sa_count[20][60] , \sa_count[20].f.unused[10] );
tran (\sa_count[20][59] , \sa_count[20].r.part1[27] );
tran (\sa_count[20][59] , \sa_count[20].f.unused[9] );
tran (\sa_count[20][58] , \sa_count[20].r.part1[26] );
tran (\sa_count[20][58] , \sa_count[20].f.unused[8] );
tran (\sa_count[20][57] , \sa_count[20].r.part1[25] );
tran (\sa_count[20][57] , \sa_count[20].f.unused[7] );
tran (\sa_count[20][56] , \sa_count[20].r.part1[24] );
tran (\sa_count[20][56] , \sa_count[20].f.unused[6] );
tran (\sa_count[20][55] , \sa_count[20].r.part1[23] );
tran (\sa_count[20][55] , \sa_count[20].f.unused[5] );
tran (\sa_count[20][54] , \sa_count[20].r.part1[22] );
tran (\sa_count[20][54] , \sa_count[20].f.unused[4] );
tran (\sa_count[20][53] , \sa_count[20].r.part1[21] );
tran (\sa_count[20][53] , \sa_count[20].f.unused[3] );
tran (\sa_count[20][52] , \sa_count[20].r.part1[20] );
tran (\sa_count[20][52] , \sa_count[20].f.unused[2] );
tran (\sa_count[20][51] , \sa_count[20].r.part1[19] );
tran (\sa_count[20][51] , \sa_count[20].f.unused[1] );
tran (\sa_count[20][50] , \sa_count[20].r.part1[18] );
tran (\sa_count[20][50] , \sa_count[20].f.unused[0] );
tran (\sa_count[20][49] , \sa_count[20].r.part1[17] );
tran (\sa_count[20][49] , \sa_count[20].f.upper[17] );
tran (\sa_count[20][48] , \sa_count[20].r.part1[16] );
tran (\sa_count[20][48] , \sa_count[20].f.upper[16] );
tran (\sa_count[20][47] , \sa_count[20].r.part1[15] );
tran (\sa_count[20][47] , \sa_count[20].f.upper[15] );
tran (\sa_count[20][46] , \sa_count[20].r.part1[14] );
tran (\sa_count[20][46] , \sa_count[20].f.upper[14] );
tran (\sa_count[20][45] , \sa_count[20].r.part1[13] );
tran (\sa_count[20][45] , \sa_count[20].f.upper[13] );
tran (\sa_count[20][44] , \sa_count[20].r.part1[12] );
tran (\sa_count[20][44] , \sa_count[20].f.upper[12] );
tran (\sa_count[20][43] , \sa_count[20].r.part1[11] );
tran (\sa_count[20][43] , \sa_count[20].f.upper[11] );
tran (\sa_count[20][42] , \sa_count[20].r.part1[10] );
tran (\sa_count[20][42] , \sa_count[20].f.upper[10] );
tran (\sa_count[20][41] , \sa_count[20].r.part1[9] );
tran (\sa_count[20][41] , \sa_count[20].f.upper[9] );
tran (\sa_count[20][40] , \sa_count[20].r.part1[8] );
tran (\sa_count[20][40] , \sa_count[20].f.upper[8] );
tran (\sa_count[20][39] , \sa_count[20].r.part1[7] );
tran (\sa_count[20][39] , \sa_count[20].f.upper[7] );
tran (\sa_count[20][38] , \sa_count[20].r.part1[6] );
tran (\sa_count[20][38] , \sa_count[20].f.upper[6] );
tran (\sa_count[20][37] , \sa_count[20].r.part1[5] );
tran (\sa_count[20][37] , \sa_count[20].f.upper[5] );
tran (\sa_count[20][36] , \sa_count[20].r.part1[4] );
tran (\sa_count[20][36] , \sa_count[20].f.upper[4] );
tran (\sa_count[20][35] , \sa_count[20].r.part1[3] );
tran (\sa_count[20][35] , \sa_count[20].f.upper[3] );
tran (\sa_count[20][34] , \sa_count[20].r.part1[2] );
tran (\sa_count[20][34] , \sa_count[20].f.upper[2] );
tran (\sa_count[20][33] , \sa_count[20].r.part1[1] );
tran (\sa_count[20][33] , \sa_count[20].f.upper[1] );
tran (\sa_count[20][32] , \sa_count[20].r.part1[0] );
tran (\sa_count[20][32] , \sa_count[20].f.upper[0] );
tran (\sa_count[20][31] , \sa_count[20].r.part0[31] );
tran (\sa_count[20][31] , \sa_count[20].f.lower[31] );
tran (\sa_count[20][30] , \sa_count[20].r.part0[30] );
tran (\sa_count[20][30] , \sa_count[20].f.lower[30] );
tran (\sa_count[20][29] , \sa_count[20].r.part0[29] );
tran (\sa_count[20][29] , \sa_count[20].f.lower[29] );
tran (\sa_count[20][28] , \sa_count[20].r.part0[28] );
tran (\sa_count[20][28] , \sa_count[20].f.lower[28] );
tran (\sa_count[20][27] , \sa_count[20].r.part0[27] );
tran (\sa_count[20][27] , \sa_count[20].f.lower[27] );
tran (\sa_count[20][26] , \sa_count[20].r.part0[26] );
tran (\sa_count[20][26] , \sa_count[20].f.lower[26] );
tran (\sa_count[20][25] , \sa_count[20].r.part0[25] );
tran (\sa_count[20][25] , \sa_count[20].f.lower[25] );
tran (\sa_count[20][24] , \sa_count[20].r.part0[24] );
tran (\sa_count[20][24] , \sa_count[20].f.lower[24] );
tran (\sa_count[20][23] , \sa_count[20].r.part0[23] );
tran (\sa_count[20][23] , \sa_count[20].f.lower[23] );
tran (\sa_count[20][22] , \sa_count[20].r.part0[22] );
tran (\sa_count[20][22] , \sa_count[20].f.lower[22] );
tran (\sa_count[20][21] , \sa_count[20].r.part0[21] );
tran (\sa_count[20][21] , \sa_count[20].f.lower[21] );
tran (\sa_count[20][20] , \sa_count[20].r.part0[20] );
tran (\sa_count[20][20] , \sa_count[20].f.lower[20] );
tran (\sa_count[20][19] , \sa_count[20].r.part0[19] );
tran (\sa_count[20][19] , \sa_count[20].f.lower[19] );
tran (\sa_count[20][18] , \sa_count[20].r.part0[18] );
tran (\sa_count[20][18] , \sa_count[20].f.lower[18] );
tran (\sa_count[20][17] , \sa_count[20].r.part0[17] );
tran (\sa_count[20][17] , \sa_count[20].f.lower[17] );
tran (\sa_count[20][16] , \sa_count[20].r.part0[16] );
tran (\sa_count[20][16] , \sa_count[20].f.lower[16] );
tran (\sa_count[20][15] , \sa_count[20].r.part0[15] );
tran (\sa_count[20][15] , \sa_count[20].f.lower[15] );
tran (\sa_count[20][14] , \sa_count[20].r.part0[14] );
tran (\sa_count[20][14] , \sa_count[20].f.lower[14] );
tran (\sa_count[20][13] , \sa_count[20].r.part0[13] );
tran (\sa_count[20][13] , \sa_count[20].f.lower[13] );
tran (\sa_count[20][12] , \sa_count[20].r.part0[12] );
tran (\sa_count[20][12] , \sa_count[20].f.lower[12] );
tran (\sa_count[20][11] , \sa_count[20].r.part0[11] );
tran (\sa_count[20][11] , \sa_count[20].f.lower[11] );
tran (\sa_count[20][10] , \sa_count[20].r.part0[10] );
tran (\sa_count[20][10] , \sa_count[20].f.lower[10] );
tran (\sa_count[20][9] , \sa_count[20].r.part0[9] );
tran (\sa_count[20][9] , \sa_count[20].f.lower[9] );
tran (\sa_count[20][8] , \sa_count[20].r.part0[8] );
tran (\sa_count[20][8] , \sa_count[20].f.lower[8] );
tran (\sa_count[20][7] , \sa_count[20].r.part0[7] );
tran (\sa_count[20][7] , \sa_count[20].f.lower[7] );
tran (\sa_count[20][6] , \sa_count[20].r.part0[6] );
tran (\sa_count[20][6] , \sa_count[20].f.lower[6] );
tran (\sa_count[20][5] , \sa_count[20].r.part0[5] );
tran (\sa_count[20][5] , \sa_count[20].f.lower[5] );
tran (\sa_count[20][4] , \sa_count[20].r.part0[4] );
tran (\sa_count[20][4] , \sa_count[20].f.lower[4] );
tran (\sa_count[20][3] , \sa_count[20].r.part0[3] );
tran (\sa_count[20][3] , \sa_count[20].f.lower[3] );
tran (\sa_count[20][2] , \sa_count[20].r.part0[2] );
tran (\sa_count[20][2] , \sa_count[20].f.lower[2] );
tran (\sa_count[20][1] , \sa_count[20].r.part0[1] );
tran (\sa_count[20][1] , \sa_count[20].f.lower[1] );
tran (\sa_count[20][0] , \sa_count[20].r.part0[0] );
tran (\sa_count[20][0] , \sa_count[20].f.lower[0] );
tran (\sa_count[19][63] , \sa_count[19].r.part1[31] );
tran (\sa_count[19][63] , \sa_count[19].f.unused[13] );
tran (\sa_count[19][62] , \sa_count[19].r.part1[30] );
tran (\sa_count[19][62] , \sa_count[19].f.unused[12] );
tran (\sa_count[19][61] , \sa_count[19].r.part1[29] );
tran (\sa_count[19][61] , \sa_count[19].f.unused[11] );
tran (\sa_count[19][60] , \sa_count[19].r.part1[28] );
tran (\sa_count[19][60] , \sa_count[19].f.unused[10] );
tran (\sa_count[19][59] , \sa_count[19].r.part1[27] );
tran (\sa_count[19][59] , \sa_count[19].f.unused[9] );
tran (\sa_count[19][58] , \sa_count[19].r.part1[26] );
tran (\sa_count[19][58] , \sa_count[19].f.unused[8] );
tran (\sa_count[19][57] , \sa_count[19].r.part1[25] );
tran (\sa_count[19][57] , \sa_count[19].f.unused[7] );
tran (\sa_count[19][56] , \sa_count[19].r.part1[24] );
tran (\sa_count[19][56] , \sa_count[19].f.unused[6] );
tran (\sa_count[19][55] , \sa_count[19].r.part1[23] );
tran (\sa_count[19][55] , \sa_count[19].f.unused[5] );
tran (\sa_count[19][54] , \sa_count[19].r.part1[22] );
tran (\sa_count[19][54] , \sa_count[19].f.unused[4] );
tran (\sa_count[19][53] , \sa_count[19].r.part1[21] );
tran (\sa_count[19][53] , \sa_count[19].f.unused[3] );
tran (\sa_count[19][52] , \sa_count[19].r.part1[20] );
tran (\sa_count[19][52] , \sa_count[19].f.unused[2] );
tran (\sa_count[19][51] , \sa_count[19].r.part1[19] );
tran (\sa_count[19][51] , \sa_count[19].f.unused[1] );
tran (\sa_count[19][50] , \sa_count[19].r.part1[18] );
tran (\sa_count[19][50] , \sa_count[19].f.unused[0] );
tran (\sa_count[19][49] , \sa_count[19].r.part1[17] );
tran (\sa_count[19][49] , \sa_count[19].f.upper[17] );
tran (\sa_count[19][48] , \sa_count[19].r.part1[16] );
tran (\sa_count[19][48] , \sa_count[19].f.upper[16] );
tran (\sa_count[19][47] , \sa_count[19].r.part1[15] );
tran (\sa_count[19][47] , \sa_count[19].f.upper[15] );
tran (\sa_count[19][46] , \sa_count[19].r.part1[14] );
tran (\sa_count[19][46] , \sa_count[19].f.upper[14] );
tran (\sa_count[19][45] , \sa_count[19].r.part1[13] );
tran (\sa_count[19][45] , \sa_count[19].f.upper[13] );
tran (\sa_count[19][44] , \sa_count[19].r.part1[12] );
tran (\sa_count[19][44] , \sa_count[19].f.upper[12] );
tran (\sa_count[19][43] , \sa_count[19].r.part1[11] );
tran (\sa_count[19][43] , \sa_count[19].f.upper[11] );
tran (\sa_count[19][42] , \sa_count[19].r.part1[10] );
tran (\sa_count[19][42] , \sa_count[19].f.upper[10] );
tran (\sa_count[19][41] , \sa_count[19].r.part1[9] );
tran (\sa_count[19][41] , \sa_count[19].f.upper[9] );
tran (\sa_count[19][40] , \sa_count[19].r.part1[8] );
tran (\sa_count[19][40] , \sa_count[19].f.upper[8] );
tran (\sa_count[19][39] , \sa_count[19].r.part1[7] );
tran (\sa_count[19][39] , \sa_count[19].f.upper[7] );
tran (\sa_count[19][38] , \sa_count[19].r.part1[6] );
tran (\sa_count[19][38] , \sa_count[19].f.upper[6] );
tran (\sa_count[19][37] , \sa_count[19].r.part1[5] );
tran (\sa_count[19][37] , \sa_count[19].f.upper[5] );
tran (\sa_count[19][36] , \sa_count[19].r.part1[4] );
tran (\sa_count[19][36] , \sa_count[19].f.upper[4] );
tran (\sa_count[19][35] , \sa_count[19].r.part1[3] );
tran (\sa_count[19][35] , \sa_count[19].f.upper[3] );
tran (\sa_count[19][34] , \sa_count[19].r.part1[2] );
tran (\sa_count[19][34] , \sa_count[19].f.upper[2] );
tran (\sa_count[19][33] , \sa_count[19].r.part1[1] );
tran (\sa_count[19][33] , \sa_count[19].f.upper[1] );
tran (\sa_count[19][32] , \sa_count[19].r.part1[0] );
tran (\sa_count[19][32] , \sa_count[19].f.upper[0] );
tran (\sa_count[19][31] , \sa_count[19].r.part0[31] );
tran (\sa_count[19][31] , \sa_count[19].f.lower[31] );
tran (\sa_count[19][30] , \sa_count[19].r.part0[30] );
tran (\sa_count[19][30] , \sa_count[19].f.lower[30] );
tran (\sa_count[19][29] , \sa_count[19].r.part0[29] );
tran (\sa_count[19][29] , \sa_count[19].f.lower[29] );
tran (\sa_count[19][28] , \sa_count[19].r.part0[28] );
tran (\sa_count[19][28] , \sa_count[19].f.lower[28] );
tran (\sa_count[19][27] , \sa_count[19].r.part0[27] );
tran (\sa_count[19][27] , \sa_count[19].f.lower[27] );
tran (\sa_count[19][26] , \sa_count[19].r.part0[26] );
tran (\sa_count[19][26] , \sa_count[19].f.lower[26] );
tran (\sa_count[19][25] , \sa_count[19].r.part0[25] );
tran (\sa_count[19][25] , \sa_count[19].f.lower[25] );
tran (\sa_count[19][24] , \sa_count[19].r.part0[24] );
tran (\sa_count[19][24] , \sa_count[19].f.lower[24] );
tran (\sa_count[19][23] , \sa_count[19].r.part0[23] );
tran (\sa_count[19][23] , \sa_count[19].f.lower[23] );
tran (\sa_count[19][22] , \sa_count[19].r.part0[22] );
tran (\sa_count[19][22] , \sa_count[19].f.lower[22] );
tran (\sa_count[19][21] , \sa_count[19].r.part0[21] );
tran (\sa_count[19][21] , \sa_count[19].f.lower[21] );
tran (\sa_count[19][20] , \sa_count[19].r.part0[20] );
tran (\sa_count[19][20] , \sa_count[19].f.lower[20] );
tran (\sa_count[19][19] , \sa_count[19].r.part0[19] );
tran (\sa_count[19][19] , \sa_count[19].f.lower[19] );
tran (\sa_count[19][18] , \sa_count[19].r.part0[18] );
tran (\sa_count[19][18] , \sa_count[19].f.lower[18] );
tran (\sa_count[19][17] , \sa_count[19].r.part0[17] );
tran (\sa_count[19][17] , \sa_count[19].f.lower[17] );
tran (\sa_count[19][16] , \sa_count[19].r.part0[16] );
tran (\sa_count[19][16] , \sa_count[19].f.lower[16] );
tran (\sa_count[19][15] , \sa_count[19].r.part0[15] );
tran (\sa_count[19][15] , \sa_count[19].f.lower[15] );
tran (\sa_count[19][14] , \sa_count[19].r.part0[14] );
tran (\sa_count[19][14] , \sa_count[19].f.lower[14] );
tran (\sa_count[19][13] , \sa_count[19].r.part0[13] );
tran (\sa_count[19][13] , \sa_count[19].f.lower[13] );
tran (\sa_count[19][12] , \sa_count[19].r.part0[12] );
tran (\sa_count[19][12] , \sa_count[19].f.lower[12] );
tran (\sa_count[19][11] , \sa_count[19].r.part0[11] );
tran (\sa_count[19][11] , \sa_count[19].f.lower[11] );
tran (\sa_count[19][10] , \sa_count[19].r.part0[10] );
tran (\sa_count[19][10] , \sa_count[19].f.lower[10] );
tran (\sa_count[19][9] , \sa_count[19].r.part0[9] );
tran (\sa_count[19][9] , \sa_count[19].f.lower[9] );
tran (\sa_count[19][8] , \sa_count[19].r.part0[8] );
tran (\sa_count[19][8] , \sa_count[19].f.lower[8] );
tran (\sa_count[19][7] , \sa_count[19].r.part0[7] );
tran (\sa_count[19][7] , \sa_count[19].f.lower[7] );
tran (\sa_count[19][6] , \sa_count[19].r.part0[6] );
tran (\sa_count[19][6] , \sa_count[19].f.lower[6] );
tran (\sa_count[19][5] , \sa_count[19].r.part0[5] );
tran (\sa_count[19][5] , \sa_count[19].f.lower[5] );
tran (\sa_count[19][4] , \sa_count[19].r.part0[4] );
tran (\sa_count[19][4] , \sa_count[19].f.lower[4] );
tran (\sa_count[19][3] , \sa_count[19].r.part0[3] );
tran (\sa_count[19][3] , \sa_count[19].f.lower[3] );
tran (\sa_count[19][2] , \sa_count[19].r.part0[2] );
tran (\sa_count[19][2] , \sa_count[19].f.lower[2] );
tran (\sa_count[19][1] , \sa_count[19].r.part0[1] );
tran (\sa_count[19][1] , \sa_count[19].f.lower[1] );
tran (\sa_count[19][0] , \sa_count[19].r.part0[0] );
tran (\sa_count[19][0] , \sa_count[19].f.lower[0] );
tran (\sa_count[18][63] , \sa_count[18].r.part1[31] );
tran (\sa_count[18][63] , \sa_count[18].f.unused[13] );
tran (\sa_count[18][62] , \sa_count[18].r.part1[30] );
tran (\sa_count[18][62] , \sa_count[18].f.unused[12] );
tran (\sa_count[18][61] , \sa_count[18].r.part1[29] );
tran (\sa_count[18][61] , \sa_count[18].f.unused[11] );
tran (\sa_count[18][60] , \sa_count[18].r.part1[28] );
tran (\sa_count[18][60] , \sa_count[18].f.unused[10] );
tran (\sa_count[18][59] , \sa_count[18].r.part1[27] );
tran (\sa_count[18][59] , \sa_count[18].f.unused[9] );
tran (\sa_count[18][58] , \sa_count[18].r.part1[26] );
tran (\sa_count[18][58] , \sa_count[18].f.unused[8] );
tran (\sa_count[18][57] , \sa_count[18].r.part1[25] );
tran (\sa_count[18][57] , \sa_count[18].f.unused[7] );
tran (\sa_count[18][56] , \sa_count[18].r.part1[24] );
tran (\sa_count[18][56] , \sa_count[18].f.unused[6] );
tran (\sa_count[18][55] , \sa_count[18].r.part1[23] );
tran (\sa_count[18][55] , \sa_count[18].f.unused[5] );
tran (\sa_count[18][54] , \sa_count[18].r.part1[22] );
tran (\sa_count[18][54] , \sa_count[18].f.unused[4] );
tran (\sa_count[18][53] , \sa_count[18].r.part1[21] );
tran (\sa_count[18][53] , \sa_count[18].f.unused[3] );
tran (\sa_count[18][52] , \sa_count[18].r.part1[20] );
tran (\sa_count[18][52] , \sa_count[18].f.unused[2] );
tran (\sa_count[18][51] , \sa_count[18].r.part1[19] );
tran (\sa_count[18][51] , \sa_count[18].f.unused[1] );
tran (\sa_count[18][50] , \sa_count[18].r.part1[18] );
tran (\sa_count[18][50] , \sa_count[18].f.unused[0] );
tran (\sa_count[18][49] , \sa_count[18].r.part1[17] );
tran (\sa_count[18][49] , \sa_count[18].f.upper[17] );
tran (\sa_count[18][48] , \sa_count[18].r.part1[16] );
tran (\sa_count[18][48] , \sa_count[18].f.upper[16] );
tran (\sa_count[18][47] , \sa_count[18].r.part1[15] );
tran (\sa_count[18][47] , \sa_count[18].f.upper[15] );
tran (\sa_count[18][46] , \sa_count[18].r.part1[14] );
tran (\sa_count[18][46] , \sa_count[18].f.upper[14] );
tran (\sa_count[18][45] , \sa_count[18].r.part1[13] );
tran (\sa_count[18][45] , \sa_count[18].f.upper[13] );
tran (\sa_count[18][44] , \sa_count[18].r.part1[12] );
tran (\sa_count[18][44] , \sa_count[18].f.upper[12] );
tran (\sa_count[18][43] , \sa_count[18].r.part1[11] );
tran (\sa_count[18][43] , \sa_count[18].f.upper[11] );
tran (\sa_count[18][42] , \sa_count[18].r.part1[10] );
tran (\sa_count[18][42] , \sa_count[18].f.upper[10] );
tran (\sa_count[18][41] , \sa_count[18].r.part1[9] );
tran (\sa_count[18][41] , \sa_count[18].f.upper[9] );
tran (\sa_count[18][40] , \sa_count[18].r.part1[8] );
tran (\sa_count[18][40] , \sa_count[18].f.upper[8] );
tran (\sa_count[18][39] , \sa_count[18].r.part1[7] );
tran (\sa_count[18][39] , \sa_count[18].f.upper[7] );
tran (\sa_count[18][38] , \sa_count[18].r.part1[6] );
tran (\sa_count[18][38] , \sa_count[18].f.upper[6] );
tran (\sa_count[18][37] , \sa_count[18].r.part1[5] );
tran (\sa_count[18][37] , \sa_count[18].f.upper[5] );
tran (\sa_count[18][36] , \sa_count[18].r.part1[4] );
tran (\sa_count[18][36] , \sa_count[18].f.upper[4] );
tran (\sa_count[18][35] , \sa_count[18].r.part1[3] );
tran (\sa_count[18][35] , \sa_count[18].f.upper[3] );
tran (\sa_count[18][34] , \sa_count[18].r.part1[2] );
tran (\sa_count[18][34] , \sa_count[18].f.upper[2] );
tran (\sa_count[18][33] , \sa_count[18].r.part1[1] );
tran (\sa_count[18][33] , \sa_count[18].f.upper[1] );
tran (\sa_count[18][32] , \sa_count[18].r.part1[0] );
tran (\sa_count[18][32] , \sa_count[18].f.upper[0] );
tran (\sa_count[18][31] , \sa_count[18].r.part0[31] );
tran (\sa_count[18][31] , \sa_count[18].f.lower[31] );
tran (\sa_count[18][30] , \sa_count[18].r.part0[30] );
tran (\sa_count[18][30] , \sa_count[18].f.lower[30] );
tran (\sa_count[18][29] , \sa_count[18].r.part0[29] );
tran (\sa_count[18][29] , \sa_count[18].f.lower[29] );
tran (\sa_count[18][28] , \sa_count[18].r.part0[28] );
tran (\sa_count[18][28] , \sa_count[18].f.lower[28] );
tran (\sa_count[18][27] , \sa_count[18].r.part0[27] );
tran (\sa_count[18][27] , \sa_count[18].f.lower[27] );
tran (\sa_count[18][26] , \sa_count[18].r.part0[26] );
tran (\sa_count[18][26] , \sa_count[18].f.lower[26] );
tran (\sa_count[18][25] , \sa_count[18].r.part0[25] );
tran (\sa_count[18][25] , \sa_count[18].f.lower[25] );
tran (\sa_count[18][24] , \sa_count[18].r.part0[24] );
tran (\sa_count[18][24] , \sa_count[18].f.lower[24] );
tran (\sa_count[18][23] , \sa_count[18].r.part0[23] );
tran (\sa_count[18][23] , \sa_count[18].f.lower[23] );
tran (\sa_count[18][22] , \sa_count[18].r.part0[22] );
tran (\sa_count[18][22] , \sa_count[18].f.lower[22] );
tran (\sa_count[18][21] , \sa_count[18].r.part0[21] );
tran (\sa_count[18][21] , \sa_count[18].f.lower[21] );
tran (\sa_count[18][20] , \sa_count[18].r.part0[20] );
tran (\sa_count[18][20] , \sa_count[18].f.lower[20] );
tran (\sa_count[18][19] , \sa_count[18].r.part0[19] );
tran (\sa_count[18][19] , \sa_count[18].f.lower[19] );
tran (\sa_count[18][18] , \sa_count[18].r.part0[18] );
tran (\sa_count[18][18] , \sa_count[18].f.lower[18] );
tran (\sa_count[18][17] , \sa_count[18].r.part0[17] );
tran (\sa_count[18][17] , \sa_count[18].f.lower[17] );
tran (\sa_count[18][16] , \sa_count[18].r.part0[16] );
tran (\sa_count[18][16] , \sa_count[18].f.lower[16] );
tran (\sa_count[18][15] , \sa_count[18].r.part0[15] );
tran (\sa_count[18][15] , \sa_count[18].f.lower[15] );
tran (\sa_count[18][14] , \sa_count[18].r.part0[14] );
tran (\sa_count[18][14] , \sa_count[18].f.lower[14] );
tran (\sa_count[18][13] , \sa_count[18].r.part0[13] );
tran (\sa_count[18][13] , \sa_count[18].f.lower[13] );
tran (\sa_count[18][12] , \sa_count[18].r.part0[12] );
tran (\sa_count[18][12] , \sa_count[18].f.lower[12] );
tran (\sa_count[18][11] , \sa_count[18].r.part0[11] );
tran (\sa_count[18][11] , \sa_count[18].f.lower[11] );
tran (\sa_count[18][10] , \sa_count[18].r.part0[10] );
tran (\sa_count[18][10] , \sa_count[18].f.lower[10] );
tran (\sa_count[18][9] , \sa_count[18].r.part0[9] );
tran (\sa_count[18][9] , \sa_count[18].f.lower[9] );
tran (\sa_count[18][8] , \sa_count[18].r.part0[8] );
tran (\sa_count[18][8] , \sa_count[18].f.lower[8] );
tran (\sa_count[18][7] , \sa_count[18].r.part0[7] );
tran (\sa_count[18][7] , \sa_count[18].f.lower[7] );
tran (\sa_count[18][6] , \sa_count[18].r.part0[6] );
tran (\sa_count[18][6] , \sa_count[18].f.lower[6] );
tran (\sa_count[18][5] , \sa_count[18].r.part0[5] );
tran (\sa_count[18][5] , \sa_count[18].f.lower[5] );
tran (\sa_count[18][4] , \sa_count[18].r.part0[4] );
tran (\sa_count[18][4] , \sa_count[18].f.lower[4] );
tran (\sa_count[18][3] , \sa_count[18].r.part0[3] );
tran (\sa_count[18][3] , \sa_count[18].f.lower[3] );
tran (\sa_count[18][2] , \sa_count[18].r.part0[2] );
tran (\sa_count[18][2] , \sa_count[18].f.lower[2] );
tran (\sa_count[18][1] , \sa_count[18].r.part0[1] );
tran (\sa_count[18][1] , \sa_count[18].f.lower[1] );
tran (\sa_count[18][0] , \sa_count[18].r.part0[0] );
tran (\sa_count[18][0] , \sa_count[18].f.lower[0] );
tran (\sa_count[17][63] , \sa_count[17].r.part1[31] );
tran (\sa_count[17][63] , \sa_count[17].f.unused[13] );
tran (\sa_count[17][62] , \sa_count[17].r.part1[30] );
tran (\sa_count[17][62] , \sa_count[17].f.unused[12] );
tran (\sa_count[17][61] , \sa_count[17].r.part1[29] );
tran (\sa_count[17][61] , \sa_count[17].f.unused[11] );
tran (\sa_count[17][60] , \sa_count[17].r.part1[28] );
tran (\sa_count[17][60] , \sa_count[17].f.unused[10] );
tran (\sa_count[17][59] , \sa_count[17].r.part1[27] );
tran (\sa_count[17][59] , \sa_count[17].f.unused[9] );
tran (\sa_count[17][58] , \sa_count[17].r.part1[26] );
tran (\sa_count[17][58] , \sa_count[17].f.unused[8] );
tran (\sa_count[17][57] , \sa_count[17].r.part1[25] );
tran (\sa_count[17][57] , \sa_count[17].f.unused[7] );
tran (\sa_count[17][56] , \sa_count[17].r.part1[24] );
tran (\sa_count[17][56] , \sa_count[17].f.unused[6] );
tran (\sa_count[17][55] , \sa_count[17].r.part1[23] );
tran (\sa_count[17][55] , \sa_count[17].f.unused[5] );
tran (\sa_count[17][54] , \sa_count[17].r.part1[22] );
tran (\sa_count[17][54] , \sa_count[17].f.unused[4] );
tran (\sa_count[17][53] , \sa_count[17].r.part1[21] );
tran (\sa_count[17][53] , \sa_count[17].f.unused[3] );
tran (\sa_count[17][52] , \sa_count[17].r.part1[20] );
tran (\sa_count[17][52] , \sa_count[17].f.unused[2] );
tran (\sa_count[17][51] , \sa_count[17].r.part1[19] );
tran (\sa_count[17][51] , \sa_count[17].f.unused[1] );
tran (\sa_count[17][50] , \sa_count[17].r.part1[18] );
tran (\sa_count[17][50] , \sa_count[17].f.unused[0] );
tran (\sa_count[17][49] , \sa_count[17].r.part1[17] );
tran (\sa_count[17][49] , \sa_count[17].f.upper[17] );
tran (\sa_count[17][48] , \sa_count[17].r.part1[16] );
tran (\sa_count[17][48] , \sa_count[17].f.upper[16] );
tran (\sa_count[17][47] , \sa_count[17].r.part1[15] );
tran (\sa_count[17][47] , \sa_count[17].f.upper[15] );
tran (\sa_count[17][46] , \sa_count[17].r.part1[14] );
tran (\sa_count[17][46] , \sa_count[17].f.upper[14] );
tran (\sa_count[17][45] , \sa_count[17].r.part1[13] );
tran (\sa_count[17][45] , \sa_count[17].f.upper[13] );
tran (\sa_count[17][44] , \sa_count[17].r.part1[12] );
tran (\sa_count[17][44] , \sa_count[17].f.upper[12] );
tran (\sa_count[17][43] , \sa_count[17].r.part1[11] );
tran (\sa_count[17][43] , \sa_count[17].f.upper[11] );
tran (\sa_count[17][42] , \sa_count[17].r.part1[10] );
tran (\sa_count[17][42] , \sa_count[17].f.upper[10] );
tran (\sa_count[17][41] , \sa_count[17].r.part1[9] );
tran (\sa_count[17][41] , \sa_count[17].f.upper[9] );
tran (\sa_count[17][40] , \sa_count[17].r.part1[8] );
tran (\sa_count[17][40] , \sa_count[17].f.upper[8] );
tran (\sa_count[17][39] , \sa_count[17].r.part1[7] );
tran (\sa_count[17][39] , \sa_count[17].f.upper[7] );
tran (\sa_count[17][38] , \sa_count[17].r.part1[6] );
tran (\sa_count[17][38] , \sa_count[17].f.upper[6] );
tran (\sa_count[17][37] , \sa_count[17].r.part1[5] );
tran (\sa_count[17][37] , \sa_count[17].f.upper[5] );
tran (\sa_count[17][36] , \sa_count[17].r.part1[4] );
tran (\sa_count[17][36] , \sa_count[17].f.upper[4] );
tran (\sa_count[17][35] , \sa_count[17].r.part1[3] );
tran (\sa_count[17][35] , \sa_count[17].f.upper[3] );
tran (\sa_count[17][34] , \sa_count[17].r.part1[2] );
tran (\sa_count[17][34] , \sa_count[17].f.upper[2] );
tran (\sa_count[17][33] , \sa_count[17].r.part1[1] );
tran (\sa_count[17][33] , \sa_count[17].f.upper[1] );
tran (\sa_count[17][32] , \sa_count[17].r.part1[0] );
tran (\sa_count[17][32] , \sa_count[17].f.upper[0] );
tran (\sa_count[17][31] , \sa_count[17].r.part0[31] );
tran (\sa_count[17][31] , \sa_count[17].f.lower[31] );
tran (\sa_count[17][30] , \sa_count[17].r.part0[30] );
tran (\sa_count[17][30] , \sa_count[17].f.lower[30] );
tran (\sa_count[17][29] , \sa_count[17].r.part0[29] );
tran (\sa_count[17][29] , \sa_count[17].f.lower[29] );
tran (\sa_count[17][28] , \sa_count[17].r.part0[28] );
tran (\sa_count[17][28] , \sa_count[17].f.lower[28] );
tran (\sa_count[17][27] , \sa_count[17].r.part0[27] );
tran (\sa_count[17][27] , \sa_count[17].f.lower[27] );
tran (\sa_count[17][26] , \sa_count[17].r.part0[26] );
tran (\sa_count[17][26] , \sa_count[17].f.lower[26] );
tran (\sa_count[17][25] , \sa_count[17].r.part0[25] );
tran (\sa_count[17][25] , \sa_count[17].f.lower[25] );
tran (\sa_count[17][24] , \sa_count[17].r.part0[24] );
tran (\sa_count[17][24] , \sa_count[17].f.lower[24] );
tran (\sa_count[17][23] , \sa_count[17].r.part0[23] );
tran (\sa_count[17][23] , \sa_count[17].f.lower[23] );
tran (\sa_count[17][22] , \sa_count[17].r.part0[22] );
tran (\sa_count[17][22] , \sa_count[17].f.lower[22] );
tran (\sa_count[17][21] , \sa_count[17].r.part0[21] );
tran (\sa_count[17][21] , \sa_count[17].f.lower[21] );
tran (\sa_count[17][20] , \sa_count[17].r.part0[20] );
tran (\sa_count[17][20] , \sa_count[17].f.lower[20] );
tran (\sa_count[17][19] , \sa_count[17].r.part0[19] );
tran (\sa_count[17][19] , \sa_count[17].f.lower[19] );
tran (\sa_count[17][18] , \sa_count[17].r.part0[18] );
tran (\sa_count[17][18] , \sa_count[17].f.lower[18] );
tran (\sa_count[17][17] , \sa_count[17].r.part0[17] );
tran (\sa_count[17][17] , \sa_count[17].f.lower[17] );
tran (\sa_count[17][16] , \sa_count[17].r.part0[16] );
tran (\sa_count[17][16] , \sa_count[17].f.lower[16] );
tran (\sa_count[17][15] , \sa_count[17].r.part0[15] );
tran (\sa_count[17][15] , \sa_count[17].f.lower[15] );
tran (\sa_count[17][14] , \sa_count[17].r.part0[14] );
tran (\sa_count[17][14] , \sa_count[17].f.lower[14] );
tran (\sa_count[17][13] , \sa_count[17].r.part0[13] );
tran (\sa_count[17][13] , \sa_count[17].f.lower[13] );
tran (\sa_count[17][12] , \sa_count[17].r.part0[12] );
tran (\sa_count[17][12] , \sa_count[17].f.lower[12] );
tran (\sa_count[17][11] , \sa_count[17].r.part0[11] );
tran (\sa_count[17][11] , \sa_count[17].f.lower[11] );
tran (\sa_count[17][10] , \sa_count[17].r.part0[10] );
tran (\sa_count[17][10] , \sa_count[17].f.lower[10] );
tran (\sa_count[17][9] , \sa_count[17].r.part0[9] );
tran (\sa_count[17][9] , \sa_count[17].f.lower[9] );
tran (\sa_count[17][8] , \sa_count[17].r.part0[8] );
tran (\sa_count[17][8] , \sa_count[17].f.lower[8] );
tran (\sa_count[17][7] , \sa_count[17].r.part0[7] );
tran (\sa_count[17][7] , \sa_count[17].f.lower[7] );
tran (\sa_count[17][6] , \sa_count[17].r.part0[6] );
tran (\sa_count[17][6] , \sa_count[17].f.lower[6] );
tran (\sa_count[17][5] , \sa_count[17].r.part0[5] );
tran (\sa_count[17][5] , \sa_count[17].f.lower[5] );
tran (\sa_count[17][4] , \sa_count[17].r.part0[4] );
tran (\sa_count[17][4] , \sa_count[17].f.lower[4] );
tran (\sa_count[17][3] , \sa_count[17].r.part0[3] );
tran (\sa_count[17][3] , \sa_count[17].f.lower[3] );
tran (\sa_count[17][2] , \sa_count[17].r.part0[2] );
tran (\sa_count[17][2] , \sa_count[17].f.lower[2] );
tran (\sa_count[17][1] , \sa_count[17].r.part0[1] );
tran (\sa_count[17][1] , \sa_count[17].f.lower[1] );
tran (\sa_count[17][0] , \sa_count[17].r.part0[0] );
tran (\sa_count[17][0] , \sa_count[17].f.lower[0] );
tran (\sa_count[16][63] , \sa_count[16].r.part1[31] );
tran (\sa_count[16][63] , \sa_count[16].f.unused[13] );
tran (\sa_count[16][62] , \sa_count[16].r.part1[30] );
tran (\sa_count[16][62] , \sa_count[16].f.unused[12] );
tran (\sa_count[16][61] , \sa_count[16].r.part1[29] );
tran (\sa_count[16][61] , \sa_count[16].f.unused[11] );
tran (\sa_count[16][60] , \sa_count[16].r.part1[28] );
tran (\sa_count[16][60] , \sa_count[16].f.unused[10] );
tran (\sa_count[16][59] , \sa_count[16].r.part1[27] );
tran (\sa_count[16][59] , \sa_count[16].f.unused[9] );
tran (\sa_count[16][58] , \sa_count[16].r.part1[26] );
tran (\sa_count[16][58] , \sa_count[16].f.unused[8] );
tran (\sa_count[16][57] , \sa_count[16].r.part1[25] );
tran (\sa_count[16][57] , \sa_count[16].f.unused[7] );
tran (\sa_count[16][56] , \sa_count[16].r.part1[24] );
tran (\sa_count[16][56] , \sa_count[16].f.unused[6] );
tran (\sa_count[16][55] , \sa_count[16].r.part1[23] );
tran (\sa_count[16][55] , \sa_count[16].f.unused[5] );
tran (\sa_count[16][54] , \sa_count[16].r.part1[22] );
tran (\sa_count[16][54] , \sa_count[16].f.unused[4] );
tran (\sa_count[16][53] , \sa_count[16].r.part1[21] );
tran (\sa_count[16][53] , \sa_count[16].f.unused[3] );
tran (\sa_count[16][52] , \sa_count[16].r.part1[20] );
tran (\sa_count[16][52] , \sa_count[16].f.unused[2] );
tran (\sa_count[16][51] , \sa_count[16].r.part1[19] );
tran (\sa_count[16][51] , \sa_count[16].f.unused[1] );
tran (\sa_count[16][50] , \sa_count[16].r.part1[18] );
tran (\sa_count[16][50] , \sa_count[16].f.unused[0] );
tran (\sa_count[16][49] , \sa_count[16].r.part1[17] );
tran (\sa_count[16][49] , \sa_count[16].f.upper[17] );
tran (\sa_count[16][48] , \sa_count[16].r.part1[16] );
tran (\sa_count[16][48] , \sa_count[16].f.upper[16] );
tran (\sa_count[16][47] , \sa_count[16].r.part1[15] );
tran (\sa_count[16][47] , \sa_count[16].f.upper[15] );
tran (\sa_count[16][46] , \sa_count[16].r.part1[14] );
tran (\sa_count[16][46] , \sa_count[16].f.upper[14] );
tran (\sa_count[16][45] , \sa_count[16].r.part1[13] );
tran (\sa_count[16][45] , \sa_count[16].f.upper[13] );
tran (\sa_count[16][44] , \sa_count[16].r.part1[12] );
tran (\sa_count[16][44] , \sa_count[16].f.upper[12] );
tran (\sa_count[16][43] , \sa_count[16].r.part1[11] );
tran (\sa_count[16][43] , \sa_count[16].f.upper[11] );
tran (\sa_count[16][42] , \sa_count[16].r.part1[10] );
tran (\sa_count[16][42] , \sa_count[16].f.upper[10] );
tran (\sa_count[16][41] , \sa_count[16].r.part1[9] );
tran (\sa_count[16][41] , \sa_count[16].f.upper[9] );
tran (\sa_count[16][40] , \sa_count[16].r.part1[8] );
tran (\sa_count[16][40] , \sa_count[16].f.upper[8] );
tran (\sa_count[16][39] , \sa_count[16].r.part1[7] );
tran (\sa_count[16][39] , \sa_count[16].f.upper[7] );
tran (\sa_count[16][38] , \sa_count[16].r.part1[6] );
tran (\sa_count[16][38] , \sa_count[16].f.upper[6] );
tran (\sa_count[16][37] , \sa_count[16].r.part1[5] );
tran (\sa_count[16][37] , \sa_count[16].f.upper[5] );
tran (\sa_count[16][36] , \sa_count[16].r.part1[4] );
tran (\sa_count[16][36] , \sa_count[16].f.upper[4] );
tran (\sa_count[16][35] , \sa_count[16].r.part1[3] );
tran (\sa_count[16][35] , \sa_count[16].f.upper[3] );
tran (\sa_count[16][34] , \sa_count[16].r.part1[2] );
tran (\sa_count[16][34] , \sa_count[16].f.upper[2] );
tran (\sa_count[16][33] , \sa_count[16].r.part1[1] );
tran (\sa_count[16][33] , \sa_count[16].f.upper[1] );
tran (\sa_count[16][32] , \sa_count[16].r.part1[0] );
tran (\sa_count[16][32] , \sa_count[16].f.upper[0] );
tran (\sa_count[16][31] , \sa_count[16].r.part0[31] );
tran (\sa_count[16][31] , \sa_count[16].f.lower[31] );
tran (\sa_count[16][30] , \sa_count[16].r.part0[30] );
tran (\sa_count[16][30] , \sa_count[16].f.lower[30] );
tran (\sa_count[16][29] , \sa_count[16].r.part0[29] );
tran (\sa_count[16][29] , \sa_count[16].f.lower[29] );
tran (\sa_count[16][28] , \sa_count[16].r.part0[28] );
tran (\sa_count[16][28] , \sa_count[16].f.lower[28] );
tran (\sa_count[16][27] , \sa_count[16].r.part0[27] );
tran (\sa_count[16][27] , \sa_count[16].f.lower[27] );
tran (\sa_count[16][26] , \sa_count[16].r.part0[26] );
tran (\sa_count[16][26] , \sa_count[16].f.lower[26] );
tran (\sa_count[16][25] , \sa_count[16].r.part0[25] );
tran (\sa_count[16][25] , \sa_count[16].f.lower[25] );
tran (\sa_count[16][24] , \sa_count[16].r.part0[24] );
tran (\sa_count[16][24] , \sa_count[16].f.lower[24] );
tran (\sa_count[16][23] , \sa_count[16].r.part0[23] );
tran (\sa_count[16][23] , \sa_count[16].f.lower[23] );
tran (\sa_count[16][22] , \sa_count[16].r.part0[22] );
tran (\sa_count[16][22] , \sa_count[16].f.lower[22] );
tran (\sa_count[16][21] , \sa_count[16].r.part0[21] );
tran (\sa_count[16][21] , \sa_count[16].f.lower[21] );
tran (\sa_count[16][20] , \sa_count[16].r.part0[20] );
tran (\sa_count[16][20] , \sa_count[16].f.lower[20] );
tran (\sa_count[16][19] , \sa_count[16].r.part0[19] );
tran (\sa_count[16][19] , \sa_count[16].f.lower[19] );
tran (\sa_count[16][18] , \sa_count[16].r.part0[18] );
tran (\sa_count[16][18] , \sa_count[16].f.lower[18] );
tran (\sa_count[16][17] , \sa_count[16].r.part0[17] );
tran (\sa_count[16][17] , \sa_count[16].f.lower[17] );
tran (\sa_count[16][16] , \sa_count[16].r.part0[16] );
tran (\sa_count[16][16] , \sa_count[16].f.lower[16] );
tran (\sa_count[16][15] , \sa_count[16].r.part0[15] );
tran (\sa_count[16][15] , \sa_count[16].f.lower[15] );
tran (\sa_count[16][14] , \sa_count[16].r.part0[14] );
tran (\sa_count[16][14] , \sa_count[16].f.lower[14] );
tran (\sa_count[16][13] , \sa_count[16].r.part0[13] );
tran (\sa_count[16][13] , \sa_count[16].f.lower[13] );
tran (\sa_count[16][12] , \sa_count[16].r.part0[12] );
tran (\sa_count[16][12] , \sa_count[16].f.lower[12] );
tran (\sa_count[16][11] , \sa_count[16].r.part0[11] );
tran (\sa_count[16][11] , \sa_count[16].f.lower[11] );
tran (\sa_count[16][10] , \sa_count[16].r.part0[10] );
tran (\sa_count[16][10] , \sa_count[16].f.lower[10] );
tran (\sa_count[16][9] , \sa_count[16].r.part0[9] );
tran (\sa_count[16][9] , \sa_count[16].f.lower[9] );
tran (\sa_count[16][8] , \sa_count[16].r.part0[8] );
tran (\sa_count[16][8] , \sa_count[16].f.lower[8] );
tran (\sa_count[16][7] , \sa_count[16].r.part0[7] );
tran (\sa_count[16][7] , \sa_count[16].f.lower[7] );
tran (\sa_count[16][6] , \sa_count[16].r.part0[6] );
tran (\sa_count[16][6] , \sa_count[16].f.lower[6] );
tran (\sa_count[16][5] , \sa_count[16].r.part0[5] );
tran (\sa_count[16][5] , \sa_count[16].f.lower[5] );
tran (\sa_count[16][4] , \sa_count[16].r.part0[4] );
tran (\sa_count[16][4] , \sa_count[16].f.lower[4] );
tran (\sa_count[16][3] , \sa_count[16].r.part0[3] );
tran (\sa_count[16][3] , \sa_count[16].f.lower[3] );
tran (\sa_count[16][2] , \sa_count[16].r.part0[2] );
tran (\sa_count[16][2] , \sa_count[16].f.lower[2] );
tran (\sa_count[16][1] , \sa_count[16].r.part0[1] );
tran (\sa_count[16][1] , \sa_count[16].f.lower[1] );
tran (\sa_count[16][0] , \sa_count[16].r.part0[0] );
tran (\sa_count[16][0] , \sa_count[16].f.lower[0] );
tran (\sa_count[15][63] , \sa_count[15].r.part1[31] );
tran (\sa_count[15][63] , \sa_count[15].f.unused[13] );
tran (\sa_count[15][62] , \sa_count[15].r.part1[30] );
tran (\sa_count[15][62] , \sa_count[15].f.unused[12] );
tran (\sa_count[15][61] , \sa_count[15].r.part1[29] );
tran (\sa_count[15][61] , \sa_count[15].f.unused[11] );
tran (\sa_count[15][60] , \sa_count[15].r.part1[28] );
tran (\sa_count[15][60] , \sa_count[15].f.unused[10] );
tran (\sa_count[15][59] , \sa_count[15].r.part1[27] );
tran (\sa_count[15][59] , \sa_count[15].f.unused[9] );
tran (\sa_count[15][58] , \sa_count[15].r.part1[26] );
tran (\sa_count[15][58] , \sa_count[15].f.unused[8] );
tran (\sa_count[15][57] , \sa_count[15].r.part1[25] );
tran (\sa_count[15][57] , \sa_count[15].f.unused[7] );
tran (\sa_count[15][56] , \sa_count[15].r.part1[24] );
tran (\sa_count[15][56] , \sa_count[15].f.unused[6] );
tran (\sa_count[15][55] , \sa_count[15].r.part1[23] );
tran (\sa_count[15][55] , \sa_count[15].f.unused[5] );
tran (\sa_count[15][54] , \sa_count[15].r.part1[22] );
tran (\sa_count[15][54] , \sa_count[15].f.unused[4] );
tran (\sa_count[15][53] , \sa_count[15].r.part1[21] );
tran (\sa_count[15][53] , \sa_count[15].f.unused[3] );
tran (\sa_count[15][52] , \sa_count[15].r.part1[20] );
tran (\sa_count[15][52] , \sa_count[15].f.unused[2] );
tran (\sa_count[15][51] , \sa_count[15].r.part1[19] );
tran (\sa_count[15][51] , \sa_count[15].f.unused[1] );
tran (\sa_count[15][50] , \sa_count[15].r.part1[18] );
tran (\sa_count[15][50] , \sa_count[15].f.unused[0] );
tran (\sa_count[15][49] , \sa_count[15].r.part1[17] );
tran (\sa_count[15][49] , \sa_count[15].f.upper[17] );
tran (\sa_count[15][48] , \sa_count[15].r.part1[16] );
tran (\sa_count[15][48] , \sa_count[15].f.upper[16] );
tran (\sa_count[15][47] , \sa_count[15].r.part1[15] );
tran (\sa_count[15][47] , \sa_count[15].f.upper[15] );
tran (\sa_count[15][46] , \sa_count[15].r.part1[14] );
tran (\sa_count[15][46] , \sa_count[15].f.upper[14] );
tran (\sa_count[15][45] , \sa_count[15].r.part1[13] );
tran (\sa_count[15][45] , \sa_count[15].f.upper[13] );
tran (\sa_count[15][44] , \sa_count[15].r.part1[12] );
tran (\sa_count[15][44] , \sa_count[15].f.upper[12] );
tran (\sa_count[15][43] , \sa_count[15].r.part1[11] );
tran (\sa_count[15][43] , \sa_count[15].f.upper[11] );
tran (\sa_count[15][42] , \sa_count[15].r.part1[10] );
tran (\sa_count[15][42] , \sa_count[15].f.upper[10] );
tran (\sa_count[15][41] , \sa_count[15].r.part1[9] );
tran (\sa_count[15][41] , \sa_count[15].f.upper[9] );
tran (\sa_count[15][40] , \sa_count[15].r.part1[8] );
tran (\sa_count[15][40] , \sa_count[15].f.upper[8] );
tran (\sa_count[15][39] , \sa_count[15].r.part1[7] );
tran (\sa_count[15][39] , \sa_count[15].f.upper[7] );
tran (\sa_count[15][38] , \sa_count[15].r.part1[6] );
tran (\sa_count[15][38] , \sa_count[15].f.upper[6] );
tran (\sa_count[15][37] , \sa_count[15].r.part1[5] );
tran (\sa_count[15][37] , \sa_count[15].f.upper[5] );
tran (\sa_count[15][36] , \sa_count[15].r.part1[4] );
tran (\sa_count[15][36] , \sa_count[15].f.upper[4] );
tran (\sa_count[15][35] , \sa_count[15].r.part1[3] );
tran (\sa_count[15][35] , \sa_count[15].f.upper[3] );
tran (\sa_count[15][34] , \sa_count[15].r.part1[2] );
tran (\sa_count[15][34] , \sa_count[15].f.upper[2] );
tran (\sa_count[15][33] , \sa_count[15].r.part1[1] );
tran (\sa_count[15][33] , \sa_count[15].f.upper[1] );
tran (\sa_count[15][32] , \sa_count[15].r.part1[0] );
tran (\sa_count[15][32] , \sa_count[15].f.upper[0] );
tran (\sa_count[15][31] , \sa_count[15].r.part0[31] );
tran (\sa_count[15][31] , \sa_count[15].f.lower[31] );
tran (\sa_count[15][30] , \sa_count[15].r.part0[30] );
tran (\sa_count[15][30] , \sa_count[15].f.lower[30] );
tran (\sa_count[15][29] , \sa_count[15].r.part0[29] );
tran (\sa_count[15][29] , \sa_count[15].f.lower[29] );
tran (\sa_count[15][28] , \sa_count[15].r.part0[28] );
tran (\sa_count[15][28] , \sa_count[15].f.lower[28] );
tran (\sa_count[15][27] , \sa_count[15].r.part0[27] );
tran (\sa_count[15][27] , \sa_count[15].f.lower[27] );
tran (\sa_count[15][26] , \sa_count[15].r.part0[26] );
tran (\sa_count[15][26] , \sa_count[15].f.lower[26] );
tran (\sa_count[15][25] , \sa_count[15].r.part0[25] );
tran (\sa_count[15][25] , \sa_count[15].f.lower[25] );
tran (\sa_count[15][24] , \sa_count[15].r.part0[24] );
tran (\sa_count[15][24] , \sa_count[15].f.lower[24] );
tran (\sa_count[15][23] , \sa_count[15].r.part0[23] );
tran (\sa_count[15][23] , \sa_count[15].f.lower[23] );
tran (\sa_count[15][22] , \sa_count[15].r.part0[22] );
tran (\sa_count[15][22] , \sa_count[15].f.lower[22] );
tran (\sa_count[15][21] , \sa_count[15].r.part0[21] );
tran (\sa_count[15][21] , \sa_count[15].f.lower[21] );
tran (\sa_count[15][20] , \sa_count[15].r.part0[20] );
tran (\sa_count[15][20] , \sa_count[15].f.lower[20] );
tran (\sa_count[15][19] , \sa_count[15].r.part0[19] );
tran (\sa_count[15][19] , \sa_count[15].f.lower[19] );
tran (\sa_count[15][18] , \sa_count[15].r.part0[18] );
tran (\sa_count[15][18] , \sa_count[15].f.lower[18] );
tran (\sa_count[15][17] , \sa_count[15].r.part0[17] );
tran (\sa_count[15][17] , \sa_count[15].f.lower[17] );
tran (\sa_count[15][16] , \sa_count[15].r.part0[16] );
tran (\sa_count[15][16] , \sa_count[15].f.lower[16] );
tran (\sa_count[15][15] , \sa_count[15].r.part0[15] );
tran (\sa_count[15][15] , \sa_count[15].f.lower[15] );
tran (\sa_count[15][14] , \sa_count[15].r.part0[14] );
tran (\sa_count[15][14] , \sa_count[15].f.lower[14] );
tran (\sa_count[15][13] , \sa_count[15].r.part0[13] );
tran (\sa_count[15][13] , \sa_count[15].f.lower[13] );
tran (\sa_count[15][12] , \sa_count[15].r.part0[12] );
tran (\sa_count[15][12] , \sa_count[15].f.lower[12] );
tran (\sa_count[15][11] , \sa_count[15].r.part0[11] );
tran (\sa_count[15][11] , \sa_count[15].f.lower[11] );
tran (\sa_count[15][10] , \sa_count[15].r.part0[10] );
tran (\sa_count[15][10] , \sa_count[15].f.lower[10] );
tran (\sa_count[15][9] , \sa_count[15].r.part0[9] );
tran (\sa_count[15][9] , \sa_count[15].f.lower[9] );
tran (\sa_count[15][8] , \sa_count[15].r.part0[8] );
tran (\sa_count[15][8] , \sa_count[15].f.lower[8] );
tran (\sa_count[15][7] , \sa_count[15].r.part0[7] );
tran (\sa_count[15][7] , \sa_count[15].f.lower[7] );
tran (\sa_count[15][6] , \sa_count[15].r.part0[6] );
tran (\sa_count[15][6] , \sa_count[15].f.lower[6] );
tran (\sa_count[15][5] , \sa_count[15].r.part0[5] );
tran (\sa_count[15][5] , \sa_count[15].f.lower[5] );
tran (\sa_count[15][4] , \sa_count[15].r.part0[4] );
tran (\sa_count[15][4] , \sa_count[15].f.lower[4] );
tran (\sa_count[15][3] , \sa_count[15].r.part0[3] );
tran (\sa_count[15][3] , \sa_count[15].f.lower[3] );
tran (\sa_count[15][2] , \sa_count[15].r.part0[2] );
tran (\sa_count[15][2] , \sa_count[15].f.lower[2] );
tran (\sa_count[15][1] , \sa_count[15].r.part0[1] );
tran (\sa_count[15][1] , \sa_count[15].f.lower[1] );
tran (\sa_count[15][0] , \sa_count[15].r.part0[0] );
tran (\sa_count[15][0] , \sa_count[15].f.lower[0] );
tran (\sa_count[14][63] , \sa_count[14].r.part1[31] );
tran (\sa_count[14][63] , \sa_count[14].f.unused[13] );
tran (\sa_count[14][62] , \sa_count[14].r.part1[30] );
tran (\sa_count[14][62] , \sa_count[14].f.unused[12] );
tran (\sa_count[14][61] , \sa_count[14].r.part1[29] );
tran (\sa_count[14][61] , \sa_count[14].f.unused[11] );
tran (\sa_count[14][60] , \sa_count[14].r.part1[28] );
tran (\sa_count[14][60] , \sa_count[14].f.unused[10] );
tran (\sa_count[14][59] , \sa_count[14].r.part1[27] );
tran (\sa_count[14][59] , \sa_count[14].f.unused[9] );
tran (\sa_count[14][58] , \sa_count[14].r.part1[26] );
tran (\sa_count[14][58] , \sa_count[14].f.unused[8] );
tran (\sa_count[14][57] , \sa_count[14].r.part1[25] );
tran (\sa_count[14][57] , \sa_count[14].f.unused[7] );
tran (\sa_count[14][56] , \sa_count[14].r.part1[24] );
tran (\sa_count[14][56] , \sa_count[14].f.unused[6] );
tran (\sa_count[14][55] , \sa_count[14].r.part1[23] );
tran (\sa_count[14][55] , \sa_count[14].f.unused[5] );
tran (\sa_count[14][54] , \sa_count[14].r.part1[22] );
tran (\sa_count[14][54] , \sa_count[14].f.unused[4] );
tran (\sa_count[14][53] , \sa_count[14].r.part1[21] );
tran (\sa_count[14][53] , \sa_count[14].f.unused[3] );
tran (\sa_count[14][52] , \sa_count[14].r.part1[20] );
tran (\sa_count[14][52] , \sa_count[14].f.unused[2] );
tran (\sa_count[14][51] , \sa_count[14].r.part1[19] );
tran (\sa_count[14][51] , \sa_count[14].f.unused[1] );
tran (\sa_count[14][50] , \sa_count[14].r.part1[18] );
tran (\sa_count[14][50] , \sa_count[14].f.unused[0] );
tran (\sa_count[14][49] , \sa_count[14].r.part1[17] );
tran (\sa_count[14][49] , \sa_count[14].f.upper[17] );
tran (\sa_count[14][48] , \sa_count[14].r.part1[16] );
tran (\sa_count[14][48] , \sa_count[14].f.upper[16] );
tran (\sa_count[14][47] , \sa_count[14].r.part1[15] );
tran (\sa_count[14][47] , \sa_count[14].f.upper[15] );
tran (\sa_count[14][46] , \sa_count[14].r.part1[14] );
tran (\sa_count[14][46] , \sa_count[14].f.upper[14] );
tran (\sa_count[14][45] , \sa_count[14].r.part1[13] );
tran (\sa_count[14][45] , \sa_count[14].f.upper[13] );
tran (\sa_count[14][44] , \sa_count[14].r.part1[12] );
tran (\sa_count[14][44] , \sa_count[14].f.upper[12] );
tran (\sa_count[14][43] , \sa_count[14].r.part1[11] );
tran (\sa_count[14][43] , \sa_count[14].f.upper[11] );
tran (\sa_count[14][42] , \sa_count[14].r.part1[10] );
tran (\sa_count[14][42] , \sa_count[14].f.upper[10] );
tran (\sa_count[14][41] , \sa_count[14].r.part1[9] );
tran (\sa_count[14][41] , \sa_count[14].f.upper[9] );
tran (\sa_count[14][40] , \sa_count[14].r.part1[8] );
tran (\sa_count[14][40] , \sa_count[14].f.upper[8] );
tran (\sa_count[14][39] , \sa_count[14].r.part1[7] );
tran (\sa_count[14][39] , \sa_count[14].f.upper[7] );
tran (\sa_count[14][38] , \sa_count[14].r.part1[6] );
tran (\sa_count[14][38] , \sa_count[14].f.upper[6] );
tran (\sa_count[14][37] , \sa_count[14].r.part1[5] );
tran (\sa_count[14][37] , \sa_count[14].f.upper[5] );
tran (\sa_count[14][36] , \sa_count[14].r.part1[4] );
tran (\sa_count[14][36] , \sa_count[14].f.upper[4] );
tran (\sa_count[14][35] , \sa_count[14].r.part1[3] );
tran (\sa_count[14][35] , \sa_count[14].f.upper[3] );
tran (\sa_count[14][34] , \sa_count[14].r.part1[2] );
tran (\sa_count[14][34] , \sa_count[14].f.upper[2] );
tran (\sa_count[14][33] , \sa_count[14].r.part1[1] );
tran (\sa_count[14][33] , \sa_count[14].f.upper[1] );
tran (\sa_count[14][32] , \sa_count[14].r.part1[0] );
tran (\sa_count[14][32] , \sa_count[14].f.upper[0] );
tran (\sa_count[14][31] , \sa_count[14].r.part0[31] );
tran (\sa_count[14][31] , \sa_count[14].f.lower[31] );
tran (\sa_count[14][30] , \sa_count[14].r.part0[30] );
tran (\sa_count[14][30] , \sa_count[14].f.lower[30] );
tran (\sa_count[14][29] , \sa_count[14].r.part0[29] );
tran (\sa_count[14][29] , \sa_count[14].f.lower[29] );
tran (\sa_count[14][28] , \sa_count[14].r.part0[28] );
tran (\sa_count[14][28] , \sa_count[14].f.lower[28] );
tran (\sa_count[14][27] , \sa_count[14].r.part0[27] );
tran (\sa_count[14][27] , \sa_count[14].f.lower[27] );
tran (\sa_count[14][26] , \sa_count[14].r.part0[26] );
tran (\sa_count[14][26] , \sa_count[14].f.lower[26] );
tran (\sa_count[14][25] , \sa_count[14].r.part0[25] );
tran (\sa_count[14][25] , \sa_count[14].f.lower[25] );
tran (\sa_count[14][24] , \sa_count[14].r.part0[24] );
tran (\sa_count[14][24] , \sa_count[14].f.lower[24] );
tran (\sa_count[14][23] , \sa_count[14].r.part0[23] );
tran (\sa_count[14][23] , \sa_count[14].f.lower[23] );
tran (\sa_count[14][22] , \sa_count[14].r.part0[22] );
tran (\sa_count[14][22] , \sa_count[14].f.lower[22] );
tran (\sa_count[14][21] , \sa_count[14].r.part0[21] );
tran (\sa_count[14][21] , \sa_count[14].f.lower[21] );
tran (\sa_count[14][20] , \sa_count[14].r.part0[20] );
tran (\sa_count[14][20] , \sa_count[14].f.lower[20] );
tran (\sa_count[14][19] , \sa_count[14].r.part0[19] );
tran (\sa_count[14][19] , \sa_count[14].f.lower[19] );
tran (\sa_count[14][18] , \sa_count[14].r.part0[18] );
tran (\sa_count[14][18] , \sa_count[14].f.lower[18] );
tran (\sa_count[14][17] , \sa_count[14].r.part0[17] );
tran (\sa_count[14][17] , \sa_count[14].f.lower[17] );
tran (\sa_count[14][16] , \sa_count[14].r.part0[16] );
tran (\sa_count[14][16] , \sa_count[14].f.lower[16] );
tran (\sa_count[14][15] , \sa_count[14].r.part0[15] );
tran (\sa_count[14][15] , \sa_count[14].f.lower[15] );
tran (\sa_count[14][14] , \sa_count[14].r.part0[14] );
tran (\sa_count[14][14] , \sa_count[14].f.lower[14] );
tran (\sa_count[14][13] , \sa_count[14].r.part0[13] );
tran (\sa_count[14][13] , \sa_count[14].f.lower[13] );
tran (\sa_count[14][12] , \sa_count[14].r.part0[12] );
tran (\sa_count[14][12] , \sa_count[14].f.lower[12] );
tran (\sa_count[14][11] , \sa_count[14].r.part0[11] );
tran (\sa_count[14][11] , \sa_count[14].f.lower[11] );
tran (\sa_count[14][10] , \sa_count[14].r.part0[10] );
tran (\sa_count[14][10] , \sa_count[14].f.lower[10] );
tran (\sa_count[14][9] , \sa_count[14].r.part0[9] );
tran (\sa_count[14][9] , \sa_count[14].f.lower[9] );
tran (\sa_count[14][8] , \sa_count[14].r.part0[8] );
tran (\sa_count[14][8] , \sa_count[14].f.lower[8] );
tran (\sa_count[14][7] , \sa_count[14].r.part0[7] );
tran (\sa_count[14][7] , \sa_count[14].f.lower[7] );
tran (\sa_count[14][6] , \sa_count[14].r.part0[6] );
tran (\sa_count[14][6] , \sa_count[14].f.lower[6] );
tran (\sa_count[14][5] , \sa_count[14].r.part0[5] );
tran (\sa_count[14][5] , \sa_count[14].f.lower[5] );
tran (\sa_count[14][4] , \sa_count[14].r.part0[4] );
tran (\sa_count[14][4] , \sa_count[14].f.lower[4] );
tran (\sa_count[14][3] , \sa_count[14].r.part0[3] );
tran (\sa_count[14][3] , \sa_count[14].f.lower[3] );
tran (\sa_count[14][2] , \sa_count[14].r.part0[2] );
tran (\sa_count[14][2] , \sa_count[14].f.lower[2] );
tran (\sa_count[14][1] , \sa_count[14].r.part0[1] );
tran (\sa_count[14][1] , \sa_count[14].f.lower[1] );
tran (\sa_count[14][0] , \sa_count[14].r.part0[0] );
tran (\sa_count[14][0] , \sa_count[14].f.lower[0] );
tran (\sa_count[13][63] , \sa_count[13].r.part1[31] );
tran (\sa_count[13][63] , \sa_count[13].f.unused[13] );
tran (\sa_count[13][62] , \sa_count[13].r.part1[30] );
tran (\sa_count[13][62] , \sa_count[13].f.unused[12] );
tran (\sa_count[13][61] , \sa_count[13].r.part1[29] );
tran (\sa_count[13][61] , \sa_count[13].f.unused[11] );
tran (\sa_count[13][60] , \sa_count[13].r.part1[28] );
tran (\sa_count[13][60] , \sa_count[13].f.unused[10] );
tran (\sa_count[13][59] , \sa_count[13].r.part1[27] );
tran (\sa_count[13][59] , \sa_count[13].f.unused[9] );
tran (\sa_count[13][58] , \sa_count[13].r.part1[26] );
tran (\sa_count[13][58] , \sa_count[13].f.unused[8] );
tran (\sa_count[13][57] , \sa_count[13].r.part1[25] );
tran (\sa_count[13][57] , \sa_count[13].f.unused[7] );
tran (\sa_count[13][56] , \sa_count[13].r.part1[24] );
tran (\sa_count[13][56] , \sa_count[13].f.unused[6] );
tran (\sa_count[13][55] , \sa_count[13].r.part1[23] );
tran (\sa_count[13][55] , \sa_count[13].f.unused[5] );
tran (\sa_count[13][54] , \sa_count[13].r.part1[22] );
tran (\sa_count[13][54] , \sa_count[13].f.unused[4] );
tran (\sa_count[13][53] , \sa_count[13].r.part1[21] );
tran (\sa_count[13][53] , \sa_count[13].f.unused[3] );
tran (\sa_count[13][52] , \sa_count[13].r.part1[20] );
tran (\sa_count[13][52] , \sa_count[13].f.unused[2] );
tran (\sa_count[13][51] , \sa_count[13].r.part1[19] );
tran (\sa_count[13][51] , \sa_count[13].f.unused[1] );
tran (\sa_count[13][50] , \sa_count[13].r.part1[18] );
tran (\sa_count[13][50] , \sa_count[13].f.unused[0] );
tran (\sa_count[13][49] , \sa_count[13].r.part1[17] );
tran (\sa_count[13][49] , \sa_count[13].f.upper[17] );
tran (\sa_count[13][48] , \sa_count[13].r.part1[16] );
tran (\sa_count[13][48] , \sa_count[13].f.upper[16] );
tran (\sa_count[13][47] , \sa_count[13].r.part1[15] );
tran (\sa_count[13][47] , \sa_count[13].f.upper[15] );
tran (\sa_count[13][46] , \sa_count[13].r.part1[14] );
tran (\sa_count[13][46] , \sa_count[13].f.upper[14] );
tran (\sa_count[13][45] , \sa_count[13].r.part1[13] );
tran (\sa_count[13][45] , \sa_count[13].f.upper[13] );
tran (\sa_count[13][44] , \sa_count[13].r.part1[12] );
tran (\sa_count[13][44] , \sa_count[13].f.upper[12] );
tran (\sa_count[13][43] , \sa_count[13].r.part1[11] );
tran (\sa_count[13][43] , \sa_count[13].f.upper[11] );
tran (\sa_count[13][42] , \sa_count[13].r.part1[10] );
tran (\sa_count[13][42] , \sa_count[13].f.upper[10] );
tran (\sa_count[13][41] , \sa_count[13].r.part1[9] );
tran (\sa_count[13][41] , \sa_count[13].f.upper[9] );
tran (\sa_count[13][40] , \sa_count[13].r.part1[8] );
tran (\sa_count[13][40] , \sa_count[13].f.upper[8] );
tran (\sa_count[13][39] , \sa_count[13].r.part1[7] );
tran (\sa_count[13][39] , \sa_count[13].f.upper[7] );
tran (\sa_count[13][38] , \sa_count[13].r.part1[6] );
tran (\sa_count[13][38] , \sa_count[13].f.upper[6] );
tran (\sa_count[13][37] , \sa_count[13].r.part1[5] );
tran (\sa_count[13][37] , \sa_count[13].f.upper[5] );
tran (\sa_count[13][36] , \sa_count[13].r.part1[4] );
tran (\sa_count[13][36] , \sa_count[13].f.upper[4] );
tran (\sa_count[13][35] , \sa_count[13].r.part1[3] );
tran (\sa_count[13][35] , \sa_count[13].f.upper[3] );
tran (\sa_count[13][34] , \sa_count[13].r.part1[2] );
tran (\sa_count[13][34] , \sa_count[13].f.upper[2] );
tran (\sa_count[13][33] , \sa_count[13].r.part1[1] );
tran (\sa_count[13][33] , \sa_count[13].f.upper[1] );
tran (\sa_count[13][32] , \sa_count[13].r.part1[0] );
tran (\sa_count[13][32] , \sa_count[13].f.upper[0] );
tran (\sa_count[13][31] , \sa_count[13].r.part0[31] );
tran (\sa_count[13][31] , \sa_count[13].f.lower[31] );
tran (\sa_count[13][30] , \sa_count[13].r.part0[30] );
tran (\sa_count[13][30] , \sa_count[13].f.lower[30] );
tran (\sa_count[13][29] , \sa_count[13].r.part0[29] );
tran (\sa_count[13][29] , \sa_count[13].f.lower[29] );
tran (\sa_count[13][28] , \sa_count[13].r.part0[28] );
tran (\sa_count[13][28] , \sa_count[13].f.lower[28] );
tran (\sa_count[13][27] , \sa_count[13].r.part0[27] );
tran (\sa_count[13][27] , \sa_count[13].f.lower[27] );
tran (\sa_count[13][26] , \sa_count[13].r.part0[26] );
tran (\sa_count[13][26] , \sa_count[13].f.lower[26] );
tran (\sa_count[13][25] , \sa_count[13].r.part0[25] );
tran (\sa_count[13][25] , \sa_count[13].f.lower[25] );
tran (\sa_count[13][24] , \sa_count[13].r.part0[24] );
tran (\sa_count[13][24] , \sa_count[13].f.lower[24] );
tran (\sa_count[13][23] , \sa_count[13].r.part0[23] );
tran (\sa_count[13][23] , \sa_count[13].f.lower[23] );
tran (\sa_count[13][22] , \sa_count[13].r.part0[22] );
tran (\sa_count[13][22] , \sa_count[13].f.lower[22] );
tran (\sa_count[13][21] , \sa_count[13].r.part0[21] );
tran (\sa_count[13][21] , \sa_count[13].f.lower[21] );
tran (\sa_count[13][20] , \sa_count[13].r.part0[20] );
tran (\sa_count[13][20] , \sa_count[13].f.lower[20] );
tran (\sa_count[13][19] , \sa_count[13].r.part0[19] );
tran (\sa_count[13][19] , \sa_count[13].f.lower[19] );
tran (\sa_count[13][18] , \sa_count[13].r.part0[18] );
tran (\sa_count[13][18] , \sa_count[13].f.lower[18] );
tran (\sa_count[13][17] , \sa_count[13].r.part0[17] );
tran (\sa_count[13][17] , \sa_count[13].f.lower[17] );
tran (\sa_count[13][16] , \sa_count[13].r.part0[16] );
tran (\sa_count[13][16] , \sa_count[13].f.lower[16] );
tran (\sa_count[13][15] , \sa_count[13].r.part0[15] );
tran (\sa_count[13][15] , \sa_count[13].f.lower[15] );
tran (\sa_count[13][14] , \sa_count[13].r.part0[14] );
tran (\sa_count[13][14] , \sa_count[13].f.lower[14] );
tran (\sa_count[13][13] , \sa_count[13].r.part0[13] );
tran (\sa_count[13][13] , \sa_count[13].f.lower[13] );
tran (\sa_count[13][12] , \sa_count[13].r.part0[12] );
tran (\sa_count[13][12] , \sa_count[13].f.lower[12] );
tran (\sa_count[13][11] , \sa_count[13].r.part0[11] );
tran (\sa_count[13][11] , \sa_count[13].f.lower[11] );
tran (\sa_count[13][10] , \sa_count[13].r.part0[10] );
tran (\sa_count[13][10] , \sa_count[13].f.lower[10] );
tran (\sa_count[13][9] , \sa_count[13].r.part0[9] );
tran (\sa_count[13][9] , \sa_count[13].f.lower[9] );
tran (\sa_count[13][8] , \sa_count[13].r.part0[8] );
tran (\sa_count[13][8] , \sa_count[13].f.lower[8] );
tran (\sa_count[13][7] , \sa_count[13].r.part0[7] );
tran (\sa_count[13][7] , \sa_count[13].f.lower[7] );
tran (\sa_count[13][6] , \sa_count[13].r.part0[6] );
tran (\sa_count[13][6] , \sa_count[13].f.lower[6] );
tran (\sa_count[13][5] , \sa_count[13].r.part0[5] );
tran (\sa_count[13][5] , \sa_count[13].f.lower[5] );
tran (\sa_count[13][4] , \sa_count[13].r.part0[4] );
tran (\sa_count[13][4] , \sa_count[13].f.lower[4] );
tran (\sa_count[13][3] , \sa_count[13].r.part0[3] );
tran (\sa_count[13][3] , \sa_count[13].f.lower[3] );
tran (\sa_count[13][2] , \sa_count[13].r.part0[2] );
tran (\sa_count[13][2] , \sa_count[13].f.lower[2] );
tran (\sa_count[13][1] , \sa_count[13].r.part0[1] );
tran (\sa_count[13][1] , \sa_count[13].f.lower[1] );
tran (\sa_count[13][0] , \sa_count[13].r.part0[0] );
tran (\sa_count[13][0] , \sa_count[13].f.lower[0] );
tran (\sa_count[12][63] , \sa_count[12].r.part1[31] );
tran (\sa_count[12][63] , \sa_count[12].f.unused[13] );
tran (\sa_count[12][62] , \sa_count[12].r.part1[30] );
tran (\sa_count[12][62] , \sa_count[12].f.unused[12] );
tran (\sa_count[12][61] , \sa_count[12].r.part1[29] );
tran (\sa_count[12][61] , \sa_count[12].f.unused[11] );
tran (\sa_count[12][60] , \sa_count[12].r.part1[28] );
tran (\sa_count[12][60] , \sa_count[12].f.unused[10] );
tran (\sa_count[12][59] , \sa_count[12].r.part1[27] );
tran (\sa_count[12][59] , \sa_count[12].f.unused[9] );
tran (\sa_count[12][58] , \sa_count[12].r.part1[26] );
tran (\sa_count[12][58] , \sa_count[12].f.unused[8] );
tran (\sa_count[12][57] , \sa_count[12].r.part1[25] );
tran (\sa_count[12][57] , \sa_count[12].f.unused[7] );
tran (\sa_count[12][56] , \sa_count[12].r.part1[24] );
tran (\sa_count[12][56] , \sa_count[12].f.unused[6] );
tran (\sa_count[12][55] , \sa_count[12].r.part1[23] );
tran (\sa_count[12][55] , \sa_count[12].f.unused[5] );
tran (\sa_count[12][54] , \sa_count[12].r.part1[22] );
tran (\sa_count[12][54] , \sa_count[12].f.unused[4] );
tran (\sa_count[12][53] , \sa_count[12].r.part1[21] );
tran (\sa_count[12][53] , \sa_count[12].f.unused[3] );
tran (\sa_count[12][52] , \sa_count[12].r.part1[20] );
tran (\sa_count[12][52] , \sa_count[12].f.unused[2] );
tran (\sa_count[12][51] , \sa_count[12].r.part1[19] );
tran (\sa_count[12][51] , \sa_count[12].f.unused[1] );
tran (\sa_count[12][50] , \sa_count[12].r.part1[18] );
tran (\sa_count[12][50] , \sa_count[12].f.unused[0] );
tran (\sa_count[12][49] , \sa_count[12].r.part1[17] );
tran (\sa_count[12][49] , \sa_count[12].f.upper[17] );
tran (\sa_count[12][48] , \sa_count[12].r.part1[16] );
tran (\sa_count[12][48] , \sa_count[12].f.upper[16] );
tran (\sa_count[12][47] , \sa_count[12].r.part1[15] );
tran (\sa_count[12][47] , \sa_count[12].f.upper[15] );
tran (\sa_count[12][46] , \sa_count[12].r.part1[14] );
tran (\sa_count[12][46] , \sa_count[12].f.upper[14] );
tran (\sa_count[12][45] , \sa_count[12].r.part1[13] );
tran (\sa_count[12][45] , \sa_count[12].f.upper[13] );
tran (\sa_count[12][44] , \sa_count[12].r.part1[12] );
tran (\sa_count[12][44] , \sa_count[12].f.upper[12] );
tran (\sa_count[12][43] , \sa_count[12].r.part1[11] );
tran (\sa_count[12][43] , \sa_count[12].f.upper[11] );
tran (\sa_count[12][42] , \sa_count[12].r.part1[10] );
tran (\sa_count[12][42] , \sa_count[12].f.upper[10] );
tran (\sa_count[12][41] , \sa_count[12].r.part1[9] );
tran (\sa_count[12][41] , \sa_count[12].f.upper[9] );
tran (\sa_count[12][40] , \sa_count[12].r.part1[8] );
tran (\sa_count[12][40] , \sa_count[12].f.upper[8] );
tran (\sa_count[12][39] , \sa_count[12].r.part1[7] );
tran (\sa_count[12][39] , \sa_count[12].f.upper[7] );
tran (\sa_count[12][38] , \sa_count[12].r.part1[6] );
tran (\sa_count[12][38] , \sa_count[12].f.upper[6] );
tran (\sa_count[12][37] , \sa_count[12].r.part1[5] );
tran (\sa_count[12][37] , \sa_count[12].f.upper[5] );
tran (\sa_count[12][36] , \sa_count[12].r.part1[4] );
tran (\sa_count[12][36] , \sa_count[12].f.upper[4] );
tran (\sa_count[12][35] , \sa_count[12].r.part1[3] );
tran (\sa_count[12][35] , \sa_count[12].f.upper[3] );
tran (\sa_count[12][34] , \sa_count[12].r.part1[2] );
tran (\sa_count[12][34] , \sa_count[12].f.upper[2] );
tran (\sa_count[12][33] , \sa_count[12].r.part1[1] );
tran (\sa_count[12][33] , \sa_count[12].f.upper[1] );
tran (\sa_count[12][32] , \sa_count[12].r.part1[0] );
tran (\sa_count[12][32] , \sa_count[12].f.upper[0] );
tran (\sa_count[12][31] , \sa_count[12].r.part0[31] );
tran (\sa_count[12][31] , \sa_count[12].f.lower[31] );
tran (\sa_count[12][30] , \sa_count[12].r.part0[30] );
tran (\sa_count[12][30] , \sa_count[12].f.lower[30] );
tran (\sa_count[12][29] , \sa_count[12].r.part0[29] );
tran (\sa_count[12][29] , \sa_count[12].f.lower[29] );
tran (\sa_count[12][28] , \sa_count[12].r.part0[28] );
tran (\sa_count[12][28] , \sa_count[12].f.lower[28] );
tran (\sa_count[12][27] , \sa_count[12].r.part0[27] );
tran (\sa_count[12][27] , \sa_count[12].f.lower[27] );
tran (\sa_count[12][26] , \sa_count[12].r.part0[26] );
tran (\sa_count[12][26] , \sa_count[12].f.lower[26] );
tran (\sa_count[12][25] , \sa_count[12].r.part0[25] );
tran (\sa_count[12][25] , \sa_count[12].f.lower[25] );
tran (\sa_count[12][24] , \sa_count[12].r.part0[24] );
tran (\sa_count[12][24] , \sa_count[12].f.lower[24] );
tran (\sa_count[12][23] , \sa_count[12].r.part0[23] );
tran (\sa_count[12][23] , \sa_count[12].f.lower[23] );
tran (\sa_count[12][22] , \sa_count[12].r.part0[22] );
tran (\sa_count[12][22] , \sa_count[12].f.lower[22] );
tran (\sa_count[12][21] , \sa_count[12].r.part0[21] );
tran (\sa_count[12][21] , \sa_count[12].f.lower[21] );
tran (\sa_count[12][20] , \sa_count[12].r.part0[20] );
tran (\sa_count[12][20] , \sa_count[12].f.lower[20] );
tran (\sa_count[12][19] , \sa_count[12].r.part0[19] );
tran (\sa_count[12][19] , \sa_count[12].f.lower[19] );
tran (\sa_count[12][18] , \sa_count[12].r.part0[18] );
tran (\sa_count[12][18] , \sa_count[12].f.lower[18] );
tran (\sa_count[12][17] , \sa_count[12].r.part0[17] );
tran (\sa_count[12][17] , \sa_count[12].f.lower[17] );
tran (\sa_count[12][16] , \sa_count[12].r.part0[16] );
tran (\sa_count[12][16] , \sa_count[12].f.lower[16] );
tran (\sa_count[12][15] , \sa_count[12].r.part0[15] );
tran (\sa_count[12][15] , \sa_count[12].f.lower[15] );
tran (\sa_count[12][14] , \sa_count[12].r.part0[14] );
tran (\sa_count[12][14] , \sa_count[12].f.lower[14] );
tran (\sa_count[12][13] , \sa_count[12].r.part0[13] );
tran (\sa_count[12][13] , \sa_count[12].f.lower[13] );
tran (\sa_count[12][12] , \sa_count[12].r.part0[12] );
tran (\sa_count[12][12] , \sa_count[12].f.lower[12] );
tran (\sa_count[12][11] , \sa_count[12].r.part0[11] );
tran (\sa_count[12][11] , \sa_count[12].f.lower[11] );
tran (\sa_count[12][10] , \sa_count[12].r.part0[10] );
tran (\sa_count[12][10] , \sa_count[12].f.lower[10] );
tran (\sa_count[12][9] , \sa_count[12].r.part0[9] );
tran (\sa_count[12][9] , \sa_count[12].f.lower[9] );
tran (\sa_count[12][8] , \sa_count[12].r.part0[8] );
tran (\sa_count[12][8] , \sa_count[12].f.lower[8] );
tran (\sa_count[12][7] , \sa_count[12].r.part0[7] );
tran (\sa_count[12][7] , \sa_count[12].f.lower[7] );
tran (\sa_count[12][6] , \sa_count[12].r.part0[6] );
tran (\sa_count[12][6] , \sa_count[12].f.lower[6] );
tran (\sa_count[12][5] , \sa_count[12].r.part0[5] );
tran (\sa_count[12][5] , \sa_count[12].f.lower[5] );
tran (\sa_count[12][4] , \sa_count[12].r.part0[4] );
tran (\sa_count[12][4] , \sa_count[12].f.lower[4] );
tran (\sa_count[12][3] , \sa_count[12].r.part0[3] );
tran (\sa_count[12][3] , \sa_count[12].f.lower[3] );
tran (\sa_count[12][2] , \sa_count[12].r.part0[2] );
tran (\sa_count[12][2] , \sa_count[12].f.lower[2] );
tran (\sa_count[12][1] , \sa_count[12].r.part0[1] );
tran (\sa_count[12][1] , \sa_count[12].f.lower[1] );
tran (\sa_count[12][0] , \sa_count[12].r.part0[0] );
tran (\sa_count[12][0] , \sa_count[12].f.lower[0] );
tran (\sa_count[11][63] , \sa_count[11].r.part1[31] );
tran (\sa_count[11][63] , \sa_count[11].f.unused[13] );
tran (\sa_count[11][62] , \sa_count[11].r.part1[30] );
tran (\sa_count[11][62] , \sa_count[11].f.unused[12] );
tran (\sa_count[11][61] , \sa_count[11].r.part1[29] );
tran (\sa_count[11][61] , \sa_count[11].f.unused[11] );
tran (\sa_count[11][60] , \sa_count[11].r.part1[28] );
tran (\sa_count[11][60] , \sa_count[11].f.unused[10] );
tran (\sa_count[11][59] , \sa_count[11].r.part1[27] );
tran (\sa_count[11][59] , \sa_count[11].f.unused[9] );
tran (\sa_count[11][58] , \sa_count[11].r.part1[26] );
tran (\sa_count[11][58] , \sa_count[11].f.unused[8] );
tran (\sa_count[11][57] , \sa_count[11].r.part1[25] );
tran (\sa_count[11][57] , \sa_count[11].f.unused[7] );
tran (\sa_count[11][56] , \sa_count[11].r.part1[24] );
tran (\sa_count[11][56] , \sa_count[11].f.unused[6] );
tran (\sa_count[11][55] , \sa_count[11].r.part1[23] );
tran (\sa_count[11][55] , \sa_count[11].f.unused[5] );
tran (\sa_count[11][54] , \sa_count[11].r.part1[22] );
tran (\sa_count[11][54] , \sa_count[11].f.unused[4] );
tran (\sa_count[11][53] , \sa_count[11].r.part1[21] );
tran (\sa_count[11][53] , \sa_count[11].f.unused[3] );
tran (\sa_count[11][52] , \sa_count[11].r.part1[20] );
tran (\sa_count[11][52] , \sa_count[11].f.unused[2] );
tran (\sa_count[11][51] , \sa_count[11].r.part1[19] );
tran (\sa_count[11][51] , \sa_count[11].f.unused[1] );
tran (\sa_count[11][50] , \sa_count[11].r.part1[18] );
tran (\sa_count[11][50] , \sa_count[11].f.unused[0] );
tran (\sa_count[11][49] , \sa_count[11].r.part1[17] );
tran (\sa_count[11][49] , \sa_count[11].f.upper[17] );
tran (\sa_count[11][48] , \sa_count[11].r.part1[16] );
tran (\sa_count[11][48] , \sa_count[11].f.upper[16] );
tran (\sa_count[11][47] , \sa_count[11].r.part1[15] );
tran (\sa_count[11][47] , \sa_count[11].f.upper[15] );
tran (\sa_count[11][46] , \sa_count[11].r.part1[14] );
tran (\sa_count[11][46] , \sa_count[11].f.upper[14] );
tran (\sa_count[11][45] , \sa_count[11].r.part1[13] );
tran (\sa_count[11][45] , \sa_count[11].f.upper[13] );
tran (\sa_count[11][44] , \sa_count[11].r.part1[12] );
tran (\sa_count[11][44] , \sa_count[11].f.upper[12] );
tran (\sa_count[11][43] , \sa_count[11].r.part1[11] );
tran (\sa_count[11][43] , \sa_count[11].f.upper[11] );
tran (\sa_count[11][42] , \sa_count[11].r.part1[10] );
tran (\sa_count[11][42] , \sa_count[11].f.upper[10] );
tran (\sa_count[11][41] , \sa_count[11].r.part1[9] );
tran (\sa_count[11][41] , \sa_count[11].f.upper[9] );
tran (\sa_count[11][40] , \sa_count[11].r.part1[8] );
tran (\sa_count[11][40] , \sa_count[11].f.upper[8] );
tran (\sa_count[11][39] , \sa_count[11].r.part1[7] );
tran (\sa_count[11][39] , \sa_count[11].f.upper[7] );
tran (\sa_count[11][38] , \sa_count[11].r.part1[6] );
tran (\sa_count[11][38] , \sa_count[11].f.upper[6] );
tran (\sa_count[11][37] , \sa_count[11].r.part1[5] );
tran (\sa_count[11][37] , \sa_count[11].f.upper[5] );
tran (\sa_count[11][36] , \sa_count[11].r.part1[4] );
tran (\sa_count[11][36] , \sa_count[11].f.upper[4] );
tran (\sa_count[11][35] , \sa_count[11].r.part1[3] );
tran (\sa_count[11][35] , \sa_count[11].f.upper[3] );
tran (\sa_count[11][34] , \sa_count[11].r.part1[2] );
tran (\sa_count[11][34] , \sa_count[11].f.upper[2] );
tran (\sa_count[11][33] , \sa_count[11].r.part1[1] );
tran (\sa_count[11][33] , \sa_count[11].f.upper[1] );
tran (\sa_count[11][32] , \sa_count[11].r.part1[0] );
tran (\sa_count[11][32] , \sa_count[11].f.upper[0] );
tran (\sa_count[11][31] , \sa_count[11].r.part0[31] );
tran (\sa_count[11][31] , \sa_count[11].f.lower[31] );
tran (\sa_count[11][30] , \sa_count[11].r.part0[30] );
tran (\sa_count[11][30] , \sa_count[11].f.lower[30] );
tran (\sa_count[11][29] , \sa_count[11].r.part0[29] );
tran (\sa_count[11][29] , \sa_count[11].f.lower[29] );
tran (\sa_count[11][28] , \sa_count[11].r.part0[28] );
tran (\sa_count[11][28] , \sa_count[11].f.lower[28] );
tran (\sa_count[11][27] , \sa_count[11].r.part0[27] );
tran (\sa_count[11][27] , \sa_count[11].f.lower[27] );
tran (\sa_count[11][26] , \sa_count[11].r.part0[26] );
tran (\sa_count[11][26] , \sa_count[11].f.lower[26] );
tran (\sa_count[11][25] , \sa_count[11].r.part0[25] );
tran (\sa_count[11][25] , \sa_count[11].f.lower[25] );
tran (\sa_count[11][24] , \sa_count[11].r.part0[24] );
tran (\sa_count[11][24] , \sa_count[11].f.lower[24] );
tran (\sa_count[11][23] , \sa_count[11].r.part0[23] );
tran (\sa_count[11][23] , \sa_count[11].f.lower[23] );
tran (\sa_count[11][22] , \sa_count[11].r.part0[22] );
tran (\sa_count[11][22] , \sa_count[11].f.lower[22] );
tran (\sa_count[11][21] , \sa_count[11].r.part0[21] );
tran (\sa_count[11][21] , \sa_count[11].f.lower[21] );
tran (\sa_count[11][20] , \sa_count[11].r.part0[20] );
tran (\sa_count[11][20] , \sa_count[11].f.lower[20] );
tran (\sa_count[11][19] , \sa_count[11].r.part0[19] );
tran (\sa_count[11][19] , \sa_count[11].f.lower[19] );
tran (\sa_count[11][18] , \sa_count[11].r.part0[18] );
tran (\sa_count[11][18] , \sa_count[11].f.lower[18] );
tran (\sa_count[11][17] , \sa_count[11].r.part0[17] );
tran (\sa_count[11][17] , \sa_count[11].f.lower[17] );
tran (\sa_count[11][16] , \sa_count[11].r.part0[16] );
tran (\sa_count[11][16] , \sa_count[11].f.lower[16] );
tran (\sa_count[11][15] , \sa_count[11].r.part0[15] );
tran (\sa_count[11][15] , \sa_count[11].f.lower[15] );
tran (\sa_count[11][14] , \sa_count[11].r.part0[14] );
tran (\sa_count[11][14] , \sa_count[11].f.lower[14] );
tran (\sa_count[11][13] , \sa_count[11].r.part0[13] );
tran (\sa_count[11][13] , \sa_count[11].f.lower[13] );
tran (\sa_count[11][12] , \sa_count[11].r.part0[12] );
tran (\sa_count[11][12] , \sa_count[11].f.lower[12] );
tran (\sa_count[11][11] , \sa_count[11].r.part0[11] );
tran (\sa_count[11][11] , \sa_count[11].f.lower[11] );
tran (\sa_count[11][10] , \sa_count[11].r.part0[10] );
tran (\sa_count[11][10] , \sa_count[11].f.lower[10] );
tran (\sa_count[11][9] , \sa_count[11].r.part0[9] );
tran (\sa_count[11][9] , \sa_count[11].f.lower[9] );
tran (\sa_count[11][8] , \sa_count[11].r.part0[8] );
tran (\sa_count[11][8] , \sa_count[11].f.lower[8] );
tran (\sa_count[11][7] , \sa_count[11].r.part0[7] );
tran (\sa_count[11][7] , \sa_count[11].f.lower[7] );
tran (\sa_count[11][6] , \sa_count[11].r.part0[6] );
tran (\sa_count[11][6] , \sa_count[11].f.lower[6] );
tran (\sa_count[11][5] , \sa_count[11].r.part0[5] );
tran (\sa_count[11][5] , \sa_count[11].f.lower[5] );
tran (\sa_count[11][4] , \sa_count[11].r.part0[4] );
tran (\sa_count[11][4] , \sa_count[11].f.lower[4] );
tran (\sa_count[11][3] , \sa_count[11].r.part0[3] );
tran (\sa_count[11][3] , \sa_count[11].f.lower[3] );
tran (\sa_count[11][2] , \sa_count[11].r.part0[2] );
tran (\sa_count[11][2] , \sa_count[11].f.lower[2] );
tran (\sa_count[11][1] , \sa_count[11].r.part0[1] );
tran (\sa_count[11][1] , \sa_count[11].f.lower[1] );
tran (\sa_count[11][0] , \sa_count[11].r.part0[0] );
tran (\sa_count[11][0] , \sa_count[11].f.lower[0] );
tran (\sa_count[10][63] , \sa_count[10].r.part1[31] );
tran (\sa_count[10][63] , \sa_count[10].f.unused[13] );
tran (\sa_count[10][62] , \sa_count[10].r.part1[30] );
tran (\sa_count[10][62] , \sa_count[10].f.unused[12] );
tran (\sa_count[10][61] , \sa_count[10].r.part1[29] );
tran (\sa_count[10][61] , \sa_count[10].f.unused[11] );
tran (\sa_count[10][60] , \sa_count[10].r.part1[28] );
tran (\sa_count[10][60] , \sa_count[10].f.unused[10] );
tran (\sa_count[10][59] , \sa_count[10].r.part1[27] );
tran (\sa_count[10][59] , \sa_count[10].f.unused[9] );
tran (\sa_count[10][58] , \sa_count[10].r.part1[26] );
tran (\sa_count[10][58] , \sa_count[10].f.unused[8] );
tran (\sa_count[10][57] , \sa_count[10].r.part1[25] );
tran (\sa_count[10][57] , \sa_count[10].f.unused[7] );
tran (\sa_count[10][56] , \sa_count[10].r.part1[24] );
tran (\sa_count[10][56] , \sa_count[10].f.unused[6] );
tran (\sa_count[10][55] , \sa_count[10].r.part1[23] );
tran (\sa_count[10][55] , \sa_count[10].f.unused[5] );
tran (\sa_count[10][54] , \sa_count[10].r.part1[22] );
tran (\sa_count[10][54] , \sa_count[10].f.unused[4] );
tran (\sa_count[10][53] , \sa_count[10].r.part1[21] );
tran (\sa_count[10][53] , \sa_count[10].f.unused[3] );
tran (\sa_count[10][52] , \sa_count[10].r.part1[20] );
tran (\sa_count[10][52] , \sa_count[10].f.unused[2] );
tran (\sa_count[10][51] , \sa_count[10].r.part1[19] );
tran (\sa_count[10][51] , \sa_count[10].f.unused[1] );
tran (\sa_count[10][50] , \sa_count[10].r.part1[18] );
tran (\sa_count[10][50] , \sa_count[10].f.unused[0] );
tran (\sa_count[10][49] , \sa_count[10].r.part1[17] );
tran (\sa_count[10][49] , \sa_count[10].f.upper[17] );
tran (\sa_count[10][48] , \sa_count[10].r.part1[16] );
tran (\sa_count[10][48] , \sa_count[10].f.upper[16] );
tran (\sa_count[10][47] , \sa_count[10].r.part1[15] );
tran (\sa_count[10][47] , \sa_count[10].f.upper[15] );
tran (\sa_count[10][46] , \sa_count[10].r.part1[14] );
tran (\sa_count[10][46] , \sa_count[10].f.upper[14] );
tran (\sa_count[10][45] , \sa_count[10].r.part1[13] );
tran (\sa_count[10][45] , \sa_count[10].f.upper[13] );
tran (\sa_count[10][44] , \sa_count[10].r.part1[12] );
tran (\sa_count[10][44] , \sa_count[10].f.upper[12] );
tran (\sa_count[10][43] , \sa_count[10].r.part1[11] );
tran (\sa_count[10][43] , \sa_count[10].f.upper[11] );
tran (\sa_count[10][42] , \sa_count[10].r.part1[10] );
tran (\sa_count[10][42] , \sa_count[10].f.upper[10] );
tran (\sa_count[10][41] , \sa_count[10].r.part1[9] );
tran (\sa_count[10][41] , \sa_count[10].f.upper[9] );
tran (\sa_count[10][40] , \sa_count[10].r.part1[8] );
tran (\sa_count[10][40] , \sa_count[10].f.upper[8] );
tran (\sa_count[10][39] , \sa_count[10].r.part1[7] );
tran (\sa_count[10][39] , \sa_count[10].f.upper[7] );
tran (\sa_count[10][38] , \sa_count[10].r.part1[6] );
tran (\sa_count[10][38] , \sa_count[10].f.upper[6] );
tran (\sa_count[10][37] , \sa_count[10].r.part1[5] );
tran (\sa_count[10][37] , \sa_count[10].f.upper[5] );
tran (\sa_count[10][36] , \sa_count[10].r.part1[4] );
tran (\sa_count[10][36] , \sa_count[10].f.upper[4] );
tran (\sa_count[10][35] , \sa_count[10].r.part1[3] );
tran (\sa_count[10][35] , \sa_count[10].f.upper[3] );
tran (\sa_count[10][34] , \sa_count[10].r.part1[2] );
tran (\sa_count[10][34] , \sa_count[10].f.upper[2] );
tran (\sa_count[10][33] , \sa_count[10].r.part1[1] );
tran (\sa_count[10][33] , \sa_count[10].f.upper[1] );
tran (\sa_count[10][32] , \sa_count[10].r.part1[0] );
tran (\sa_count[10][32] , \sa_count[10].f.upper[0] );
tran (\sa_count[10][31] , \sa_count[10].r.part0[31] );
tran (\sa_count[10][31] , \sa_count[10].f.lower[31] );
tran (\sa_count[10][30] , \sa_count[10].r.part0[30] );
tran (\sa_count[10][30] , \sa_count[10].f.lower[30] );
tran (\sa_count[10][29] , \sa_count[10].r.part0[29] );
tran (\sa_count[10][29] , \sa_count[10].f.lower[29] );
tran (\sa_count[10][28] , \sa_count[10].r.part0[28] );
tran (\sa_count[10][28] , \sa_count[10].f.lower[28] );
tran (\sa_count[10][27] , \sa_count[10].r.part0[27] );
tran (\sa_count[10][27] , \sa_count[10].f.lower[27] );
tran (\sa_count[10][26] , \sa_count[10].r.part0[26] );
tran (\sa_count[10][26] , \sa_count[10].f.lower[26] );
tran (\sa_count[10][25] , \sa_count[10].r.part0[25] );
tran (\sa_count[10][25] , \sa_count[10].f.lower[25] );
tran (\sa_count[10][24] , \sa_count[10].r.part0[24] );
tran (\sa_count[10][24] , \sa_count[10].f.lower[24] );
tran (\sa_count[10][23] , \sa_count[10].r.part0[23] );
tran (\sa_count[10][23] , \sa_count[10].f.lower[23] );
tran (\sa_count[10][22] , \sa_count[10].r.part0[22] );
tran (\sa_count[10][22] , \sa_count[10].f.lower[22] );
tran (\sa_count[10][21] , \sa_count[10].r.part0[21] );
tran (\sa_count[10][21] , \sa_count[10].f.lower[21] );
tran (\sa_count[10][20] , \sa_count[10].r.part0[20] );
tran (\sa_count[10][20] , \sa_count[10].f.lower[20] );
tran (\sa_count[10][19] , \sa_count[10].r.part0[19] );
tran (\sa_count[10][19] , \sa_count[10].f.lower[19] );
tran (\sa_count[10][18] , \sa_count[10].r.part0[18] );
tran (\sa_count[10][18] , \sa_count[10].f.lower[18] );
tran (\sa_count[10][17] , \sa_count[10].r.part0[17] );
tran (\sa_count[10][17] , \sa_count[10].f.lower[17] );
tran (\sa_count[10][16] , \sa_count[10].r.part0[16] );
tran (\sa_count[10][16] , \sa_count[10].f.lower[16] );
tran (\sa_count[10][15] , \sa_count[10].r.part0[15] );
tran (\sa_count[10][15] , \sa_count[10].f.lower[15] );
tran (\sa_count[10][14] , \sa_count[10].r.part0[14] );
tran (\sa_count[10][14] , \sa_count[10].f.lower[14] );
tran (\sa_count[10][13] , \sa_count[10].r.part0[13] );
tran (\sa_count[10][13] , \sa_count[10].f.lower[13] );
tran (\sa_count[10][12] , \sa_count[10].r.part0[12] );
tran (\sa_count[10][12] , \sa_count[10].f.lower[12] );
tran (\sa_count[10][11] , \sa_count[10].r.part0[11] );
tran (\sa_count[10][11] , \sa_count[10].f.lower[11] );
tran (\sa_count[10][10] , \sa_count[10].r.part0[10] );
tran (\sa_count[10][10] , \sa_count[10].f.lower[10] );
tran (\sa_count[10][9] , \sa_count[10].r.part0[9] );
tran (\sa_count[10][9] , \sa_count[10].f.lower[9] );
tran (\sa_count[10][8] , \sa_count[10].r.part0[8] );
tran (\sa_count[10][8] , \sa_count[10].f.lower[8] );
tran (\sa_count[10][7] , \sa_count[10].r.part0[7] );
tran (\sa_count[10][7] , \sa_count[10].f.lower[7] );
tran (\sa_count[10][6] , \sa_count[10].r.part0[6] );
tran (\sa_count[10][6] , \sa_count[10].f.lower[6] );
tran (\sa_count[10][5] , \sa_count[10].r.part0[5] );
tran (\sa_count[10][5] , \sa_count[10].f.lower[5] );
tran (\sa_count[10][4] , \sa_count[10].r.part0[4] );
tran (\sa_count[10][4] , \sa_count[10].f.lower[4] );
tran (\sa_count[10][3] , \sa_count[10].r.part0[3] );
tran (\sa_count[10][3] , \sa_count[10].f.lower[3] );
tran (\sa_count[10][2] , \sa_count[10].r.part0[2] );
tran (\sa_count[10][2] , \sa_count[10].f.lower[2] );
tran (\sa_count[10][1] , \sa_count[10].r.part0[1] );
tran (\sa_count[10][1] , \sa_count[10].f.lower[1] );
tran (\sa_count[10][0] , \sa_count[10].r.part0[0] );
tran (\sa_count[10][0] , \sa_count[10].f.lower[0] );
tran (\sa_count[9][63] , \sa_count[9].r.part1[31] );
tran (\sa_count[9][63] , \sa_count[9].f.unused[13] );
tran (\sa_count[9][62] , \sa_count[9].r.part1[30] );
tran (\sa_count[9][62] , \sa_count[9].f.unused[12] );
tran (\sa_count[9][61] , \sa_count[9].r.part1[29] );
tran (\sa_count[9][61] , \sa_count[9].f.unused[11] );
tran (\sa_count[9][60] , \sa_count[9].r.part1[28] );
tran (\sa_count[9][60] , \sa_count[9].f.unused[10] );
tran (\sa_count[9][59] , \sa_count[9].r.part1[27] );
tran (\sa_count[9][59] , \sa_count[9].f.unused[9] );
tran (\sa_count[9][58] , \sa_count[9].r.part1[26] );
tran (\sa_count[9][58] , \sa_count[9].f.unused[8] );
tran (\sa_count[9][57] , \sa_count[9].r.part1[25] );
tran (\sa_count[9][57] , \sa_count[9].f.unused[7] );
tran (\sa_count[9][56] , \sa_count[9].r.part1[24] );
tran (\sa_count[9][56] , \sa_count[9].f.unused[6] );
tran (\sa_count[9][55] , \sa_count[9].r.part1[23] );
tran (\sa_count[9][55] , \sa_count[9].f.unused[5] );
tran (\sa_count[9][54] , \sa_count[9].r.part1[22] );
tran (\sa_count[9][54] , \sa_count[9].f.unused[4] );
tran (\sa_count[9][53] , \sa_count[9].r.part1[21] );
tran (\sa_count[9][53] , \sa_count[9].f.unused[3] );
tran (\sa_count[9][52] , \sa_count[9].r.part1[20] );
tran (\sa_count[9][52] , \sa_count[9].f.unused[2] );
tran (\sa_count[9][51] , \sa_count[9].r.part1[19] );
tran (\sa_count[9][51] , \sa_count[9].f.unused[1] );
tran (\sa_count[9][50] , \sa_count[9].r.part1[18] );
tran (\sa_count[9][50] , \sa_count[9].f.unused[0] );
tran (\sa_count[9][49] , \sa_count[9].r.part1[17] );
tran (\sa_count[9][49] , \sa_count[9].f.upper[17] );
tran (\sa_count[9][48] , \sa_count[9].r.part1[16] );
tran (\sa_count[9][48] , \sa_count[9].f.upper[16] );
tran (\sa_count[9][47] , \sa_count[9].r.part1[15] );
tran (\sa_count[9][47] , \sa_count[9].f.upper[15] );
tran (\sa_count[9][46] , \sa_count[9].r.part1[14] );
tran (\sa_count[9][46] , \sa_count[9].f.upper[14] );
tran (\sa_count[9][45] , \sa_count[9].r.part1[13] );
tran (\sa_count[9][45] , \sa_count[9].f.upper[13] );
tran (\sa_count[9][44] , \sa_count[9].r.part1[12] );
tran (\sa_count[9][44] , \sa_count[9].f.upper[12] );
tran (\sa_count[9][43] , \sa_count[9].r.part1[11] );
tran (\sa_count[9][43] , \sa_count[9].f.upper[11] );
tran (\sa_count[9][42] , \sa_count[9].r.part1[10] );
tran (\sa_count[9][42] , \sa_count[9].f.upper[10] );
tran (\sa_count[9][41] , \sa_count[9].r.part1[9] );
tran (\sa_count[9][41] , \sa_count[9].f.upper[9] );
tran (\sa_count[9][40] , \sa_count[9].r.part1[8] );
tran (\sa_count[9][40] , \sa_count[9].f.upper[8] );
tran (\sa_count[9][39] , \sa_count[9].r.part1[7] );
tran (\sa_count[9][39] , \sa_count[9].f.upper[7] );
tran (\sa_count[9][38] , \sa_count[9].r.part1[6] );
tran (\sa_count[9][38] , \sa_count[9].f.upper[6] );
tran (\sa_count[9][37] , \sa_count[9].r.part1[5] );
tran (\sa_count[9][37] , \sa_count[9].f.upper[5] );
tran (\sa_count[9][36] , \sa_count[9].r.part1[4] );
tran (\sa_count[9][36] , \sa_count[9].f.upper[4] );
tran (\sa_count[9][35] , \sa_count[9].r.part1[3] );
tran (\sa_count[9][35] , \sa_count[9].f.upper[3] );
tran (\sa_count[9][34] , \sa_count[9].r.part1[2] );
tran (\sa_count[9][34] , \sa_count[9].f.upper[2] );
tran (\sa_count[9][33] , \sa_count[9].r.part1[1] );
tran (\sa_count[9][33] , \sa_count[9].f.upper[1] );
tran (\sa_count[9][32] , \sa_count[9].r.part1[0] );
tran (\sa_count[9][32] , \sa_count[9].f.upper[0] );
tran (\sa_count[9][31] , \sa_count[9].r.part0[31] );
tran (\sa_count[9][31] , \sa_count[9].f.lower[31] );
tran (\sa_count[9][30] , \sa_count[9].r.part0[30] );
tran (\sa_count[9][30] , \sa_count[9].f.lower[30] );
tran (\sa_count[9][29] , \sa_count[9].r.part0[29] );
tran (\sa_count[9][29] , \sa_count[9].f.lower[29] );
tran (\sa_count[9][28] , \sa_count[9].r.part0[28] );
tran (\sa_count[9][28] , \sa_count[9].f.lower[28] );
tran (\sa_count[9][27] , \sa_count[9].r.part0[27] );
tran (\sa_count[9][27] , \sa_count[9].f.lower[27] );
tran (\sa_count[9][26] , \sa_count[9].r.part0[26] );
tran (\sa_count[9][26] , \sa_count[9].f.lower[26] );
tran (\sa_count[9][25] , \sa_count[9].r.part0[25] );
tran (\sa_count[9][25] , \sa_count[9].f.lower[25] );
tran (\sa_count[9][24] , \sa_count[9].r.part0[24] );
tran (\sa_count[9][24] , \sa_count[9].f.lower[24] );
tran (\sa_count[9][23] , \sa_count[9].r.part0[23] );
tran (\sa_count[9][23] , \sa_count[9].f.lower[23] );
tran (\sa_count[9][22] , \sa_count[9].r.part0[22] );
tran (\sa_count[9][22] , \sa_count[9].f.lower[22] );
tran (\sa_count[9][21] , \sa_count[9].r.part0[21] );
tran (\sa_count[9][21] , \sa_count[9].f.lower[21] );
tran (\sa_count[9][20] , \sa_count[9].r.part0[20] );
tran (\sa_count[9][20] , \sa_count[9].f.lower[20] );
tran (\sa_count[9][19] , \sa_count[9].r.part0[19] );
tran (\sa_count[9][19] , \sa_count[9].f.lower[19] );
tran (\sa_count[9][18] , \sa_count[9].r.part0[18] );
tran (\sa_count[9][18] , \sa_count[9].f.lower[18] );
tran (\sa_count[9][17] , \sa_count[9].r.part0[17] );
tran (\sa_count[9][17] , \sa_count[9].f.lower[17] );
tran (\sa_count[9][16] , \sa_count[9].r.part0[16] );
tran (\sa_count[9][16] , \sa_count[9].f.lower[16] );
tran (\sa_count[9][15] , \sa_count[9].r.part0[15] );
tran (\sa_count[9][15] , \sa_count[9].f.lower[15] );
tran (\sa_count[9][14] , \sa_count[9].r.part0[14] );
tran (\sa_count[9][14] , \sa_count[9].f.lower[14] );
tran (\sa_count[9][13] , \sa_count[9].r.part0[13] );
tran (\sa_count[9][13] , \sa_count[9].f.lower[13] );
tran (\sa_count[9][12] , \sa_count[9].r.part0[12] );
tran (\sa_count[9][12] , \sa_count[9].f.lower[12] );
tran (\sa_count[9][11] , \sa_count[9].r.part0[11] );
tran (\sa_count[9][11] , \sa_count[9].f.lower[11] );
tran (\sa_count[9][10] , \sa_count[9].r.part0[10] );
tran (\sa_count[9][10] , \sa_count[9].f.lower[10] );
tran (\sa_count[9][9] , \sa_count[9].r.part0[9] );
tran (\sa_count[9][9] , \sa_count[9].f.lower[9] );
tran (\sa_count[9][8] , \sa_count[9].r.part0[8] );
tran (\sa_count[9][8] , \sa_count[9].f.lower[8] );
tran (\sa_count[9][7] , \sa_count[9].r.part0[7] );
tran (\sa_count[9][7] , \sa_count[9].f.lower[7] );
tran (\sa_count[9][6] , \sa_count[9].r.part0[6] );
tran (\sa_count[9][6] , \sa_count[9].f.lower[6] );
tran (\sa_count[9][5] , \sa_count[9].r.part0[5] );
tran (\sa_count[9][5] , \sa_count[9].f.lower[5] );
tran (\sa_count[9][4] , \sa_count[9].r.part0[4] );
tran (\sa_count[9][4] , \sa_count[9].f.lower[4] );
tran (\sa_count[9][3] , \sa_count[9].r.part0[3] );
tran (\sa_count[9][3] , \sa_count[9].f.lower[3] );
tran (\sa_count[9][2] , \sa_count[9].r.part0[2] );
tran (\sa_count[9][2] , \sa_count[9].f.lower[2] );
tran (\sa_count[9][1] , \sa_count[9].r.part0[1] );
tran (\sa_count[9][1] , \sa_count[9].f.lower[1] );
tran (\sa_count[9][0] , \sa_count[9].r.part0[0] );
tran (\sa_count[9][0] , \sa_count[9].f.lower[0] );
tran (\sa_count[8][63] , \sa_count[8].r.part1[31] );
tran (\sa_count[8][63] , \sa_count[8].f.unused[13] );
tran (\sa_count[8][62] , \sa_count[8].r.part1[30] );
tran (\sa_count[8][62] , \sa_count[8].f.unused[12] );
tran (\sa_count[8][61] , \sa_count[8].r.part1[29] );
tran (\sa_count[8][61] , \sa_count[8].f.unused[11] );
tran (\sa_count[8][60] , \sa_count[8].r.part1[28] );
tran (\sa_count[8][60] , \sa_count[8].f.unused[10] );
tran (\sa_count[8][59] , \sa_count[8].r.part1[27] );
tran (\sa_count[8][59] , \sa_count[8].f.unused[9] );
tran (\sa_count[8][58] , \sa_count[8].r.part1[26] );
tran (\sa_count[8][58] , \sa_count[8].f.unused[8] );
tran (\sa_count[8][57] , \sa_count[8].r.part1[25] );
tran (\sa_count[8][57] , \sa_count[8].f.unused[7] );
tran (\sa_count[8][56] , \sa_count[8].r.part1[24] );
tran (\sa_count[8][56] , \sa_count[8].f.unused[6] );
tran (\sa_count[8][55] , \sa_count[8].r.part1[23] );
tran (\sa_count[8][55] , \sa_count[8].f.unused[5] );
tran (\sa_count[8][54] , \sa_count[8].r.part1[22] );
tran (\sa_count[8][54] , \sa_count[8].f.unused[4] );
tran (\sa_count[8][53] , \sa_count[8].r.part1[21] );
tran (\sa_count[8][53] , \sa_count[8].f.unused[3] );
tran (\sa_count[8][52] , \sa_count[8].r.part1[20] );
tran (\sa_count[8][52] , \sa_count[8].f.unused[2] );
tran (\sa_count[8][51] , \sa_count[8].r.part1[19] );
tran (\sa_count[8][51] , \sa_count[8].f.unused[1] );
tran (\sa_count[8][50] , \sa_count[8].r.part1[18] );
tran (\sa_count[8][50] , \sa_count[8].f.unused[0] );
tran (\sa_count[8][49] , \sa_count[8].r.part1[17] );
tran (\sa_count[8][49] , \sa_count[8].f.upper[17] );
tran (\sa_count[8][48] , \sa_count[8].r.part1[16] );
tran (\sa_count[8][48] , \sa_count[8].f.upper[16] );
tran (\sa_count[8][47] , \sa_count[8].r.part1[15] );
tran (\sa_count[8][47] , \sa_count[8].f.upper[15] );
tran (\sa_count[8][46] , \sa_count[8].r.part1[14] );
tran (\sa_count[8][46] , \sa_count[8].f.upper[14] );
tran (\sa_count[8][45] , \sa_count[8].r.part1[13] );
tran (\sa_count[8][45] , \sa_count[8].f.upper[13] );
tran (\sa_count[8][44] , \sa_count[8].r.part1[12] );
tran (\sa_count[8][44] , \sa_count[8].f.upper[12] );
tran (\sa_count[8][43] , \sa_count[8].r.part1[11] );
tran (\sa_count[8][43] , \sa_count[8].f.upper[11] );
tran (\sa_count[8][42] , \sa_count[8].r.part1[10] );
tran (\sa_count[8][42] , \sa_count[8].f.upper[10] );
tran (\sa_count[8][41] , \sa_count[8].r.part1[9] );
tran (\sa_count[8][41] , \sa_count[8].f.upper[9] );
tran (\sa_count[8][40] , \sa_count[8].r.part1[8] );
tran (\sa_count[8][40] , \sa_count[8].f.upper[8] );
tran (\sa_count[8][39] , \sa_count[8].r.part1[7] );
tran (\sa_count[8][39] , \sa_count[8].f.upper[7] );
tran (\sa_count[8][38] , \sa_count[8].r.part1[6] );
tran (\sa_count[8][38] , \sa_count[8].f.upper[6] );
tran (\sa_count[8][37] , \sa_count[8].r.part1[5] );
tran (\sa_count[8][37] , \sa_count[8].f.upper[5] );
tran (\sa_count[8][36] , \sa_count[8].r.part1[4] );
tran (\sa_count[8][36] , \sa_count[8].f.upper[4] );
tran (\sa_count[8][35] , \sa_count[8].r.part1[3] );
tran (\sa_count[8][35] , \sa_count[8].f.upper[3] );
tran (\sa_count[8][34] , \sa_count[8].r.part1[2] );
tran (\sa_count[8][34] , \sa_count[8].f.upper[2] );
tran (\sa_count[8][33] , \sa_count[8].r.part1[1] );
tran (\sa_count[8][33] , \sa_count[8].f.upper[1] );
tran (\sa_count[8][32] , \sa_count[8].r.part1[0] );
tran (\sa_count[8][32] , \sa_count[8].f.upper[0] );
tran (\sa_count[8][31] , \sa_count[8].r.part0[31] );
tran (\sa_count[8][31] , \sa_count[8].f.lower[31] );
tran (\sa_count[8][30] , \sa_count[8].r.part0[30] );
tran (\sa_count[8][30] , \sa_count[8].f.lower[30] );
tran (\sa_count[8][29] , \sa_count[8].r.part0[29] );
tran (\sa_count[8][29] , \sa_count[8].f.lower[29] );
tran (\sa_count[8][28] , \sa_count[8].r.part0[28] );
tran (\sa_count[8][28] , \sa_count[8].f.lower[28] );
tran (\sa_count[8][27] , \sa_count[8].r.part0[27] );
tran (\sa_count[8][27] , \sa_count[8].f.lower[27] );
tran (\sa_count[8][26] , \sa_count[8].r.part0[26] );
tran (\sa_count[8][26] , \sa_count[8].f.lower[26] );
tran (\sa_count[8][25] , \sa_count[8].r.part0[25] );
tran (\sa_count[8][25] , \sa_count[8].f.lower[25] );
tran (\sa_count[8][24] , \sa_count[8].r.part0[24] );
tran (\sa_count[8][24] , \sa_count[8].f.lower[24] );
tran (\sa_count[8][23] , \sa_count[8].r.part0[23] );
tran (\sa_count[8][23] , \sa_count[8].f.lower[23] );
tran (\sa_count[8][22] , \sa_count[8].r.part0[22] );
tran (\sa_count[8][22] , \sa_count[8].f.lower[22] );
tran (\sa_count[8][21] , \sa_count[8].r.part0[21] );
tran (\sa_count[8][21] , \sa_count[8].f.lower[21] );
tran (\sa_count[8][20] , \sa_count[8].r.part0[20] );
tran (\sa_count[8][20] , \sa_count[8].f.lower[20] );
tran (\sa_count[8][19] , \sa_count[8].r.part0[19] );
tran (\sa_count[8][19] , \sa_count[8].f.lower[19] );
tran (\sa_count[8][18] , \sa_count[8].r.part0[18] );
tran (\sa_count[8][18] , \sa_count[8].f.lower[18] );
tran (\sa_count[8][17] , \sa_count[8].r.part0[17] );
tran (\sa_count[8][17] , \sa_count[8].f.lower[17] );
tran (\sa_count[8][16] , \sa_count[8].r.part0[16] );
tran (\sa_count[8][16] , \sa_count[8].f.lower[16] );
tran (\sa_count[8][15] , \sa_count[8].r.part0[15] );
tran (\sa_count[8][15] , \sa_count[8].f.lower[15] );
tran (\sa_count[8][14] , \sa_count[8].r.part0[14] );
tran (\sa_count[8][14] , \sa_count[8].f.lower[14] );
tran (\sa_count[8][13] , \sa_count[8].r.part0[13] );
tran (\sa_count[8][13] , \sa_count[8].f.lower[13] );
tran (\sa_count[8][12] , \sa_count[8].r.part0[12] );
tran (\sa_count[8][12] , \sa_count[8].f.lower[12] );
tran (\sa_count[8][11] , \sa_count[8].r.part0[11] );
tran (\sa_count[8][11] , \sa_count[8].f.lower[11] );
tran (\sa_count[8][10] , \sa_count[8].r.part0[10] );
tran (\sa_count[8][10] , \sa_count[8].f.lower[10] );
tran (\sa_count[8][9] , \sa_count[8].r.part0[9] );
tran (\sa_count[8][9] , \sa_count[8].f.lower[9] );
tran (\sa_count[8][8] , \sa_count[8].r.part0[8] );
tran (\sa_count[8][8] , \sa_count[8].f.lower[8] );
tran (\sa_count[8][7] , \sa_count[8].r.part0[7] );
tran (\sa_count[8][7] , \sa_count[8].f.lower[7] );
tran (\sa_count[8][6] , \sa_count[8].r.part0[6] );
tran (\sa_count[8][6] , \sa_count[8].f.lower[6] );
tran (\sa_count[8][5] , \sa_count[8].r.part0[5] );
tran (\sa_count[8][5] , \sa_count[8].f.lower[5] );
tran (\sa_count[8][4] , \sa_count[8].r.part0[4] );
tran (\sa_count[8][4] , \sa_count[8].f.lower[4] );
tran (\sa_count[8][3] , \sa_count[8].r.part0[3] );
tran (\sa_count[8][3] , \sa_count[8].f.lower[3] );
tran (\sa_count[8][2] , \sa_count[8].r.part0[2] );
tran (\sa_count[8][2] , \sa_count[8].f.lower[2] );
tran (\sa_count[8][1] , \sa_count[8].r.part0[1] );
tran (\sa_count[8][1] , \sa_count[8].f.lower[1] );
tran (\sa_count[8][0] , \sa_count[8].r.part0[0] );
tran (\sa_count[8][0] , \sa_count[8].f.lower[0] );
tran (\sa_count[7][63] , \sa_count[7].r.part1[31] );
tran (\sa_count[7][63] , \sa_count[7].f.unused[13] );
tran (\sa_count[7][62] , \sa_count[7].r.part1[30] );
tran (\sa_count[7][62] , \sa_count[7].f.unused[12] );
tran (\sa_count[7][61] , \sa_count[7].r.part1[29] );
tran (\sa_count[7][61] , \sa_count[7].f.unused[11] );
tran (\sa_count[7][60] , \sa_count[7].r.part1[28] );
tran (\sa_count[7][60] , \sa_count[7].f.unused[10] );
tran (\sa_count[7][59] , \sa_count[7].r.part1[27] );
tran (\sa_count[7][59] , \sa_count[7].f.unused[9] );
tran (\sa_count[7][58] , \sa_count[7].r.part1[26] );
tran (\sa_count[7][58] , \sa_count[7].f.unused[8] );
tran (\sa_count[7][57] , \sa_count[7].r.part1[25] );
tran (\sa_count[7][57] , \sa_count[7].f.unused[7] );
tran (\sa_count[7][56] , \sa_count[7].r.part1[24] );
tran (\sa_count[7][56] , \sa_count[7].f.unused[6] );
tran (\sa_count[7][55] , \sa_count[7].r.part1[23] );
tran (\sa_count[7][55] , \sa_count[7].f.unused[5] );
tran (\sa_count[7][54] , \sa_count[7].r.part1[22] );
tran (\sa_count[7][54] , \sa_count[7].f.unused[4] );
tran (\sa_count[7][53] , \sa_count[7].r.part1[21] );
tran (\sa_count[7][53] , \sa_count[7].f.unused[3] );
tran (\sa_count[7][52] , \sa_count[7].r.part1[20] );
tran (\sa_count[7][52] , \sa_count[7].f.unused[2] );
tran (\sa_count[7][51] , \sa_count[7].r.part1[19] );
tran (\sa_count[7][51] , \sa_count[7].f.unused[1] );
tran (\sa_count[7][50] , \sa_count[7].r.part1[18] );
tran (\sa_count[7][50] , \sa_count[7].f.unused[0] );
tran (\sa_count[7][49] , \sa_count[7].r.part1[17] );
tran (\sa_count[7][49] , \sa_count[7].f.upper[17] );
tran (\sa_count[7][48] , \sa_count[7].r.part1[16] );
tran (\sa_count[7][48] , \sa_count[7].f.upper[16] );
tran (\sa_count[7][47] , \sa_count[7].r.part1[15] );
tran (\sa_count[7][47] , \sa_count[7].f.upper[15] );
tran (\sa_count[7][46] , \sa_count[7].r.part1[14] );
tran (\sa_count[7][46] , \sa_count[7].f.upper[14] );
tran (\sa_count[7][45] , \sa_count[7].r.part1[13] );
tran (\sa_count[7][45] , \sa_count[7].f.upper[13] );
tran (\sa_count[7][44] , \sa_count[7].r.part1[12] );
tran (\sa_count[7][44] , \sa_count[7].f.upper[12] );
tran (\sa_count[7][43] , \sa_count[7].r.part1[11] );
tran (\sa_count[7][43] , \sa_count[7].f.upper[11] );
tran (\sa_count[7][42] , \sa_count[7].r.part1[10] );
tran (\sa_count[7][42] , \sa_count[7].f.upper[10] );
tran (\sa_count[7][41] , \sa_count[7].r.part1[9] );
tran (\sa_count[7][41] , \sa_count[7].f.upper[9] );
tran (\sa_count[7][40] , \sa_count[7].r.part1[8] );
tran (\sa_count[7][40] , \sa_count[7].f.upper[8] );
tran (\sa_count[7][39] , \sa_count[7].r.part1[7] );
tran (\sa_count[7][39] , \sa_count[7].f.upper[7] );
tran (\sa_count[7][38] , \sa_count[7].r.part1[6] );
tran (\sa_count[7][38] , \sa_count[7].f.upper[6] );
tran (\sa_count[7][37] , \sa_count[7].r.part1[5] );
tran (\sa_count[7][37] , \sa_count[7].f.upper[5] );
tran (\sa_count[7][36] , \sa_count[7].r.part1[4] );
tran (\sa_count[7][36] , \sa_count[7].f.upper[4] );
tran (\sa_count[7][35] , \sa_count[7].r.part1[3] );
tran (\sa_count[7][35] , \sa_count[7].f.upper[3] );
tran (\sa_count[7][34] , \sa_count[7].r.part1[2] );
tran (\sa_count[7][34] , \sa_count[7].f.upper[2] );
tran (\sa_count[7][33] , \sa_count[7].r.part1[1] );
tran (\sa_count[7][33] , \sa_count[7].f.upper[1] );
tran (\sa_count[7][32] , \sa_count[7].r.part1[0] );
tran (\sa_count[7][32] , \sa_count[7].f.upper[0] );
tran (\sa_count[7][31] , \sa_count[7].r.part0[31] );
tran (\sa_count[7][31] , \sa_count[7].f.lower[31] );
tran (\sa_count[7][30] , \sa_count[7].r.part0[30] );
tran (\sa_count[7][30] , \sa_count[7].f.lower[30] );
tran (\sa_count[7][29] , \sa_count[7].r.part0[29] );
tran (\sa_count[7][29] , \sa_count[7].f.lower[29] );
tran (\sa_count[7][28] , \sa_count[7].r.part0[28] );
tran (\sa_count[7][28] , \sa_count[7].f.lower[28] );
tran (\sa_count[7][27] , \sa_count[7].r.part0[27] );
tran (\sa_count[7][27] , \sa_count[7].f.lower[27] );
tran (\sa_count[7][26] , \sa_count[7].r.part0[26] );
tran (\sa_count[7][26] , \sa_count[7].f.lower[26] );
tran (\sa_count[7][25] , \sa_count[7].r.part0[25] );
tran (\sa_count[7][25] , \sa_count[7].f.lower[25] );
tran (\sa_count[7][24] , \sa_count[7].r.part0[24] );
tran (\sa_count[7][24] , \sa_count[7].f.lower[24] );
tran (\sa_count[7][23] , \sa_count[7].r.part0[23] );
tran (\sa_count[7][23] , \sa_count[7].f.lower[23] );
tran (\sa_count[7][22] , \sa_count[7].r.part0[22] );
tran (\sa_count[7][22] , \sa_count[7].f.lower[22] );
tran (\sa_count[7][21] , \sa_count[7].r.part0[21] );
tran (\sa_count[7][21] , \sa_count[7].f.lower[21] );
tran (\sa_count[7][20] , \sa_count[7].r.part0[20] );
tran (\sa_count[7][20] , \sa_count[7].f.lower[20] );
tran (\sa_count[7][19] , \sa_count[7].r.part0[19] );
tran (\sa_count[7][19] , \sa_count[7].f.lower[19] );
tran (\sa_count[7][18] , \sa_count[7].r.part0[18] );
tran (\sa_count[7][18] , \sa_count[7].f.lower[18] );
tran (\sa_count[7][17] , \sa_count[7].r.part0[17] );
tran (\sa_count[7][17] , \sa_count[7].f.lower[17] );
tran (\sa_count[7][16] , \sa_count[7].r.part0[16] );
tran (\sa_count[7][16] , \sa_count[7].f.lower[16] );
tran (\sa_count[7][15] , \sa_count[7].r.part0[15] );
tran (\sa_count[7][15] , \sa_count[7].f.lower[15] );
tran (\sa_count[7][14] , \sa_count[7].r.part0[14] );
tran (\sa_count[7][14] , \sa_count[7].f.lower[14] );
tran (\sa_count[7][13] , \sa_count[7].r.part0[13] );
tran (\sa_count[7][13] , \sa_count[7].f.lower[13] );
tran (\sa_count[7][12] , \sa_count[7].r.part0[12] );
tran (\sa_count[7][12] , \sa_count[7].f.lower[12] );
tran (\sa_count[7][11] , \sa_count[7].r.part0[11] );
tran (\sa_count[7][11] , \sa_count[7].f.lower[11] );
tran (\sa_count[7][10] , \sa_count[7].r.part0[10] );
tran (\sa_count[7][10] , \sa_count[7].f.lower[10] );
tran (\sa_count[7][9] , \sa_count[7].r.part0[9] );
tran (\sa_count[7][9] , \sa_count[7].f.lower[9] );
tran (\sa_count[7][8] , \sa_count[7].r.part0[8] );
tran (\sa_count[7][8] , \sa_count[7].f.lower[8] );
tran (\sa_count[7][7] , \sa_count[7].r.part0[7] );
tran (\sa_count[7][7] , \sa_count[7].f.lower[7] );
tran (\sa_count[7][6] , \sa_count[7].r.part0[6] );
tran (\sa_count[7][6] , \sa_count[7].f.lower[6] );
tran (\sa_count[7][5] , \sa_count[7].r.part0[5] );
tran (\sa_count[7][5] , \sa_count[7].f.lower[5] );
tran (\sa_count[7][4] , \sa_count[7].r.part0[4] );
tran (\sa_count[7][4] , \sa_count[7].f.lower[4] );
tran (\sa_count[7][3] , \sa_count[7].r.part0[3] );
tran (\sa_count[7][3] , \sa_count[7].f.lower[3] );
tran (\sa_count[7][2] , \sa_count[7].r.part0[2] );
tran (\sa_count[7][2] , \sa_count[7].f.lower[2] );
tran (\sa_count[7][1] , \sa_count[7].r.part0[1] );
tran (\sa_count[7][1] , \sa_count[7].f.lower[1] );
tran (\sa_count[7][0] , \sa_count[7].r.part0[0] );
tran (\sa_count[7][0] , \sa_count[7].f.lower[0] );
tran (\sa_count[6][63] , \sa_count[6].r.part1[31] );
tran (\sa_count[6][63] , \sa_count[6].f.unused[13] );
tran (\sa_count[6][62] , \sa_count[6].r.part1[30] );
tran (\sa_count[6][62] , \sa_count[6].f.unused[12] );
tran (\sa_count[6][61] , \sa_count[6].r.part1[29] );
tran (\sa_count[6][61] , \sa_count[6].f.unused[11] );
tran (\sa_count[6][60] , \sa_count[6].r.part1[28] );
tran (\sa_count[6][60] , \sa_count[6].f.unused[10] );
tran (\sa_count[6][59] , \sa_count[6].r.part1[27] );
tran (\sa_count[6][59] , \sa_count[6].f.unused[9] );
tran (\sa_count[6][58] , \sa_count[6].r.part1[26] );
tran (\sa_count[6][58] , \sa_count[6].f.unused[8] );
tran (\sa_count[6][57] , \sa_count[6].r.part1[25] );
tran (\sa_count[6][57] , \sa_count[6].f.unused[7] );
tran (\sa_count[6][56] , \sa_count[6].r.part1[24] );
tran (\sa_count[6][56] , \sa_count[6].f.unused[6] );
tran (\sa_count[6][55] , \sa_count[6].r.part1[23] );
tran (\sa_count[6][55] , \sa_count[6].f.unused[5] );
tran (\sa_count[6][54] , \sa_count[6].r.part1[22] );
tran (\sa_count[6][54] , \sa_count[6].f.unused[4] );
tran (\sa_count[6][53] , \sa_count[6].r.part1[21] );
tran (\sa_count[6][53] , \sa_count[6].f.unused[3] );
tran (\sa_count[6][52] , \sa_count[6].r.part1[20] );
tran (\sa_count[6][52] , \sa_count[6].f.unused[2] );
tran (\sa_count[6][51] , \sa_count[6].r.part1[19] );
tran (\sa_count[6][51] , \sa_count[6].f.unused[1] );
tran (\sa_count[6][50] , \sa_count[6].r.part1[18] );
tran (\sa_count[6][50] , \sa_count[6].f.unused[0] );
tran (\sa_count[6][49] , \sa_count[6].r.part1[17] );
tran (\sa_count[6][49] , \sa_count[6].f.upper[17] );
tran (\sa_count[6][48] , \sa_count[6].r.part1[16] );
tran (\sa_count[6][48] , \sa_count[6].f.upper[16] );
tran (\sa_count[6][47] , \sa_count[6].r.part1[15] );
tran (\sa_count[6][47] , \sa_count[6].f.upper[15] );
tran (\sa_count[6][46] , \sa_count[6].r.part1[14] );
tran (\sa_count[6][46] , \sa_count[6].f.upper[14] );
tran (\sa_count[6][45] , \sa_count[6].r.part1[13] );
tran (\sa_count[6][45] , \sa_count[6].f.upper[13] );
tran (\sa_count[6][44] , \sa_count[6].r.part1[12] );
tran (\sa_count[6][44] , \sa_count[6].f.upper[12] );
tran (\sa_count[6][43] , \sa_count[6].r.part1[11] );
tran (\sa_count[6][43] , \sa_count[6].f.upper[11] );
tran (\sa_count[6][42] , \sa_count[6].r.part1[10] );
tran (\sa_count[6][42] , \sa_count[6].f.upper[10] );
tran (\sa_count[6][41] , \sa_count[6].r.part1[9] );
tran (\sa_count[6][41] , \sa_count[6].f.upper[9] );
tran (\sa_count[6][40] , \sa_count[6].r.part1[8] );
tran (\sa_count[6][40] , \sa_count[6].f.upper[8] );
tran (\sa_count[6][39] , \sa_count[6].r.part1[7] );
tran (\sa_count[6][39] , \sa_count[6].f.upper[7] );
tran (\sa_count[6][38] , \sa_count[6].r.part1[6] );
tran (\sa_count[6][38] , \sa_count[6].f.upper[6] );
tran (\sa_count[6][37] , \sa_count[6].r.part1[5] );
tran (\sa_count[6][37] , \sa_count[6].f.upper[5] );
tran (\sa_count[6][36] , \sa_count[6].r.part1[4] );
tran (\sa_count[6][36] , \sa_count[6].f.upper[4] );
tran (\sa_count[6][35] , \sa_count[6].r.part1[3] );
tran (\sa_count[6][35] , \sa_count[6].f.upper[3] );
tran (\sa_count[6][34] , \sa_count[6].r.part1[2] );
tran (\sa_count[6][34] , \sa_count[6].f.upper[2] );
tran (\sa_count[6][33] , \sa_count[6].r.part1[1] );
tran (\sa_count[6][33] , \sa_count[6].f.upper[1] );
tran (\sa_count[6][32] , \sa_count[6].r.part1[0] );
tran (\sa_count[6][32] , \sa_count[6].f.upper[0] );
tran (\sa_count[6][31] , \sa_count[6].r.part0[31] );
tran (\sa_count[6][31] , \sa_count[6].f.lower[31] );
tran (\sa_count[6][30] , \sa_count[6].r.part0[30] );
tran (\sa_count[6][30] , \sa_count[6].f.lower[30] );
tran (\sa_count[6][29] , \sa_count[6].r.part0[29] );
tran (\sa_count[6][29] , \sa_count[6].f.lower[29] );
tran (\sa_count[6][28] , \sa_count[6].r.part0[28] );
tran (\sa_count[6][28] , \sa_count[6].f.lower[28] );
tran (\sa_count[6][27] , \sa_count[6].r.part0[27] );
tran (\sa_count[6][27] , \sa_count[6].f.lower[27] );
tran (\sa_count[6][26] , \sa_count[6].r.part0[26] );
tran (\sa_count[6][26] , \sa_count[6].f.lower[26] );
tran (\sa_count[6][25] , \sa_count[6].r.part0[25] );
tran (\sa_count[6][25] , \sa_count[6].f.lower[25] );
tran (\sa_count[6][24] , \sa_count[6].r.part0[24] );
tran (\sa_count[6][24] , \sa_count[6].f.lower[24] );
tran (\sa_count[6][23] , \sa_count[6].r.part0[23] );
tran (\sa_count[6][23] , \sa_count[6].f.lower[23] );
tran (\sa_count[6][22] , \sa_count[6].r.part0[22] );
tran (\sa_count[6][22] , \sa_count[6].f.lower[22] );
tran (\sa_count[6][21] , \sa_count[6].r.part0[21] );
tran (\sa_count[6][21] , \sa_count[6].f.lower[21] );
tran (\sa_count[6][20] , \sa_count[6].r.part0[20] );
tran (\sa_count[6][20] , \sa_count[6].f.lower[20] );
tran (\sa_count[6][19] , \sa_count[6].r.part0[19] );
tran (\sa_count[6][19] , \sa_count[6].f.lower[19] );
tran (\sa_count[6][18] , \sa_count[6].r.part0[18] );
tran (\sa_count[6][18] , \sa_count[6].f.lower[18] );
tran (\sa_count[6][17] , \sa_count[6].r.part0[17] );
tran (\sa_count[6][17] , \sa_count[6].f.lower[17] );
tran (\sa_count[6][16] , \sa_count[6].r.part0[16] );
tran (\sa_count[6][16] , \sa_count[6].f.lower[16] );
tran (\sa_count[6][15] , \sa_count[6].r.part0[15] );
tran (\sa_count[6][15] , \sa_count[6].f.lower[15] );
tran (\sa_count[6][14] , \sa_count[6].r.part0[14] );
tran (\sa_count[6][14] , \sa_count[6].f.lower[14] );
tran (\sa_count[6][13] , \sa_count[6].r.part0[13] );
tran (\sa_count[6][13] , \sa_count[6].f.lower[13] );
tran (\sa_count[6][12] , \sa_count[6].r.part0[12] );
tran (\sa_count[6][12] , \sa_count[6].f.lower[12] );
tran (\sa_count[6][11] , \sa_count[6].r.part0[11] );
tran (\sa_count[6][11] , \sa_count[6].f.lower[11] );
tran (\sa_count[6][10] , \sa_count[6].r.part0[10] );
tran (\sa_count[6][10] , \sa_count[6].f.lower[10] );
tran (\sa_count[6][9] , \sa_count[6].r.part0[9] );
tran (\sa_count[6][9] , \sa_count[6].f.lower[9] );
tran (\sa_count[6][8] , \sa_count[6].r.part0[8] );
tran (\sa_count[6][8] , \sa_count[6].f.lower[8] );
tran (\sa_count[6][7] , \sa_count[6].r.part0[7] );
tran (\sa_count[6][7] , \sa_count[6].f.lower[7] );
tran (\sa_count[6][6] , \sa_count[6].r.part0[6] );
tran (\sa_count[6][6] , \sa_count[6].f.lower[6] );
tran (\sa_count[6][5] , \sa_count[6].r.part0[5] );
tran (\sa_count[6][5] , \sa_count[6].f.lower[5] );
tran (\sa_count[6][4] , \sa_count[6].r.part0[4] );
tran (\sa_count[6][4] , \sa_count[6].f.lower[4] );
tran (\sa_count[6][3] , \sa_count[6].r.part0[3] );
tran (\sa_count[6][3] , \sa_count[6].f.lower[3] );
tran (\sa_count[6][2] , \sa_count[6].r.part0[2] );
tran (\sa_count[6][2] , \sa_count[6].f.lower[2] );
tran (\sa_count[6][1] , \sa_count[6].r.part0[1] );
tran (\sa_count[6][1] , \sa_count[6].f.lower[1] );
tran (\sa_count[6][0] , \sa_count[6].r.part0[0] );
tran (\sa_count[6][0] , \sa_count[6].f.lower[0] );
tran (\sa_count[5][63] , \sa_count[5].r.part1[31] );
tran (\sa_count[5][63] , \sa_count[5].f.unused[13] );
tran (\sa_count[5][62] , \sa_count[5].r.part1[30] );
tran (\sa_count[5][62] , \sa_count[5].f.unused[12] );
tran (\sa_count[5][61] , \sa_count[5].r.part1[29] );
tran (\sa_count[5][61] , \sa_count[5].f.unused[11] );
tran (\sa_count[5][60] , \sa_count[5].r.part1[28] );
tran (\sa_count[5][60] , \sa_count[5].f.unused[10] );
tran (\sa_count[5][59] , \sa_count[5].r.part1[27] );
tran (\sa_count[5][59] , \sa_count[5].f.unused[9] );
tran (\sa_count[5][58] , \sa_count[5].r.part1[26] );
tran (\sa_count[5][58] , \sa_count[5].f.unused[8] );
tran (\sa_count[5][57] , \sa_count[5].r.part1[25] );
tran (\sa_count[5][57] , \sa_count[5].f.unused[7] );
tran (\sa_count[5][56] , \sa_count[5].r.part1[24] );
tran (\sa_count[5][56] , \sa_count[5].f.unused[6] );
tran (\sa_count[5][55] , \sa_count[5].r.part1[23] );
tran (\sa_count[5][55] , \sa_count[5].f.unused[5] );
tran (\sa_count[5][54] , \sa_count[5].r.part1[22] );
tran (\sa_count[5][54] , \sa_count[5].f.unused[4] );
tran (\sa_count[5][53] , \sa_count[5].r.part1[21] );
tran (\sa_count[5][53] , \sa_count[5].f.unused[3] );
tran (\sa_count[5][52] , \sa_count[5].r.part1[20] );
tran (\sa_count[5][52] , \sa_count[5].f.unused[2] );
tran (\sa_count[5][51] , \sa_count[5].r.part1[19] );
tran (\sa_count[5][51] , \sa_count[5].f.unused[1] );
tran (\sa_count[5][50] , \sa_count[5].r.part1[18] );
tran (\sa_count[5][50] , \sa_count[5].f.unused[0] );
tran (\sa_count[5][49] , \sa_count[5].r.part1[17] );
tran (\sa_count[5][49] , \sa_count[5].f.upper[17] );
tran (\sa_count[5][48] , \sa_count[5].r.part1[16] );
tran (\sa_count[5][48] , \sa_count[5].f.upper[16] );
tran (\sa_count[5][47] , \sa_count[5].r.part1[15] );
tran (\sa_count[5][47] , \sa_count[5].f.upper[15] );
tran (\sa_count[5][46] , \sa_count[5].r.part1[14] );
tran (\sa_count[5][46] , \sa_count[5].f.upper[14] );
tran (\sa_count[5][45] , \sa_count[5].r.part1[13] );
tran (\sa_count[5][45] , \sa_count[5].f.upper[13] );
tran (\sa_count[5][44] , \sa_count[5].r.part1[12] );
tran (\sa_count[5][44] , \sa_count[5].f.upper[12] );
tran (\sa_count[5][43] , \sa_count[5].r.part1[11] );
tran (\sa_count[5][43] , \sa_count[5].f.upper[11] );
tran (\sa_count[5][42] , \sa_count[5].r.part1[10] );
tran (\sa_count[5][42] , \sa_count[5].f.upper[10] );
tran (\sa_count[5][41] , \sa_count[5].r.part1[9] );
tran (\sa_count[5][41] , \sa_count[5].f.upper[9] );
tran (\sa_count[5][40] , \sa_count[5].r.part1[8] );
tran (\sa_count[5][40] , \sa_count[5].f.upper[8] );
tran (\sa_count[5][39] , \sa_count[5].r.part1[7] );
tran (\sa_count[5][39] , \sa_count[5].f.upper[7] );
tran (\sa_count[5][38] , \sa_count[5].r.part1[6] );
tran (\sa_count[5][38] , \sa_count[5].f.upper[6] );
tran (\sa_count[5][37] , \sa_count[5].r.part1[5] );
tran (\sa_count[5][37] , \sa_count[5].f.upper[5] );
tran (\sa_count[5][36] , \sa_count[5].r.part1[4] );
tran (\sa_count[5][36] , \sa_count[5].f.upper[4] );
tran (\sa_count[5][35] , \sa_count[5].r.part1[3] );
tran (\sa_count[5][35] , \sa_count[5].f.upper[3] );
tran (\sa_count[5][34] , \sa_count[5].r.part1[2] );
tran (\sa_count[5][34] , \sa_count[5].f.upper[2] );
tran (\sa_count[5][33] , \sa_count[5].r.part1[1] );
tran (\sa_count[5][33] , \sa_count[5].f.upper[1] );
tran (\sa_count[5][32] , \sa_count[5].r.part1[0] );
tran (\sa_count[5][32] , \sa_count[5].f.upper[0] );
tran (\sa_count[5][31] , \sa_count[5].r.part0[31] );
tran (\sa_count[5][31] , \sa_count[5].f.lower[31] );
tran (\sa_count[5][30] , \sa_count[5].r.part0[30] );
tran (\sa_count[5][30] , \sa_count[5].f.lower[30] );
tran (\sa_count[5][29] , \sa_count[5].r.part0[29] );
tran (\sa_count[5][29] , \sa_count[5].f.lower[29] );
tran (\sa_count[5][28] , \sa_count[5].r.part0[28] );
tran (\sa_count[5][28] , \sa_count[5].f.lower[28] );
tran (\sa_count[5][27] , \sa_count[5].r.part0[27] );
tran (\sa_count[5][27] , \sa_count[5].f.lower[27] );
tran (\sa_count[5][26] , \sa_count[5].r.part0[26] );
tran (\sa_count[5][26] , \sa_count[5].f.lower[26] );
tran (\sa_count[5][25] , \sa_count[5].r.part0[25] );
tran (\sa_count[5][25] , \sa_count[5].f.lower[25] );
tran (\sa_count[5][24] , \sa_count[5].r.part0[24] );
tran (\sa_count[5][24] , \sa_count[5].f.lower[24] );
tran (\sa_count[5][23] , \sa_count[5].r.part0[23] );
tran (\sa_count[5][23] , \sa_count[5].f.lower[23] );
tran (\sa_count[5][22] , \sa_count[5].r.part0[22] );
tran (\sa_count[5][22] , \sa_count[5].f.lower[22] );
tran (\sa_count[5][21] , \sa_count[5].r.part0[21] );
tran (\sa_count[5][21] , \sa_count[5].f.lower[21] );
tran (\sa_count[5][20] , \sa_count[5].r.part0[20] );
tran (\sa_count[5][20] , \sa_count[5].f.lower[20] );
tran (\sa_count[5][19] , \sa_count[5].r.part0[19] );
tran (\sa_count[5][19] , \sa_count[5].f.lower[19] );
tran (\sa_count[5][18] , \sa_count[5].r.part0[18] );
tran (\sa_count[5][18] , \sa_count[5].f.lower[18] );
tran (\sa_count[5][17] , \sa_count[5].r.part0[17] );
tran (\sa_count[5][17] , \sa_count[5].f.lower[17] );
tran (\sa_count[5][16] , \sa_count[5].r.part0[16] );
tran (\sa_count[5][16] , \sa_count[5].f.lower[16] );
tran (\sa_count[5][15] , \sa_count[5].r.part0[15] );
tran (\sa_count[5][15] , \sa_count[5].f.lower[15] );
tran (\sa_count[5][14] , \sa_count[5].r.part0[14] );
tran (\sa_count[5][14] , \sa_count[5].f.lower[14] );
tran (\sa_count[5][13] , \sa_count[5].r.part0[13] );
tran (\sa_count[5][13] , \sa_count[5].f.lower[13] );
tran (\sa_count[5][12] , \sa_count[5].r.part0[12] );
tran (\sa_count[5][12] , \sa_count[5].f.lower[12] );
tran (\sa_count[5][11] , \sa_count[5].r.part0[11] );
tran (\sa_count[5][11] , \sa_count[5].f.lower[11] );
tran (\sa_count[5][10] , \sa_count[5].r.part0[10] );
tran (\sa_count[5][10] , \sa_count[5].f.lower[10] );
tran (\sa_count[5][9] , \sa_count[5].r.part0[9] );
tran (\sa_count[5][9] , \sa_count[5].f.lower[9] );
tran (\sa_count[5][8] , \sa_count[5].r.part0[8] );
tran (\sa_count[5][8] , \sa_count[5].f.lower[8] );
tran (\sa_count[5][7] , \sa_count[5].r.part0[7] );
tran (\sa_count[5][7] , \sa_count[5].f.lower[7] );
tran (\sa_count[5][6] , \sa_count[5].r.part0[6] );
tran (\sa_count[5][6] , \sa_count[5].f.lower[6] );
tran (\sa_count[5][5] , \sa_count[5].r.part0[5] );
tran (\sa_count[5][5] , \sa_count[5].f.lower[5] );
tran (\sa_count[5][4] , \sa_count[5].r.part0[4] );
tran (\sa_count[5][4] , \sa_count[5].f.lower[4] );
tran (\sa_count[5][3] , \sa_count[5].r.part0[3] );
tran (\sa_count[5][3] , \sa_count[5].f.lower[3] );
tran (\sa_count[5][2] , \sa_count[5].r.part0[2] );
tran (\sa_count[5][2] , \sa_count[5].f.lower[2] );
tran (\sa_count[5][1] , \sa_count[5].r.part0[1] );
tran (\sa_count[5][1] , \sa_count[5].f.lower[1] );
tran (\sa_count[5][0] , \sa_count[5].r.part0[0] );
tran (\sa_count[5][0] , \sa_count[5].f.lower[0] );
tran (\sa_count[4][63] , \sa_count[4].r.part1[31] );
tran (\sa_count[4][63] , \sa_count[4].f.unused[13] );
tran (\sa_count[4][62] , \sa_count[4].r.part1[30] );
tran (\sa_count[4][62] , \sa_count[4].f.unused[12] );
tran (\sa_count[4][61] , \sa_count[4].r.part1[29] );
tran (\sa_count[4][61] , \sa_count[4].f.unused[11] );
tran (\sa_count[4][60] , \sa_count[4].r.part1[28] );
tran (\sa_count[4][60] , \sa_count[4].f.unused[10] );
tran (\sa_count[4][59] , \sa_count[4].r.part1[27] );
tran (\sa_count[4][59] , \sa_count[4].f.unused[9] );
tran (\sa_count[4][58] , \sa_count[4].r.part1[26] );
tran (\sa_count[4][58] , \sa_count[4].f.unused[8] );
tran (\sa_count[4][57] , \sa_count[4].r.part1[25] );
tran (\sa_count[4][57] , \sa_count[4].f.unused[7] );
tran (\sa_count[4][56] , \sa_count[4].r.part1[24] );
tran (\sa_count[4][56] , \sa_count[4].f.unused[6] );
tran (\sa_count[4][55] , \sa_count[4].r.part1[23] );
tran (\sa_count[4][55] , \sa_count[4].f.unused[5] );
tran (\sa_count[4][54] , \sa_count[4].r.part1[22] );
tran (\sa_count[4][54] , \sa_count[4].f.unused[4] );
tran (\sa_count[4][53] , \sa_count[4].r.part1[21] );
tran (\sa_count[4][53] , \sa_count[4].f.unused[3] );
tran (\sa_count[4][52] , \sa_count[4].r.part1[20] );
tran (\sa_count[4][52] , \sa_count[4].f.unused[2] );
tran (\sa_count[4][51] , \sa_count[4].r.part1[19] );
tran (\sa_count[4][51] , \sa_count[4].f.unused[1] );
tran (\sa_count[4][50] , \sa_count[4].r.part1[18] );
tran (\sa_count[4][50] , \sa_count[4].f.unused[0] );
tran (\sa_count[4][49] , \sa_count[4].r.part1[17] );
tran (\sa_count[4][49] , \sa_count[4].f.upper[17] );
tran (\sa_count[4][48] , \sa_count[4].r.part1[16] );
tran (\sa_count[4][48] , \sa_count[4].f.upper[16] );
tran (\sa_count[4][47] , \sa_count[4].r.part1[15] );
tran (\sa_count[4][47] , \sa_count[4].f.upper[15] );
tran (\sa_count[4][46] , \sa_count[4].r.part1[14] );
tran (\sa_count[4][46] , \sa_count[4].f.upper[14] );
tran (\sa_count[4][45] , \sa_count[4].r.part1[13] );
tran (\sa_count[4][45] , \sa_count[4].f.upper[13] );
tran (\sa_count[4][44] , \sa_count[4].r.part1[12] );
tran (\sa_count[4][44] , \sa_count[4].f.upper[12] );
tran (\sa_count[4][43] , \sa_count[4].r.part1[11] );
tran (\sa_count[4][43] , \sa_count[4].f.upper[11] );
tran (\sa_count[4][42] , \sa_count[4].r.part1[10] );
tran (\sa_count[4][42] , \sa_count[4].f.upper[10] );
tran (\sa_count[4][41] , \sa_count[4].r.part1[9] );
tran (\sa_count[4][41] , \sa_count[4].f.upper[9] );
tran (\sa_count[4][40] , \sa_count[4].r.part1[8] );
tran (\sa_count[4][40] , \sa_count[4].f.upper[8] );
tran (\sa_count[4][39] , \sa_count[4].r.part1[7] );
tran (\sa_count[4][39] , \sa_count[4].f.upper[7] );
tran (\sa_count[4][38] , \sa_count[4].r.part1[6] );
tran (\sa_count[4][38] , \sa_count[4].f.upper[6] );
tran (\sa_count[4][37] , \sa_count[4].r.part1[5] );
tran (\sa_count[4][37] , \sa_count[4].f.upper[5] );
tran (\sa_count[4][36] , \sa_count[4].r.part1[4] );
tran (\sa_count[4][36] , \sa_count[4].f.upper[4] );
tran (\sa_count[4][35] , \sa_count[4].r.part1[3] );
tran (\sa_count[4][35] , \sa_count[4].f.upper[3] );
tran (\sa_count[4][34] , \sa_count[4].r.part1[2] );
tran (\sa_count[4][34] , \sa_count[4].f.upper[2] );
tran (\sa_count[4][33] , \sa_count[4].r.part1[1] );
tran (\sa_count[4][33] , \sa_count[4].f.upper[1] );
tran (\sa_count[4][32] , \sa_count[4].r.part1[0] );
tran (\sa_count[4][32] , \sa_count[4].f.upper[0] );
tran (\sa_count[4][31] , \sa_count[4].r.part0[31] );
tran (\sa_count[4][31] , \sa_count[4].f.lower[31] );
tran (\sa_count[4][30] , \sa_count[4].r.part0[30] );
tran (\sa_count[4][30] , \sa_count[4].f.lower[30] );
tran (\sa_count[4][29] , \sa_count[4].r.part0[29] );
tran (\sa_count[4][29] , \sa_count[4].f.lower[29] );
tran (\sa_count[4][28] , \sa_count[4].r.part0[28] );
tran (\sa_count[4][28] , \sa_count[4].f.lower[28] );
tran (\sa_count[4][27] , \sa_count[4].r.part0[27] );
tran (\sa_count[4][27] , \sa_count[4].f.lower[27] );
tran (\sa_count[4][26] , \sa_count[4].r.part0[26] );
tran (\sa_count[4][26] , \sa_count[4].f.lower[26] );
tran (\sa_count[4][25] , \sa_count[4].r.part0[25] );
tran (\sa_count[4][25] , \sa_count[4].f.lower[25] );
tran (\sa_count[4][24] , \sa_count[4].r.part0[24] );
tran (\sa_count[4][24] , \sa_count[4].f.lower[24] );
tran (\sa_count[4][23] , \sa_count[4].r.part0[23] );
tran (\sa_count[4][23] , \sa_count[4].f.lower[23] );
tran (\sa_count[4][22] , \sa_count[4].r.part0[22] );
tran (\sa_count[4][22] , \sa_count[4].f.lower[22] );
tran (\sa_count[4][21] , \sa_count[4].r.part0[21] );
tran (\sa_count[4][21] , \sa_count[4].f.lower[21] );
tran (\sa_count[4][20] , \sa_count[4].r.part0[20] );
tran (\sa_count[4][20] , \sa_count[4].f.lower[20] );
tran (\sa_count[4][19] , \sa_count[4].r.part0[19] );
tran (\sa_count[4][19] , \sa_count[4].f.lower[19] );
tran (\sa_count[4][18] , \sa_count[4].r.part0[18] );
tran (\sa_count[4][18] , \sa_count[4].f.lower[18] );
tran (\sa_count[4][17] , \sa_count[4].r.part0[17] );
tran (\sa_count[4][17] , \sa_count[4].f.lower[17] );
tran (\sa_count[4][16] , \sa_count[4].r.part0[16] );
tran (\sa_count[4][16] , \sa_count[4].f.lower[16] );
tran (\sa_count[4][15] , \sa_count[4].r.part0[15] );
tran (\sa_count[4][15] , \sa_count[4].f.lower[15] );
tran (\sa_count[4][14] , \sa_count[4].r.part0[14] );
tran (\sa_count[4][14] , \sa_count[4].f.lower[14] );
tran (\sa_count[4][13] , \sa_count[4].r.part0[13] );
tran (\sa_count[4][13] , \sa_count[4].f.lower[13] );
tran (\sa_count[4][12] , \sa_count[4].r.part0[12] );
tran (\sa_count[4][12] , \sa_count[4].f.lower[12] );
tran (\sa_count[4][11] , \sa_count[4].r.part0[11] );
tran (\sa_count[4][11] , \sa_count[4].f.lower[11] );
tran (\sa_count[4][10] , \sa_count[4].r.part0[10] );
tran (\sa_count[4][10] , \sa_count[4].f.lower[10] );
tran (\sa_count[4][9] , \sa_count[4].r.part0[9] );
tran (\sa_count[4][9] , \sa_count[4].f.lower[9] );
tran (\sa_count[4][8] , \sa_count[4].r.part0[8] );
tran (\sa_count[4][8] , \sa_count[4].f.lower[8] );
tran (\sa_count[4][7] , \sa_count[4].r.part0[7] );
tran (\sa_count[4][7] , \sa_count[4].f.lower[7] );
tran (\sa_count[4][6] , \sa_count[4].r.part0[6] );
tran (\sa_count[4][6] , \sa_count[4].f.lower[6] );
tran (\sa_count[4][5] , \sa_count[4].r.part0[5] );
tran (\sa_count[4][5] , \sa_count[4].f.lower[5] );
tran (\sa_count[4][4] , \sa_count[4].r.part0[4] );
tran (\sa_count[4][4] , \sa_count[4].f.lower[4] );
tran (\sa_count[4][3] , \sa_count[4].r.part0[3] );
tran (\sa_count[4][3] , \sa_count[4].f.lower[3] );
tran (\sa_count[4][2] , \sa_count[4].r.part0[2] );
tran (\sa_count[4][2] , \sa_count[4].f.lower[2] );
tran (\sa_count[4][1] , \sa_count[4].r.part0[1] );
tran (\sa_count[4][1] , \sa_count[4].f.lower[1] );
tran (\sa_count[4][0] , \sa_count[4].r.part0[0] );
tran (\sa_count[4][0] , \sa_count[4].f.lower[0] );
tran (\sa_count[3][63] , \sa_count[3].r.part1[31] );
tran (\sa_count[3][63] , \sa_count[3].f.unused[13] );
tran (\sa_count[3][62] , \sa_count[3].r.part1[30] );
tran (\sa_count[3][62] , \sa_count[3].f.unused[12] );
tran (\sa_count[3][61] , \sa_count[3].r.part1[29] );
tran (\sa_count[3][61] , \sa_count[3].f.unused[11] );
tran (\sa_count[3][60] , \sa_count[3].r.part1[28] );
tran (\sa_count[3][60] , \sa_count[3].f.unused[10] );
tran (\sa_count[3][59] , \sa_count[3].r.part1[27] );
tran (\sa_count[3][59] , \sa_count[3].f.unused[9] );
tran (\sa_count[3][58] , \sa_count[3].r.part1[26] );
tran (\sa_count[3][58] , \sa_count[3].f.unused[8] );
tran (\sa_count[3][57] , \sa_count[3].r.part1[25] );
tran (\sa_count[3][57] , \sa_count[3].f.unused[7] );
tran (\sa_count[3][56] , \sa_count[3].r.part1[24] );
tran (\sa_count[3][56] , \sa_count[3].f.unused[6] );
tran (\sa_count[3][55] , \sa_count[3].r.part1[23] );
tran (\sa_count[3][55] , \sa_count[3].f.unused[5] );
tran (\sa_count[3][54] , \sa_count[3].r.part1[22] );
tran (\sa_count[3][54] , \sa_count[3].f.unused[4] );
tran (\sa_count[3][53] , \sa_count[3].r.part1[21] );
tran (\sa_count[3][53] , \sa_count[3].f.unused[3] );
tran (\sa_count[3][52] , \sa_count[3].r.part1[20] );
tran (\sa_count[3][52] , \sa_count[3].f.unused[2] );
tran (\sa_count[3][51] , \sa_count[3].r.part1[19] );
tran (\sa_count[3][51] , \sa_count[3].f.unused[1] );
tran (\sa_count[3][50] , \sa_count[3].r.part1[18] );
tran (\sa_count[3][50] , \sa_count[3].f.unused[0] );
tran (\sa_count[3][49] , \sa_count[3].r.part1[17] );
tran (\sa_count[3][49] , \sa_count[3].f.upper[17] );
tran (\sa_count[3][48] , \sa_count[3].r.part1[16] );
tran (\sa_count[3][48] , \sa_count[3].f.upper[16] );
tran (\sa_count[3][47] , \sa_count[3].r.part1[15] );
tran (\sa_count[3][47] , \sa_count[3].f.upper[15] );
tran (\sa_count[3][46] , \sa_count[3].r.part1[14] );
tran (\sa_count[3][46] , \sa_count[3].f.upper[14] );
tran (\sa_count[3][45] , \sa_count[3].r.part1[13] );
tran (\sa_count[3][45] , \sa_count[3].f.upper[13] );
tran (\sa_count[3][44] , \sa_count[3].r.part1[12] );
tran (\sa_count[3][44] , \sa_count[3].f.upper[12] );
tran (\sa_count[3][43] , \sa_count[3].r.part1[11] );
tran (\sa_count[3][43] , \sa_count[3].f.upper[11] );
tran (\sa_count[3][42] , \sa_count[3].r.part1[10] );
tran (\sa_count[3][42] , \sa_count[3].f.upper[10] );
tran (\sa_count[3][41] , \sa_count[3].r.part1[9] );
tran (\sa_count[3][41] , \sa_count[3].f.upper[9] );
tran (\sa_count[3][40] , \sa_count[3].r.part1[8] );
tran (\sa_count[3][40] , \sa_count[3].f.upper[8] );
tran (\sa_count[3][39] , \sa_count[3].r.part1[7] );
tran (\sa_count[3][39] , \sa_count[3].f.upper[7] );
tran (\sa_count[3][38] , \sa_count[3].r.part1[6] );
tran (\sa_count[3][38] , \sa_count[3].f.upper[6] );
tran (\sa_count[3][37] , \sa_count[3].r.part1[5] );
tran (\sa_count[3][37] , \sa_count[3].f.upper[5] );
tran (\sa_count[3][36] , \sa_count[3].r.part1[4] );
tran (\sa_count[3][36] , \sa_count[3].f.upper[4] );
tran (\sa_count[3][35] , \sa_count[3].r.part1[3] );
tran (\sa_count[3][35] , \sa_count[3].f.upper[3] );
tran (\sa_count[3][34] , \sa_count[3].r.part1[2] );
tran (\sa_count[3][34] , \sa_count[3].f.upper[2] );
tran (\sa_count[3][33] , \sa_count[3].r.part1[1] );
tran (\sa_count[3][33] , \sa_count[3].f.upper[1] );
tran (\sa_count[3][32] , \sa_count[3].r.part1[0] );
tran (\sa_count[3][32] , \sa_count[3].f.upper[0] );
tran (\sa_count[3][31] , \sa_count[3].r.part0[31] );
tran (\sa_count[3][31] , \sa_count[3].f.lower[31] );
tran (\sa_count[3][30] , \sa_count[3].r.part0[30] );
tran (\sa_count[3][30] , \sa_count[3].f.lower[30] );
tran (\sa_count[3][29] , \sa_count[3].r.part0[29] );
tran (\sa_count[3][29] , \sa_count[3].f.lower[29] );
tran (\sa_count[3][28] , \sa_count[3].r.part0[28] );
tran (\sa_count[3][28] , \sa_count[3].f.lower[28] );
tran (\sa_count[3][27] , \sa_count[3].r.part0[27] );
tran (\sa_count[3][27] , \sa_count[3].f.lower[27] );
tran (\sa_count[3][26] , \sa_count[3].r.part0[26] );
tran (\sa_count[3][26] , \sa_count[3].f.lower[26] );
tran (\sa_count[3][25] , \sa_count[3].r.part0[25] );
tran (\sa_count[3][25] , \sa_count[3].f.lower[25] );
tran (\sa_count[3][24] , \sa_count[3].r.part0[24] );
tran (\sa_count[3][24] , \sa_count[3].f.lower[24] );
tran (\sa_count[3][23] , \sa_count[3].r.part0[23] );
tran (\sa_count[3][23] , \sa_count[3].f.lower[23] );
tran (\sa_count[3][22] , \sa_count[3].r.part0[22] );
tran (\sa_count[3][22] , \sa_count[3].f.lower[22] );
tran (\sa_count[3][21] , \sa_count[3].r.part0[21] );
tran (\sa_count[3][21] , \sa_count[3].f.lower[21] );
tran (\sa_count[3][20] , \sa_count[3].r.part0[20] );
tran (\sa_count[3][20] , \sa_count[3].f.lower[20] );
tran (\sa_count[3][19] , \sa_count[3].r.part0[19] );
tran (\sa_count[3][19] , \sa_count[3].f.lower[19] );
tran (\sa_count[3][18] , \sa_count[3].r.part0[18] );
tran (\sa_count[3][18] , \sa_count[3].f.lower[18] );
tran (\sa_count[3][17] , \sa_count[3].r.part0[17] );
tran (\sa_count[3][17] , \sa_count[3].f.lower[17] );
tran (\sa_count[3][16] , \sa_count[3].r.part0[16] );
tran (\sa_count[3][16] , \sa_count[3].f.lower[16] );
tran (\sa_count[3][15] , \sa_count[3].r.part0[15] );
tran (\sa_count[3][15] , \sa_count[3].f.lower[15] );
tran (\sa_count[3][14] , \sa_count[3].r.part0[14] );
tran (\sa_count[3][14] , \sa_count[3].f.lower[14] );
tran (\sa_count[3][13] , \sa_count[3].r.part0[13] );
tran (\sa_count[3][13] , \sa_count[3].f.lower[13] );
tran (\sa_count[3][12] , \sa_count[3].r.part0[12] );
tran (\sa_count[3][12] , \sa_count[3].f.lower[12] );
tran (\sa_count[3][11] , \sa_count[3].r.part0[11] );
tran (\sa_count[3][11] , \sa_count[3].f.lower[11] );
tran (\sa_count[3][10] , \sa_count[3].r.part0[10] );
tran (\sa_count[3][10] , \sa_count[3].f.lower[10] );
tran (\sa_count[3][9] , \sa_count[3].r.part0[9] );
tran (\sa_count[3][9] , \sa_count[3].f.lower[9] );
tran (\sa_count[3][8] , \sa_count[3].r.part0[8] );
tran (\sa_count[3][8] , \sa_count[3].f.lower[8] );
tran (\sa_count[3][7] , \sa_count[3].r.part0[7] );
tran (\sa_count[3][7] , \sa_count[3].f.lower[7] );
tran (\sa_count[3][6] , \sa_count[3].r.part0[6] );
tran (\sa_count[3][6] , \sa_count[3].f.lower[6] );
tran (\sa_count[3][5] , \sa_count[3].r.part0[5] );
tran (\sa_count[3][5] , \sa_count[3].f.lower[5] );
tran (\sa_count[3][4] , \sa_count[3].r.part0[4] );
tran (\sa_count[3][4] , \sa_count[3].f.lower[4] );
tran (\sa_count[3][3] , \sa_count[3].r.part0[3] );
tran (\sa_count[3][3] , \sa_count[3].f.lower[3] );
tran (\sa_count[3][2] , \sa_count[3].r.part0[2] );
tran (\sa_count[3][2] , \sa_count[3].f.lower[2] );
tran (\sa_count[3][1] , \sa_count[3].r.part0[1] );
tran (\sa_count[3][1] , \sa_count[3].f.lower[1] );
tran (\sa_count[3][0] , \sa_count[3].r.part0[0] );
tran (\sa_count[3][0] , \sa_count[3].f.lower[0] );
tran (\sa_count[2][63] , \sa_count[2].r.part1[31] );
tran (\sa_count[2][63] , \sa_count[2].f.unused[13] );
tran (\sa_count[2][62] , \sa_count[2].r.part1[30] );
tran (\sa_count[2][62] , \sa_count[2].f.unused[12] );
tran (\sa_count[2][61] , \sa_count[2].r.part1[29] );
tran (\sa_count[2][61] , \sa_count[2].f.unused[11] );
tran (\sa_count[2][60] , \sa_count[2].r.part1[28] );
tran (\sa_count[2][60] , \sa_count[2].f.unused[10] );
tran (\sa_count[2][59] , \sa_count[2].r.part1[27] );
tran (\sa_count[2][59] , \sa_count[2].f.unused[9] );
tran (\sa_count[2][58] , \sa_count[2].r.part1[26] );
tran (\sa_count[2][58] , \sa_count[2].f.unused[8] );
tran (\sa_count[2][57] , \sa_count[2].r.part1[25] );
tran (\sa_count[2][57] , \sa_count[2].f.unused[7] );
tran (\sa_count[2][56] , \sa_count[2].r.part1[24] );
tran (\sa_count[2][56] , \sa_count[2].f.unused[6] );
tran (\sa_count[2][55] , \sa_count[2].r.part1[23] );
tran (\sa_count[2][55] , \sa_count[2].f.unused[5] );
tran (\sa_count[2][54] , \sa_count[2].r.part1[22] );
tran (\sa_count[2][54] , \sa_count[2].f.unused[4] );
tran (\sa_count[2][53] , \sa_count[2].r.part1[21] );
tran (\sa_count[2][53] , \sa_count[2].f.unused[3] );
tran (\sa_count[2][52] , \sa_count[2].r.part1[20] );
tran (\sa_count[2][52] , \sa_count[2].f.unused[2] );
tran (\sa_count[2][51] , \sa_count[2].r.part1[19] );
tran (\sa_count[2][51] , \sa_count[2].f.unused[1] );
tran (\sa_count[2][50] , \sa_count[2].r.part1[18] );
tran (\sa_count[2][50] , \sa_count[2].f.unused[0] );
tran (\sa_count[2][49] , \sa_count[2].r.part1[17] );
tran (\sa_count[2][49] , \sa_count[2].f.upper[17] );
tran (\sa_count[2][48] , \sa_count[2].r.part1[16] );
tran (\sa_count[2][48] , \sa_count[2].f.upper[16] );
tran (\sa_count[2][47] , \sa_count[2].r.part1[15] );
tran (\sa_count[2][47] , \sa_count[2].f.upper[15] );
tran (\sa_count[2][46] , \sa_count[2].r.part1[14] );
tran (\sa_count[2][46] , \sa_count[2].f.upper[14] );
tran (\sa_count[2][45] , \sa_count[2].r.part1[13] );
tran (\sa_count[2][45] , \sa_count[2].f.upper[13] );
tran (\sa_count[2][44] , \sa_count[2].r.part1[12] );
tran (\sa_count[2][44] , \sa_count[2].f.upper[12] );
tran (\sa_count[2][43] , \sa_count[2].r.part1[11] );
tran (\sa_count[2][43] , \sa_count[2].f.upper[11] );
tran (\sa_count[2][42] , \sa_count[2].r.part1[10] );
tran (\sa_count[2][42] , \sa_count[2].f.upper[10] );
tran (\sa_count[2][41] , \sa_count[2].r.part1[9] );
tran (\sa_count[2][41] , \sa_count[2].f.upper[9] );
tran (\sa_count[2][40] , \sa_count[2].r.part1[8] );
tran (\sa_count[2][40] , \sa_count[2].f.upper[8] );
tran (\sa_count[2][39] , \sa_count[2].r.part1[7] );
tran (\sa_count[2][39] , \sa_count[2].f.upper[7] );
tran (\sa_count[2][38] , \sa_count[2].r.part1[6] );
tran (\sa_count[2][38] , \sa_count[2].f.upper[6] );
tran (\sa_count[2][37] , \sa_count[2].r.part1[5] );
tran (\sa_count[2][37] , \sa_count[2].f.upper[5] );
tran (\sa_count[2][36] , \sa_count[2].r.part1[4] );
tran (\sa_count[2][36] , \sa_count[2].f.upper[4] );
tran (\sa_count[2][35] , \sa_count[2].r.part1[3] );
tran (\sa_count[2][35] , \sa_count[2].f.upper[3] );
tran (\sa_count[2][34] , \sa_count[2].r.part1[2] );
tran (\sa_count[2][34] , \sa_count[2].f.upper[2] );
tran (\sa_count[2][33] , \sa_count[2].r.part1[1] );
tran (\sa_count[2][33] , \sa_count[2].f.upper[1] );
tran (\sa_count[2][32] , \sa_count[2].r.part1[0] );
tran (\sa_count[2][32] , \sa_count[2].f.upper[0] );
tran (\sa_count[2][31] , \sa_count[2].r.part0[31] );
tran (\sa_count[2][31] , \sa_count[2].f.lower[31] );
tran (\sa_count[2][30] , \sa_count[2].r.part0[30] );
tran (\sa_count[2][30] , \sa_count[2].f.lower[30] );
tran (\sa_count[2][29] , \sa_count[2].r.part0[29] );
tran (\sa_count[2][29] , \sa_count[2].f.lower[29] );
tran (\sa_count[2][28] , \sa_count[2].r.part0[28] );
tran (\sa_count[2][28] , \sa_count[2].f.lower[28] );
tran (\sa_count[2][27] , \sa_count[2].r.part0[27] );
tran (\sa_count[2][27] , \sa_count[2].f.lower[27] );
tran (\sa_count[2][26] , \sa_count[2].r.part0[26] );
tran (\sa_count[2][26] , \sa_count[2].f.lower[26] );
tran (\sa_count[2][25] , \sa_count[2].r.part0[25] );
tran (\sa_count[2][25] , \sa_count[2].f.lower[25] );
tran (\sa_count[2][24] , \sa_count[2].r.part0[24] );
tran (\sa_count[2][24] , \sa_count[2].f.lower[24] );
tran (\sa_count[2][23] , \sa_count[2].r.part0[23] );
tran (\sa_count[2][23] , \sa_count[2].f.lower[23] );
tran (\sa_count[2][22] , \sa_count[2].r.part0[22] );
tran (\sa_count[2][22] , \sa_count[2].f.lower[22] );
tran (\sa_count[2][21] , \sa_count[2].r.part0[21] );
tran (\sa_count[2][21] , \sa_count[2].f.lower[21] );
tran (\sa_count[2][20] , \sa_count[2].r.part0[20] );
tran (\sa_count[2][20] , \sa_count[2].f.lower[20] );
tran (\sa_count[2][19] , \sa_count[2].r.part0[19] );
tran (\sa_count[2][19] , \sa_count[2].f.lower[19] );
tran (\sa_count[2][18] , \sa_count[2].r.part0[18] );
tran (\sa_count[2][18] , \sa_count[2].f.lower[18] );
tran (\sa_count[2][17] , \sa_count[2].r.part0[17] );
tran (\sa_count[2][17] , \sa_count[2].f.lower[17] );
tran (\sa_count[2][16] , \sa_count[2].r.part0[16] );
tran (\sa_count[2][16] , \sa_count[2].f.lower[16] );
tran (\sa_count[2][15] , \sa_count[2].r.part0[15] );
tran (\sa_count[2][15] , \sa_count[2].f.lower[15] );
tran (\sa_count[2][14] , \sa_count[2].r.part0[14] );
tran (\sa_count[2][14] , \sa_count[2].f.lower[14] );
tran (\sa_count[2][13] , \sa_count[2].r.part0[13] );
tran (\sa_count[2][13] , \sa_count[2].f.lower[13] );
tran (\sa_count[2][12] , \sa_count[2].r.part0[12] );
tran (\sa_count[2][12] , \sa_count[2].f.lower[12] );
tran (\sa_count[2][11] , \sa_count[2].r.part0[11] );
tran (\sa_count[2][11] , \sa_count[2].f.lower[11] );
tran (\sa_count[2][10] , \sa_count[2].r.part0[10] );
tran (\sa_count[2][10] , \sa_count[2].f.lower[10] );
tran (\sa_count[2][9] , \sa_count[2].r.part0[9] );
tran (\sa_count[2][9] , \sa_count[2].f.lower[9] );
tran (\sa_count[2][8] , \sa_count[2].r.part0[8] );
tran (\sa_count[2][8] , \sa_count[2].f.lower[8] );
tran (\sa_count[2][7] , \sa_count[2].r.part0[7] );
tran (\sa_count[2][7] , \sa_count[2].f.lower[7] );
tran (\sa_count[2][6] , \sa_count[2].r.part0[6] );
tran (\sa_count[2][6] , \sa_count[2].f.lower[6] );
tran (\sa_count[2][5] , \sa_count[2].r.part0[5] );
tran (\sa_count[2][5] , \sa_count[2].f.lower[5] );
tran (\sa_count[2][4] , \sa_count[2].r.part0[4] );
tran (\sa_count[2][4] , \sa_count[2].f.lower[4] );
tran (\sa_count[2][3] , \sa_count[2].r.part0[3] );
tran (\sa_count[2][3] , \sa_count[2].f.lower[3] );
tran (\sa_count[2][2] , \sa_count[2].r.part0[2] );
tran (\sa_count[2][2] , \sa_count[2].f.lower[2] );
tran (\sa_count[2][1] , \sa_count[2].r.part0[1] );
tran (\sa_count[2][1] , \sa_count[2].f.lower[1] );
tran (\sa_count[2][0] , \sa_count[2].r.part0[0] );
tran (\sa_count[2][0] , \sa_count[2].f.lower[0] );
tran (\sa_count[1][63] , \sa_count[1].r.part1[31] );
tran (\sa_count[1][63] , \sa_count[1].f.unused[13] );
tran (\sa_count[1][62] , \sa_count[1].r.part1[30] );
tran (\sa_count[1][62] , \sa_count[1].f.unused[12] );
tran (\sa_count[1][61] , \sa_count[1].r.part1[29] );
tran (\sa_count[1][61] , \sa_count[1].f.unused[11] );
tran (\sa_count[1][60] , \sa_count[1].r.part1[28] );
tran (\sa_count[1][60] , \sa_count[1].f.unused[10] );
tran (\sa_count[1][59] , \sa_count[1].r.part1[27] );
tran (\sa_count[1][59] , \sa_count[1].f.unused[9] );
tran (\sa_count[1][58] , \sa_count[1].r.part1[26] );
tran (\sa_count[1][58] , \sa_count[1].f.unused[8] );
tran (\sa_count[1][57] , \sa_count[1].r.part1[25] );
tran (\sa_count[1][57] , \sa_count[1].f.unused[7] );
tran (\sa_count[1][56] , \sa_count[1].r.part1[24] );
tran (\sa_count[1][56] , \sa_count[1].f.unused[6] );
tran (\sa_count[1][55] , \sa_count[1].r.part1[23] );
tran (\sa_count[1][55] , \sa_count[1].f.unused[5] );
tran (\sa_count[1][54] , \sa_count[1].r.part1[22] );
tran (\sa_count[1][54] , \sa_count[1].f.unused[4] );
tran (\sa_count[1][53] , \sa_count[1].r.part1[21] );
tran (\sa_count[1][53] , \sa_count[1].f.unused[3] );
tran (\sa_count[1][52] , \sa_count[1].r.part1[20] );
tran (\sa_count[1][52] , \sa_count[1].f.unused[2] );
tran (\sa_count[1][51] , \sa_count[1].r.part1[19] );
tran (\sa_count[1][51] , \sa_count[1].f.unused[1] );
tran (\sa_count[1][50] , \sa_count[1].r.part1[18] );
tran (\sa_count[1][50] , \sa_count[1].f.unused[0] );
tran (\sa_count[1][49] , \sa_count[1].r.part1[17] );
tran (\sa_count[1][49] , \sa_count[1].f.upper[17] );
tran (\sa_count[1][48] , \sa_count[1].r.part1[16] );
tran (\sa_count[1][48] , \sa_count[1].f.upper[16] );
tran (\sa_count[1][47] , \sa_count[1].r.part1[15] );
tran (\sa_count[1][47] , \sa_count[1].f.upper[15] );
tran (\sa_count[1][46] , \sa_count[1].r.part1[14] );
tran (\sa_count[1][46] , \sa_count[1].f.upper[14] );
tran (\sa_count[1][45] , \sa_count[1].r.part1[13] );
tran (\sa_count[1][45] , \sa_count[1].f.upper[13] );
tran (\sa_count[1][44] , \sa_count[1].r.part1[12] );
tran (\sa_count[1][44] , \sa_count[1].f.upper[12] );
tran (\sa_count[1][43] , \sa_count[1].r.part1[11] );
tran (\sa_count[1][43] , \sa_count[1].f.upper[11] );
tran (\sa_count[1][42] , \sa_count[1].r.part1[10] );
tran (\sa_count[1][42] , \sa_count[1].f.upper[10] );
tran (\sa_count[1][41] , \sa_count[1].r.part1[9] );
tran (\sa_count[1][41] , \sa_count[1].f.upper[9] );
tran (\sa_count[1][40] , \sa_count[1].r.part1[8] );
tran (\sa_count[1][40] , \sa_count[1].f.upper[8] );
tran (\sa_count[1][39] , \sa_count[1].r.part1[7] );
tran (\sa_count[1][39] , \sa_count[1].f.upper[7] );
tran (\sa_count[1][38] , \sa_count[1].r.part1[6] );
tran (\sa_count[1][38] , \sa_count[1].f.upper[6] );
tran (\sa_count[1][37] , \sa_count[1].r.part1[5] );
tran (\sa_count[1][37] , \sa_count[1].f.upper[5] );
tran (\sa_count[1][36] , \sa_count[1].r.part1[4] );
tran (\sa_count[1][36] , \sa_count[1].f.upper[4] );
tran (\sa_count[1][35] , \sa_count[1].r.part1[3] );
tran (\sa_count[1][35] , \sa_count[1].f.upper[3] );
tran (\sa_count[1][34] , \sa_count[1].r.part1[2] );
tran (\sa_count[1][34] , \sa_count[1].f.upper[2] );
tran (\sa_count[1][33] , \sa_count[1].r.part1[1] );
tran (\sa_count[1][33] , \sa_count[1].f.upper[1] );
tran (\sa_count[1][32] , \sa_count[1].r.part1[0] );
tran (\sa_count[1][32] , \sa_count[1].f.upper[0] );
tran (\sa_count[1][31] , \sa_count[1].r.part0[31] );
tran (\sa_count[1][31] , \sa_count[1].f.lower[31] );
tran (\sa_count[1][30] , \sa_count[1].r.part0[30] );
tran (\sa_count[1][30] , \sa_count[1].f.lower[30] );
tran (\sa_count[1][29] , \sa_count[1].r.part0[29] );
tran (\sa_count[1][29] , \sa_count[1].f.lower[29] );
tran (\sa_count[1][28] , \sa_count[1].r.part0[28] );
tran (\sa_count[1][28] , \sa_count[1].f.lower[28] );
tran (\sa_count[1][27] , \sa_count[1].r.part0[27] );
tran (\sa_count[1][27] , \sa_count[1].f.lower[27] );
tran (\sa_count[1][26] , \sa_count[1].r.part0[26] );
tran (\sa_count[1][26] , \sa_count[1].f.lower[26] );
tran (\sa_count[1][25] , \sa_count[1].r.part0[25] );
tran (\sa_count[1][25] , \sa_count[1].f.lower[25] );
tran (\sa_count[1][24] , \sa_count[1].r.part0[24] );
tran (\sa_count[1][24] , \sa_count[1].f.lower[24] );
tran (\sa_count[1][23] , \sa_count[1].r.part0[23] );
tran (\sa_count[1][23] , \sa_count[1].f.lower[23] );
tran (\sa_count[1][22] , \sa_count[1].r.part0[22] );
tran (\sa_count[1][22] , \sa_count[1].f.lower[22] );
tran (\sa_count[1][21] , \sa_count[1].r.part0[21] );
tran (\sa_count[1][21] , \sa_count[1].f.lower[21] );
tran (\sa_count[1][20] , \sa_count[1].r.part0[20] );
tran (\sa_count[1][20] , \sa_count[1].f.lower[20] );
tran (\sa_count[1][19] , \sa_count[1].r.part0[19] );
tran (\sa_count[1][19] , \sa_count[1].f.lower[19] );
tran (\sa_count[1][18] , \sa_count[1].r.part0[18] );
tran (\sa_count[1][18] , \sa_count[1].f.lower[18] );
tran (\sa_count[1][17] , \sa_count[1].r.part0[17] );
tran (\sa_count[1][17] , \sa_count[1].f.lower[17] );
tran (\sa_count[1][16] , \sa_count[1].r.part0[16] );
tran (\sa_count[1][16] , \sa_count[1].f.lower[16] );
tran (\sa_count[1][15] , \sa_count[1].r.part0[15] );
tran (\sa_count[1][15] , \sa_count[1].f.lower[15] );
tran (\sa_count[1][14] , \sa_count[1].r.part0[14] );
tran (\sa_count[1][14] , \sa_count[1].f.lower[14] );
tran (\sa_count[1][13] , \sa_count[1].r.part0[13] );
tran (\sa_count[1][13] , \sa_count[1].f.lower[13] );
tran (\sa_count[1][12] , \sa_count[1].r.part0[12] );
tran (\sa_count[1][12] , \sa_count[1].f.lower[12] );
tran (\sa_count[1][11] , \sa_count[1].r.part0[11] );
tran (\sa_count[1][11] , \sa_count[1].f.lower[11] );
tran (\sa_count[1][10] , \sa_count[1].r.part0[10] );
tran (\sa_count[1][10] , \sa_count[1].f.lower[10] );
tran (\sa_count[1][9] , \sa_count[1].r.part0[9] );
tran (\sa_count[1][9] , \sa_count[1].f.lower[9] );
tran (\sa_count[1][8] , \sa_count[1].r.part0[8] );
tran (\sa_count[1][8] , \sa_count[1].f.lower[8] );
tran (\sa_count[1][7] , \sa_count[1].r.part0[7] );
tran (\sa_count[1][7] , \sa_count[1].f.lower[7] );
tran (\sa_count[1][6] , \sa_count[1].r.part0[6] );
tran (\sa_count[1][6] , \sa_count[1].f.lower[6] );
tran (\sa_count[1][5] , \sa_count[1].r.part0[5] );
tran (\sa_count[1][5] , \sa_count[1].f.lower[5] );
tran (\sa_count[1][4] , \sa_count[1].r.part0[4] );
tran (\sa_count[1][4] , \sa_count[1].f.lower[4] );
tran (\sa_count[1][3] , \sa_count[1].r.part0[3] );
tran (\sa_count[1][3] , \sa_count[1].f.lower[3] );
tran (\sa_count[1][2] , \sa_count[1].r.part0[2] );
tran (\sa_count[1][2] , \sa_count[1].f.lower[2] );
tran (\sa_count[1][1] , \sa_count[1].r.part0[1] );
tran (\sa_count[1][1] , \sa_count[1].f.lower[1] );
tran (\sa_count[1][0] , \sa_count[1].r.part0[0] );
tran (\sa_count[1][0] , \sa_count[1].f.lower[0] );
tran (\sa_count[0][63] , \sa_count[0].r.part1[31] );
tran (\sa_count[0][63] , \sa_count[0].f.unused[13] );
tran (\sa_count[0][62] , \sa_count[0].r.part1[30] );
tran (\sa_count[0][62] , \sa_count[0].f.unused[12] );
tran (\sa_count[0][61] , \sa_count[0].r.part1[29] );
tran (\sa_count[0][61] , \sa_count[0].f.unused[11] );
tran (\sa_count[0][60] , \sa_count[0].r.part1[28] );
tran (\sa_count[0][60] , \sa_count[0].f.unused[10] );
tran (\sa_count[0][59] , \sa_count[0].r.part1[27] );
tran (\sa_count[0][59] , \sa_count[0].f.unused[9] );
tran (\sa_count[0][58] , \sa_count[0].r.part1[26] );
tran (\sa_count[0][58] , \sa_count[0].f.unused[8] );
tran (\sa_count[0][57] , \sa_count[0].r.part1[25] );
tran (\sa_count[0][57] , \sa_count[0].f.unused[7] );
tran (\sa_count[0][56] , \sa_count[0].r.part1[24] );
tran (\sa_count[0][56] , \sa_count[0].f.unused[6] );
tran (\sa_count[0][55] , \sa_count[0].r.part1[23] );
tran (\sa_count[0][55] , \sa_count[0].f.unused[5] );
tran (\sa_count[0][54] , \sa_count[0].r.part1[22] );
tran (\sa_count[0][54] , \sa_count[0].f.unused[4] );
tran (\sa_count[0][53] , \sa_count[0].r.part1[21] );
tran (\sa_count[0][53] , \sa_count[0].f.unused[3] );
tran (\sa_count[0][52] , \sa_count[0].r.part1[20] );
tran (\sa_count[0][52] , \sa_count[0].f.unused[2] );
tran (\sa_count[0][51] , \sa_count[0].r.part1[19] );
tran (\sa_count[0][51] , \sa_count[0].f.unused[1] );
tran (\sa_count[0][50] , \sa_count[0].r.part1[18] );
tran (\sa_count[0][50] , \sa_count[0].f.unused[0] );
tran (\sa_count[0][49] , \sa_count[0].r.part1[17] );
tran (\sa_count[0][49] , \sa_count[0].f.upper[17] );
tran (\sa_count[0][48] , \sa_count[0].r.part1[16] );
tran (\sa_count[0][48] , \sa_count[0].f.upper[16] );
tran (\sa_count[0][47] , \sa_count[0].r.part1[15] );
tran (\sa_count[0][47] , \sa_count[0].f.upper[15] );
tran (\sa_count[0][46] , \sa_count[0].r.part1[14] );
tran (\sa_count[0][46] , \sa_count[0].f.upper[14] );
tran (\sa_count[0][45] , \sa_count[0].r.part1[13] );
tran (\sa_count[0][45] , \sa_count[0].f.upper[13] );
tran (\sa_count[0][44] , \sa_count[0].r.part1[12] );
tran (\sa_count[0][44] , \sa_count[0].f.upper[12] );
tran (\sa_count[0][43] , \sa_count[0].r.part1[11] );
tran (\sa_count[0][43] , \sa_count[0].f.upper[11] );
tran (\sa_count[0][42] , \sa_count[0].r.part1[10] );
tran (\sa_count[0][42] , \sa_count[0].f.upper[10] );
tran (\sa_count[0][41] , \sa_count[0].r.part1[9] );
tran (\sa_count[0][41] , \sa_count[0].f.upper[9] );
tran (\sa_count[0][40] , \sa_count[0].r.part1[8] );
tran (\sa_count[0][40] , \sa_count[0].f.upper[8] );
tran (\sa_count[0][39] , \sa_count[0].r.part1[7] );
tran (\sa_count[0][39] , \sa_count[0].f.upper[7] );
tran (\sa_count[0][38] , \sa_count[0].r.part1[6] );
tran (\sa_count[0][38] , \sa_count[0].f.upper[6] );
tran (\sa_count[0][37] , \sa_count[0].r.part1[5] );
tran (\sa_count[0][37] , \sa_count[0].f.upper[5] );
tran (\sa_count[0][36] , \sa_count[0].r.part1[4] );
tran (\sa_count[0][36] , \sa_count[0].f.upper[4] );
tran (\sa_count[0][35] , \sa_count[0].r.part1[3] );
tran (\sa_count[0][35] , \sa_count[0].f.upper[3] );
tran (\sa_count[0][34] , \sa_count[0].r.part1[2] );
tran (\sa_count[0][34] , \sa_count[0].f.upper[2] );
tran (\sa_count[0][33] , \sa_count[0].r.part1[1] );
tran (\sa_count[0][33] , \sa_count[0].f.upper[1] );
tran (\sa_count[0][32] , \sa_count[0].r.part1[0] );
tran (\sa_count[0][32] , \sa_count[0].f.upper[0] );
tran (\sa_count[0][31] , \sa_count[0].r.part0[31] );
tran (\sa_count[0][31] , \sa_count[0].f.lower[31] );
tran (\sa_count[0][30] , \sa_count[0].r.part0[30] );
tran (\sa_count[0][30] , \sa_count[0].f.lower[30] );
tran (\sa_count[0][29] , \sa_count[0].r.part0[29] );
tran (\sa_count[0][29] , \sa_count[0].f.lower[29] );
tran (\sa_count[0][28] , \sa_count[0].r.part0[28] );
tran (\sa_count[0][28] , \sa_count[0].f.lower[28] );
tran (\sa_count[0][27] , \sa_count[0].r.part0[27] );
tran (\sa_count[0][27] , \sa_count[0].f.lower[27] );
tran (\sa_count[0][26] , \sa_count[0].r.part0[26] );
tran (\sa_count[0][26] , \sa_count[0].f.lower[26] );
tran (\sa_count[0][25] , \sa_count[0].r.part0[25] );
tran (\sa_count[0][25] , \sa_count[0].f.lower[25] );
tran (\sa_count[0][24] , \sa_count[0].r.part0[24] );
tran (\sa_count[0][24] , \sa_count[0].f.lower[24] );
tran (\sa_count[0][23] , \sa_count[0].r.part0[23] );
tran (\sa_count[0][23] , \sa_count[0].f.lower[23] );
tran (\sa_count[0][22] , \sa_count[0].r.part0[22] );
tran (\sa_count[0][22] , \sa_count[0].f.lower[22] );
tran (\sa_count[0][21] , \sa_count[0].r.part0[21] );
tran (\sa_count[0][21] , \sa_count[0].f.lower[21] );
tran (\sa_count[0][20] , \sa_count[0].r.part0[20] );
tran (\sa_count[0][20] , \sa_count[0].f.lower[20] );
tran (\sa_count[0][19] , \sa_count[0].r.part0[19] );
tran (\sa_count[0][19] , \sa_count[0].f.lower[19] );
tran (\sa_count[0][18] , \sa_count[0].r.part0[18] );
tran (\sa_count[0][18] , \sa_count[0].f.lower[18] );
tran (\sa_count[0][17] , \sa_count[0].r.part0[17] );
tran (\sa_count[0][17] , \sa_count[0].f.lower[17] );
tran (\sa_count[0][16] , \sa_count[0].r.part0[16] );
tran (\sa_count[0][16] , \sa_count[0].f.lower[16] );
tran (\sa_count[0][15] , \sa_count[0].r.part0[15] );
tran (\sa_count[0][15] , \sa_count[0].f.lower[15] );
tran (\sa_count[0][14] , \sa_count[0].r.part0[14] );
tran (\sa_count[0][14] , \sa_count[0].f.lower[14] );
tran (\sa_count[0][13] , \sa_count[0].r.part0[13] );
tran (\sa_count[0][13] , \sa_count[0].f.lower[13] );
tran (\sa_count[0][12] , \sa_count[0].r.part0[12] );
tran (\sa_count[0][12] , \sa_count[0].f.lower[12] );
tran (\sa_count[0][11] , \sa_count[0].r.part0[11] );
tran (\sa_count[0][11] , \sa_count[0].f.lower[11] );
tran (\sa_count[0][10] , \sa_count[0].r.part0[10] );
tran (\sa_count[0][10] , \sa_count[0].f.lower[10] );
tran (\sa_count[0][9] , \sa_count[0].r.part0[9] );
tran (\sa_count[0][9] , \sa_count[0].f.lower[9] );
tran (\sa_count[0][8] , \sa_count[0].r.part0[8] );
tran (\sa_count[0][8] , \sa_count[0].f.lower[8] );
tran (\sa_count[0][7] , \sa_count[0].r.part0[7] );
tran (\sa_count[0][7] , \sa_count[0].f.lower[7] );
tran (\sa_count[0][6] , \sa_count[0].r.part0[6] );
tran (\sa_count[0][6] , \sa_count[0].f.lower[6] );
tran (\sa_count[0][5] , \sa_count[0].r.part0[5] );
tran (\sa_count[0][5] , \sa_count[0].f.lower[5] );
tran (\sa_count[0][4] , \sa_count[0].r.part0[4] );
tran (\sa_count[0][4] , \sa_count[0].f.lower[4] );
tran (\sa_count[0][3] , \sa_count[0].r.part0[3] );
tran (\sa_count[0][3] , \sa_count[0].f.lower[3] );
tran (\sa_count[0][2] , \sa_count[0].r.part0[2] );
tran (\sa_count[0][2] , \sa_count[0].f.lower[2] );
tran (\sa_count[0][1] , \sa_count[0].r.part0[1] );
tran (\sa_count[0][1] , \sa_count[0].f.lower[1] );
tran (\sa_count[0][0] , \sa_count[0].r.part0[0] );
tran (\sa_count[0][0] , \sa_count[0].f.lower[0] );
tran (\_zy_simnet_tvar_53[7][271] , \_zy_simnet_tvar_53[7].guid_size[0] );
tran (\_zy_simnet_tvar_53[7][270] , \_zy_simnet_tvar_53[7].label_size[5] );
tran (\_zy_simnet_tvar_53[7][269] , \_zy_simnet_tvar_53[7].label_size[4] );
tran (\_zy_simnet_tvar_53[7][268] , \_zy_simnet_tvar_53[7].label_size[3] );
tran (\_zy_simnet_tvar_53[7][267] , \_zy_simnet_tvar_53[7].label_size[2] );
tran (\_zy_simnet_tvar_53[7][266] , \_zy_simnet_tvar_53[7].label_size[1] );
tran (\_zy_simnet_tvar_53[7][265] , \_zy_simnet_tvar_53[7].label_size[0] );
tran (\_zy_simnet_tvar_53[7][264] , \_zy_simnet_tvar_53[7].label[255] );
tran (\_zy_simnet_tvar_53[7][263] , \_zy_simnet_tvar_53[7].label[254] );
tran (\_zy_simnet_tvar_53[7][262] , \_zy_simnet_tvar_53[7].label[253] );
tran (\_zy_simnet_tvar_53[7][261] , \_zy_simnet_tvar_53[7].label[252] );
tran (\_zy_simnet_tvar_53[7][260] , \_zy_simnet_tvar_53[7].label[251] );
tran (\_zy_simnet_tvar_53[7][259] , \_zy_simnet_tvar_53[7].label[250] );
tran (\_zy_simnet_tvar_53[7][258] , \_zy_simnet_tvar_53[7].label[249] );
tran (\_zy_simnet_tvar_53[7][257] , \_zy_simnet_tvar_53[7].label[248] );
tran (\_zy_simnet_tvar_53[7][256] , \_zy_simnet_tvar_53[7].label[247] );
tran (\_zy_simnet_tvar_53[7][255] , \_zy_simnet_tvar_53[7].label[246] );
tran (\_zy_simnet_tvar_53[7][254] , \_zy_simnet_tvar_53[7].label[245] );
tran (\_zy_simnet_tvar_53[7][253] , \_zy_simnet_tvar_53[7].label[244] );
tran (\_zy_simnet_tvar_53[7][252] , \_zy_simnet_tvar_53[7].label[243] );
tran (\_zy_simnet_tvar_53[7][251] , \_zy_simnet_tvar_53[7].label[242] );
tran (\_zy_simnet_tvar_53[7][250] , \_zy_simnet_tvar_53[7].label[241] );
tran (\_zy_simnet_tvar_53[7][249] , \_zy_simnet_tvar_53[7].label[240] );
tran (\_zy_simnet_tvar_53[7][248] , \_zy_simnet_tvar_53[7].label[239] );
tran (\_zy_simnet_tvar_53[7][247] , \_zy_simnet_tvar_53[7].label[238] );
tran (\_zy_simnet_tvar_53[7][246] , \_zy_simnet_tvar_53[7].label[237] );
tran (\_zy_simnet_tvar_53[7][245] , \_zy_simnet_tvar_53[7].label[236] );
tran (\_zy_simnet_tvar_53[7][244] , \_zy_simnet_tvar_53[7].label[235] );
tran (\_zy_simnet_tvar_53[7][243] , \_zy_simnet_tvar_53[7].label[234] );
tran (\_zy_simnet_tvar_53[7][242] , \_zy_simnet_tvar_53[7].label[233] );
tran (\_zy_simnet_tvar_53[7][241] , \_zy_simnet_tvar_53[7].label[232] );
tran (\_zy_simnet_tvar_53[7][240] , \_zy_simnet_tvar_53[7].label[231] );
tran (\_zy_simnet_tvar_53[7][239] , \_zy_simnet_tvar_53[7].label[230] );
tran (\_zy_simnet_tvar_53[7][238] , \_zy_simnet_tvar_53[7].label[229] );
tran (\_zy_simnet_tvar_53[7][237] , \_zy_simnet_tvar_53[7].label[228] );
tran (\_zy_simnet_tvar_53[7][236] , \_zy_simnet_tvar_53[7].label[227] );
tran (\_zy_simnet_tvar_53[7][235] , \_zy_simnet_tvar_53[7].label[226] );
tran (\_zy_simnet_tvar_53[7][234] , \_zy_simnet_tvar_53[7].label[225] );
tran (\_zy_simnet_tvar_53[7][233] , \_zy_simnet_tvar_53[7].label[224] );
tran (\_zy_simnet_tvar_53[7][232] , \_zy_simnet_tvar_53[7].label[223] );
tran (\_zy_simnet_tvar_53[7][231] , \_zy_simnet_tvar_53[7].label[222] );
tran (\_zy_simnet_tvar_53[7][230] , \_zy_simnet_tvar_53[7].label[221] );
tran (\_zy_simnet_tvar_53[7][229] , \_zy_simnet_tvar_53[7].label[220] );
tran (\_zy_simnet_tvar_53[7][228] , \_zy_simnet_tvar_53[7].label[219] );
tran (\_zy_simnet_tvar_53[7][227] , \_zy_simnet_tvar_53[7].label[218] );
tran (\_zy_simnet_tvar_53[7][226] , \_zy_simnet_tvar_53[7].label[217] );
tran (\_zy_simnet_tvar_53[7][225] , \_zy_simnet_tvar_53[7].label[216] );
tran (\_zy_simnet_tvar_53[7][224] , \_zy_simnet_tvar_53[7].label[215] );
tran (\_zy_simnet_tvar_53[7][223] , \_zy_simnet_tvar_53[7].label[214] );
tran (\_zy_simnet_tvar_53[7][222] , \_zy_simnet_tvar_53[7].label[213] );
tran (\_zy_simnet_tvar_53[7][221] , \_zy_simnet_tvar_53[7].label[212] );
tran (\_zy_simnet_tvar_53[7][220] , \_zy_simnet_tvar_53[7].label[211] );
tran (\_zy_simnet_tvar_53[7][219] , \_zy_simnet_tvar_53[7].label[210] );
tran (\_zy_simnet_tvar_53[7][218] , \_zy_simnet_tvar_53[7].label[209] );
tran (\_zy_simnet_tvar_53[7][217] , \_zy_simnet_tvar_53[7].label[208] );
tran (\_zy_simnet_tvar_53[7][216] , \_zy_simnet_tvar_53[7].label[207] );
tran (\_zy_simnet_tvar_53[7][215] , \_zy_simnet_tvar_53[7].label[206] );
tran (\_zy_simnet_tvar_53[7][214] , \_zy_simnet_tvar_53[7].label[205] );
tran (\_zy_simnet_tvar_53[7][213] , \_zy_simnet_tvar_53[7].label[204] );
tran (\_zy_simnet_tvar_53[7][212] , \_zy_simnet_tvar_53[7].label[203] );
tran (\_zy_simnet_tvar_53[7][211] , \_zy_simnet_tvar_53[7].label[202] );
tran (\_zy_simnet_tvar_53[7][210] , \_zy_simnet_tvar_53[7].label[201] );
tran (\_zy_simnet_tvar_53[7][209] , \_zy_simnet_tvar_53[7].label[200] );
tran (\_zy_simnet_tvar_53[7][208] , \_zy_simnet_tvar_53[7].label[199] );
tran (\_zy_simnet_tvar_53[7][207] , \_zy_simnet_tvar_53[7].label[198] );
tran (\_zy_simnet_tvar_53[7][206] , \_zy_simnet_tvar_53[7].label[197] );
tran (\_zy_simnet_tvar_53[7][205] , \_zy_simnet_tvar_53[7].label[196] );
tran (\_zy_simnet_tvar_53[7][204] , \_zy_simnet_tvar_53[7].label[195] );
tran (\_zy_simnet_tvar_53[7][203] , \_zy_simnet_tvar_53[7].label[194] );
tran (\_zy_simnet_tvar_53[7][202] , \_zy_simnet_tvar_53[7].label[193] );
tran (\_zy_simnet_tvar_53[7][201] , \_zy_simnet_tvar_53[7].label[192] );
tran (\_zy_simnet_tvar_53[7][200] , \_zy_simnet_tvar_53[7].label[191] );
tran (\_zy_simnet_tvar_53[7][199] , \_zy_simnet_tvar_53[7].label[190] );
tran (\_zy_simnet_tvar_53[7][198] , \_zy_simnet_tvar_53[7].label[189] );
tran (\_zy_simnet_tvar_53[7][197] , \_zy_simnet_tvar_53[7].label[188] );
tran (\_zy_simnet_tvar_53[7][196] , \_zy_simnet_tvar_53[7].label[187] );
tran (\_zy_simnet_tvar_53[7][195] , \_zy_simnet_tvar_53[7].label[186] );
tran (\_zy_simnet_tvar_53[7][194] , \_zy_simnet_tvar_53[7].label[185] );
tran (\_zy_simnet_tvar_53[7][193] , \_zy_simnet_tvar_53[7].label[184] );
tran (\_zy_simnet_tvar_53[7][192] , \_zy_simnet_tvar_53[7].label[183] );
tran (\_zy_simnet_tvar_53[7][191] , \_zy_simnet_tvar_53[7].label[182] );
tran (\_zy_simnet_tvar_53[7][190] , \_zy_simnet_tvar_53[7].label[181] );
tran (\_zy_simnet_tvar_53[7][189] , \_zy_simnet_tvar_53[7].label[180] );
tran (\_zy_simnet_tvar_53[7][188] , \_zy_simnet_tvar_53[7].label[179] );
tran (\_zy_simnet_tvar_53[7][187] , \_zy_simnet_tvar_53[7].label[178] );
tran (\_zy_simnet_tvar_53[7][186] , \_zy_simnet_tvar_53[7].label[177] );
tran (\_zy_simnet_tvar_53[7][185] , \_zy_simnet_tvar_53[7].label[176] );
tran (\_zy_simnet_tvar_53[7][184] , \_zy_simnet_tvar_53[7].label[175] );
tran (\_zy_simnet_tvar_53[7][183] , \_zy_simnet_tvar_53[7].label[174] );
tran (\_zy_simnet_tvar_53[7][182] , \_zy_simnet_tvar_53[7].label[173] );
tran (\_zy_simnet_tvar_53[7][181] , \_zy_simnet_tvar_53[7].label[172] );
tran (\_zy_simnet_tvar_53[7][180] , \_zy_simnet_tvar_53[7].label[171] );
tran (\_zy_simnet_tvar_53[7][179] , \_zy_simnet_tvar_53[7].label[170] );
tran (\_zy_simnet_tvar_53[7][178] , \_zy_simnet_tvar_53[7].label[169] );
tran (\_zy_simnet_tvar_53[7][177] , \_zy_simnet_tvar_53[7].label[168] );
tran (\_zy_simnet_tvar_53[7][176] , \_zy_simnet_tvar_53[7].label[167] );
tran (\_zy_simnet_tvar_53[7][175] , \_zy_simnet_tvar_53[7].label[166] );
tran (\_zy_simnet_tvar_53[7][174] , \_zy_simnet_tvar_53[7].label[165] );
tran (\_zy_simnet_tvar_53[7][173] , \_zy_simnet_tvar_53[7].label[164] );
tran (\_zy_simnet_tvar_53[7][172] , \_zy_simnet_tvar_53[7].label[163] );
tran (\_zy_simnet_tvar_53[7][171] , \_zy_simnet_tvar_53[7].label[162] );
tran (\_zy_simnet_tvar_53[7][170] , \_zy_simnet_tvar_53[7].label[161] );
tran (\_zy_simnet_tvar_53[7][169] , \_zy_simnet_tvar_53[7].label[160] );
tran (\_zy_simnet_tvar_53[7][168] , \_zy_simnet_tvar_53[7].label[159] );
tran (\_zy_simnet_tvar_53[7][167] , \_zy_simnet_tvar_53[7].label[158] );
tran (\_zy_simnet_tvar_53[7][166] , \_zy_simnet_tvar_53[7].label[157] );
tran (\_zy_simnet_tvar_53[7][165] , \_zy_simnet_tvar_53[7].label[156] );
tran (\_zy_simnet_tvar_53[7][164] , \_zy_simnet_tvar_53[7].label[155] );
tran (\_zy_simnet_tvar_53[7][163] , \_zy_simnet_tvar_53[7].label[154] );
tran (\_zy_simnet_tvar_53[7][162] , \_zy_simnet_tvar_53[7].label[153] );
tran (\_zy_simnet_tvar_53[7][161] , \_zy_simnet_tvar_53[7].label[152] );
tran (\_zy_simnet_tvar_53[7][160] , \_zy_simnet_tvar_53[7].label[151] );
tran (\_zy_simnet_tvar_53[7][159] , \_zy_simnet_tvar_53[7].label[150] );
tran (\_zy_simnet_tvar_53[7][158] , \_zy_simnet_tvar_53[7].label[149] );
tran (\_zy_simnet_tvar_53[7][157] , \_zy_simnet_tvar_53[7].label[148] );
tran (\_zy_simnet_tvar_53[7][156] , \_zy_simnet_tvar_53[7].label[147] );
tran (\_zy_simnet_tvar_53[7][155] , \_zy_simnet_tvar_53[7].label[146] );
tran (\_zy_simnet_tvar_53[7][154] , \_zy_simnet_tvar_53[7].label[145] );
tran (\_zy_simnet_tvar_53[7][153] , \_zy_simnet_tvar_53[7].label[144] );
tran (\_zy_simnet_tvar_53[7][152] , \_zy_simnet_tvar_53[7].label[143] );
tran (\_zy_simnet_tvar_53[7][151] , \_zy_simnet_tvar_53[7].label[142] );
tran (\_zy_simnet_tvar_53[7][150] , \_zy_simnet_tvar_53[7].label[141] );
tran (\_zy_simnet_tvar_53[7][149] , \_zy_simnet_tvar_53[7].label[140] );
tran (\_zy_simnet_tvar_53[7][148] , \_zy_simnet_tvar_53[7].label[139] );
tran (\_zy_simnet_tvar_53[7][147] , \_zy_simnet_tvar_53[7].label[138] );
tran (\_zy_simnet_tvar_53[7][146] , \_zy_simnet_tvar_53[7].label[137] );
tran (\_zy_simnet_tvar_53[7][145] , \_zy_simnet_tvar_53[7].label[136] );
tran (\_zy_simnet_tvar_53[7][144] , \_zy_simnet_tvar_53[7].label[135] );
tran (\_zy_simnet_tvar_53[7][143] , \_zy_simnet_tvar_53[7].label[134] );
tran (\_zy_simnet_tvar_53[7][142] , \_zy_simnet_tvar_53[7].label[133] );
tran (\_zy_simnet_tvar_53[7][141] , \_zy_simnet_tvar_53[7].label[132] );
tran (\_zy_simnet_tvar_53[7][140] , \_zy_simnet_tvar_53[7].label[131] );
tran (\_zy_simnet_tvar_53[7][139] , \_zy_simnet_tvar_53[7].label[130] );
tran (\_zy_simnet_tvar_53[7][138] , \_zy_simnet_tvar_53[7].label[129] );
tran (\_zy_simnet_tvar_53[7][137] , \_zy_simnet_tvar_53[7].label[128] );
tran (\_zy_simnet_tvar_53[7][136] , \_zy_simnet_tvar_53[7].label[127] );
tran (\_zy_simnet_tvar_53[7][135] , \_zy_simnet_tvar_53[7].label[126] );
tran (\_zy_simnet_tvar_53[7][134] , \_zy_simnet_tvar_53[7].label[125] );
tran (\_zy_simnet_tvar_53[7][133] , \_zy_simnet_tvar_53[7].label[124] );
tran (\_zy_simnet_tvar_53[7][132] , \_zy_simnet_tvar_53[7].label[123] );
tran (\_zy_simnet_tvar_53[7][131] , \_zy_simnet_tvar_53[7].label[122] );
tran (\_zy_simnet_tvar_53[7][130] , \_zy_simnet_tvar_53[7].label[121] );
tran (\_zy_simnet_tvar_53[7][129] , \_zy_simnet_tvar_53[7].label[120] );
tran (\_zy_simnet_tvar_53[7][128] , \_zy_simnet_tvar_53[7].label[119] );
tran (\_zy_simnet_tvar_53[7][127] , \_zy_simnet_tvar_53[7].label[118] );
tran (\_zy_simnet_tvar_53[7][126] , \_zy_simnet_tvar_53[7].label[117] );
tran (\_zy_simnet_tvar_53[7][125] , \_zy_simnet_tvar_53[7].label[116] );
tran (\_zy_simnet_tvar_53[7][124] , \_zy_simnet_tvar_53[7].label[115] );
tran (\_zy_simnet_tvar_53[7][123] , \_zy_simnet_tvar_53[7].label[114] );
tran (\_zy_simnet_tvar_53[7][122] , \_zy_simnet_tvar_53[7].label[113] );
tran (\_zy_simnet_tvar_53[7][121] , \_zy_simnet_tvar_53[7].label[112] );
tran (\_zy_simnet_tvar_53[7][120] , \_zy_simnet_tvar_53[7].label[111] );
tran (\_zy_simnet_tvar_53[7][119] , \_zy_simnet_tvar_53[7].label[110] );
tran (\_zy_simnet_tvar_53[7][118] , \_zy_simnet_tvar_53[7].label[109] );
tran (\_zy_simnet_tvar_53[7][117] , \_zy_simnet_tvar_53[7].label[108] );
tran (\_zy_simnet_tvar_53[7][116] , \_zy_simnet_tvar_53[7].label[107] );
tran (\_zy_simnet_tvar_53[7][115] , \_zy_simnet_tvar_53[7].label[106] );
tran (\_zy_simnet_tvar_53[7][114] , \_zy_simnet_tvar_53[7].label[105] );
tran (\_zy_simnet_tvar_53[7][113] , \_zy_simnet_tvar_53[7].label[104] );
tran (\_zy_simnet_tvar_53[7][112] , \_zy_simnet_tvar_53[7].label[103] );
tran (\_zy_simnet_tvar_53[7][111] , \_zy_simnet_tvar_53[7].label[102] );
tran (\_zy_simnet_tvar_53[7][110] , \_zy_simnet_tvar_53[7].label[101] );
tran (\_zy_simnet_tvar_53[7][109] , \_zy_simnet_tvar_53[7].label[100] );
tran (\_zy_simnet_tvar_53[7][108] , \_zy_simnet_tvar_53[7].label[99] );
tran (\_zy_simnet_tvar_53[7][107] , \_zy_simnet_tvar_53[7].label[98] );
tran (\_zy_simnet_tvar_53[7][106] , \_zy_simnet_tvar_53[7].label[97] );
tran (\_zy_simnet_tvar_53[7][105] , \_zy_simnet_tvar_53[7].label[96] );
tran (\_zy_simnet_tvar_53[7][104] , \_zy_simnet_tvar_53[7].label[95] );
tran (\_zy_simnet_tvar_53[7][103] , \_zy_simnet_tvar_53[7].label[94] );
tran (\_zy_simnet_tvar_53[7][102] , \_zy_simnet_tvar_53[7].label[93] );
tran (\_zy_simnet_tvar_53[7][101] , \_zy_simnet_tvar_53[7].label[92] );
tran (\_zy_simnet_tvar_53[7][100] , \_zy_simnet_tvar_53[7].label[91] );
tran (\_zy_simnet_tvar_53[7][99] , \_zy_simnet_tvar_53[7].label[90] );
tran (\_zy_simnet_tvar_53[7][98] , \_zy_simnet_tvar_53[7].label[89] );
tran (\_zy_simnet_tvar_53[7][97] , \_zy_simnet_tvar_53[7].label[88] );
tran (\_zy_simnet_tvar_53[7][96] , \_zy_simnet_tvar_53[7].label[87] );
tran (\_zy_simnet_tvar_53[7][95] , \_zy_simnet_tvar_53[7].label[86] );
tran (\_zy_simnet_tvar_53[7][94] , \_zy_simnet_tvar_53[7].label[85] );
tran (\_zy_simnet_tvar_53[7][93] , \_zy_simnet_tvar_53[7].label[84] );
tran (\_zy_simnet_tvar_53[7][92] , \_zy_simnet_tvar_53[7].label[83] );
tran (\_zy_simnet_tvar_53[7][91] , \_zy_simnet_tvar_53[7].label[82] );
tran (\_zy_simnet_tvar_53[7][90] , \_zy_simnet_tvar_53[7].label[81] );
tran (\_zy_simnet_tvar_53[7][89] , \_zy_simnet_tvar_53[7].label[80] );
tran (\_zy_simnet_tvar_53[7][88] , \_zy_simnet_tvar_53[7].label[79] );
tran (\_zy_simnet_tvar_53[7][87] , \_zy_simnet_tvar_53[7].label[78] );
tran (\_zy_simnet_tvar_53[7][86] , \_zy_simnet_tvar_53[7].label[77] );
tran (\_zy_simnet_tvar_53[7][85] , \_zy_simnet_tvar_53[7].label[76] );
tran (\_zy_simnet_tvar_53[7][84] , \_zy_simnet_tvar_53[7].label[75] );
tran (\_zy_simnet_tvar_53[7][83] , \_zy_simnet_tvar_53[7].label[74] );
tran (\_zy_simnet_tvar_53[7][82] , \_zy_simnet_tvar_53[7].label[73] );
tran (\_zy_simnet_tvar_53[7][81] , \_zy_simnet_tvar_53[7].label[72] );
tran (\_zy_simnet_tvar_53[7][80] , \_zy_simnet_tvar_53[7].label[71] );
tran (\_zy_simnet_tvar_53[7][79] , \_zy_simnet_tvar_53[7].label[70] );
tran (\_zy_simnet_tvar_53[7][78] , \_zy_simnet_tvar_53[7].label[69] );
tran (\_zy_simnet_tvar_53[7][77] , \_zy_simnet_tvar_53[7].label[68] );
tran (\_zy_simnet_tvar_53[7][76] , \_zy_simnet_tvar_53[7].label[67] );
tran (\_zy_simnet_tvar_53[7][75] , \_zy_simnet_tvar_53[7].label[66] );
tran (\_zy_simnet_tvar_53[7][74] , \_zy_simnet_tvar_53[7].label[65] );
tran (\_zy_simnet_tvar_53[7][73] , \_zy_simnet_tvar_53[7].label[64] );
tran (\_zy_simnet_tvar_53[7][72] , \_zy_simnet_tvar_53[7].label[63] );
tran (\_zy_simnet_tvar_53[7][71] , \_zy_simnet_tvar_53[7].label[62] );
tran (\_zy_simnet_tvar_53[7][70] , \_zy_simnet_tvar_53[7].label[61] );
tran (\_zy_simnet_tvar_53[7][69] , \_zy_simnet_tvar_53[7].label[60] );
tran (\_zy_simnet_tvar_53[7][68] , \_zy_simnet_tvar_53[7].label[59] );
tran (\_zy_simnet_tvar_53[7][67] , \_zy_simnet_tvar_53[7].label[58] );
tran (\_zy_simnet_tvar_53[7][66] , \_zy_simnet_tvar_53[7].label[57] );
tran (\_zy_simnet_tvar_53[7][65] , \_zy_simnet_tvar_53[7].label[56] );
tran (\_zy_simnet_tvar_53[7][64] , \_zy_simnet_tvar_53[7].label[55] );
tran (\_zy_simnet_tvar_53[7][63] , \_zy_simnet_tvar_53[7].label[54] );
tran (\_zy_simnet_tvar_53[7][62] , \_zy_simnet_tvar_53[7].label[53] );
tran (\_zy_simnet_tvar_53[7][61] , \_zy_simnet_tvar_53[7].label[52] );
tran (\_zy_simnet_tvar_53[7][60] , \_zy_simnet_tvar_53[7].label[51] );
tran (\_zy_simnet_tvar_53[7][59] , \_zy_simnet_tvar_53[7].label[50] );
tran (\_zy_simnet_tvar_53[7][58] , \_zy_simnet_tvar_53[7].label[49] );
tran (\_zy_simnet_tvar_53[7][57] , \_zy_simnet_tvar_53[7].label[48] );
tran (\_zy_simnet_tvar_53[7][56] , \_zy_simnet_tvar_53[7].label[47] );
tran (\_zy_simnet_tvar_53[7][55] , \_zy_simnet_tvar_53[7].label[46] );
tran (\_zy_simnet_tvar_53[7][54] , \_zy_simnet_tvar_53[7].label[45] );
tran (\_zy_simnet_tvar_53[7][53] , \_zy_simnet_tvar_53[7].label[44] );
tran (\_zy_simnet_tvar_53[7][52] , \_zy_simnet_tvar_53[7].label[43] );
tran (\_zy_simnet_tvar_53[7][51] , \_zy_simnet_tvar_53[7].label[42] );
tran (\_zy_simnet_tvar_53[7][50] , \_zy_simnet_tvar_53[7].label[41] );
tran (\_zy_simnet_tvar_53[7][49] , \_zy_simnet_tvar_53[7].label[40] );
tran (\_zy_simnet_tvar_53[7][48] , \_zy_simnet_tvar_53[7].label[39] );
tran (\_zy_simnet_tvar_53[7][47] , \_zy_simnet_tvar_53[7].label[38] );
tran (\_zy_simnet_tvar_53[7][46] , \_zy_simnet_tvar_53[7].label[37] );
tran (\_zy_simnet_tvar_53[7][45] , \_zy_simnet_tvar_53[7].label[36] );
tran (\_zy_simnet_tvar_53[7][44] , \_zy_simnet_tvar_53[7].label[35] );
tran (\_zy_simnet_tvar_53[7][43] , \_zy_simnet_tvar_53[7].label[34] );
tran (\_zy_simnet_tvar_53[7][42] , \_zy_simnet_tvar_53[7].label[33] );
tran (\_zy_simnet_tvar_53[7][41] , \_zy_simnet_tvar_53[7].label[32] );
tran (\_zy_simnet_tvar_53[7][40] , \_zy_simnet_tvar_53[7].label[31] );
tran (\_zy_simnet_tvar_53[7][39] , \_zy_simnet_tvar_53[7].label[30] );
tran (\_zy_simnet_tvar_53[7][38] , \_zy_simnet_tvar_53[7].label[29] );
tran (\_zy_simnet_tvar_53[7][37] , \_zy_simnet_tvar_53[7].label[28] );
tran (\_zy_simnet_tvar_53[7][36] , \_zy_simnet_tvar_53[7].label[27] );
tran (\_zy_simnet_tvar_53[7][35] , \_zy_simnet_tvar_53[7].label[26] );
tran (\_zy_simnet_tvar_53[7][34] , \_zy_simnet_tvar_53[7].label[25] );
tran (\_zy_simnet_tvar_53[7][33] , \_zy_simnet_tvar_53[7].label[24] );
tran (\_zy_simnet_tvar_53[7][32] , \_zy_simnet_tvar_53[7].label[23] );
tran (\_zy_simnet_tvar_53[7][31] , \_zy_simnet_tvar_53[7].label[22] );
tran (\_zy_simnet_tvar_53[7][30] , \_zy_simnet_tvar_53[7].label[21] );
tran (\_zy_simnet_tvar_53[7][29] , \_zy_simnet_tvar_53[7].label[20] );
tran (\_zy_simnet_tvar_53[7][28] , \_zy_simnet_tvar_53[7].label[19] );
tran (\_zy_simnet_tvar_53[7][27] , \_zy_simnet_tvar_53[7].label[18] );
tran (\_zy_simnet_tvar_53[7][26] , \_zy_simnet_tvar_53[7].label[17] );
tran (\_zy_simnet_tvar_53[7][25] , \_zy_simnet_tvar_53[7].label[16] );
tran (\_zy_simnet_tvar_53[7][24] , \_zy_simnet_tvar_53[7].label[15] );
tran (\_zy_simnet_tvar_53[7][23] , \_zy_simnet_tvar_53[7].label[14] );
tran (\_zy_simnet_tvar_53[7][22] , \_zy_simnet_tvar_53[7].label[13] );
tran (\_zy_simnet_tvar_53[7][21] , \_zy_simnet_tvar_53[7].label[12] );
tran (\_zy_simnet_tvar_53[7][20] , \_zy_simnet_tvar_53[7].label[11] );
tran (\_zy_simnet_tvar_53[7][19] , \_zy_simnet_tvar_53[7].label[10] );
tran (\_zy_simnet_tvar_53[7][18] , \_zy_simnet_tvar_53[7].label[9] );
tran (\_zy_simnet_tvar_53[7][17] , \_zy_simnet_tvar_53[7].label[8] );
tran (\_zy_simnet_tvar_53[7][16] , \_zy_simnet_tvar_53[7].label[7] );
tran (\_zy_simnet_tvar_53[7][15] , \_zy_simnet_tvar_53[7].label[6] );
tran (\_zy_simnet_tvar_53[7][14] , \_zy_simnet_tvar_53[7].label[5] );
tran (\_zy_simnet_tvar_53[7][13] , \_zy_simnet_tvar_53[7].label[4] );
tran (\_zy_simnet_tvar_53[7][12] , \_zy_simnet_tvar_53[7].label[3] );
tran (\_zy_simnet_tvar_53[7][11] , \_zy_simnet_tvar_53[7].label[2] );
tran (\_zy_simnet_tvar_53[7][10] , \_zy_simnet_tvar_53[7].label[1] );
tran (\_zy_simnet_tvar_53[7][9] , \_zy_simnet_tvar_53[7].label[0] );
tran (\_zy_simnet_tvar_53[7][8] , \_zy_simnet_tvar_53[7].delimiter_valid[0] );
tran (\_zy_simnet_tvar_53[7][7] , \_zy_simnet_tvar_53[7].delimiter[7] );
tran (\_zy_simnet_tvar_53[7][6] , \_zy_simnet_tvar_53[7].delimiter[6] );
tran (\_zy_simnet_tvar_53[7][5] , \_zy_simnet_tvar_53[7].delimiter[5] );
tran (\_zy_simnet_tvar_53[7][4] , \_zy_simnet_tvar_53[7].delimiter[4] );
tran (\_zy_simnet_tvar_53[7][3] , \_zy_simnet_tvar_53[7].delimiter[3] );
tran (\_zy_simnet_tvar_53[7][2] , \_zy_simnet_tvar_53[7].delimiter[2] );
tran (\_zy_simnet_tvar_53[7][1] , \_zy_simnet_tvar_53[7].delimiter[1] );
tran (\_zy_simnet_tvar_53[7][0] , \_zy_simnet_tvar_53[7].delimiter[0] );
tran (\_zy_simnet_tvar_53[6][271] , \_zy_simnet_tvar_53[6].guid_size[0] );
tran (\_zy_simnet_tvar_53[6][270] , \_zy_simnet_tvar_53[6].label_size[5] );
tran (\_zy_simnet_tvar_53[6][269] , \_zy_simnet_tvar_53[6].label_size[4] );
tran (\_zy_simnet_tvar_53[6][268] , \_zy_simnet_tvar_53[6].label_size[3] );
tran (\_zy_simnet_tvar_53[6][267] , \_zy_simnet_tvar_53[6].label_size[2] );
tran (\_zy_simnet_tvar_53[6][266] , \_zy_simnet_tvar_53[6].label_size[1] );
tran (\_zy_simnet_tvar_53[6][265] , \_zy_simnet_tvar_53[6].label_size[0] );
tran (\_zy_simnet_tvar_53[6][264] , \_zy_simnet_tvar_53[6].label[255] );
tran (\_zy_simnet_tvar_53[6][263] , \_zy_simnet_tvar_53[6].label[254] );
tran (\_zy_simnet_tvar_53[6][262] , \_zy_simnet_tvar_53[6].label[253] );
tran (\_zy_simnet_tvar_53[6][261] , \_zy_simnet_tvar_53[6].label[252] );
tran (\_zy_simnet_tvar_53[6][260] , \_zy_simnet_tvar_53[6].label[251] );
tran (\_zy_simnet_tvar_53[6][259] , \_zy_simnet_tvar_53[6].label[250] );
tran (\_zy_simnet_tvar_53[6][258] , \_zy_simnet_tvar_53[6].label[249] );
tran (\_zy_simnet_tvar_53[6][257] , \_zy_simnet_tvar_53[6].label[248] );
tran (\_zy_simnet_tvar_53[6][256] , \_zy_simnet_tvar_53[6].label[247] );
tran (\_zy_simnet_tvar_53[6][255] , \_zy_simnet_tvar_53[6].label[246] );
tran (\_zy_simnet_tvar_53[6][254] , \_zy_simnet_tvar_53[6].label[245] );
tran (\_zy_simnet_tvar_53[6][253] , \_zy_simnet_tvar_53[6].label[244] );
tran (\_zy_simnet_tvar_53[6][252] , \_zy_simnet_tvar_53[6].label[243] );
tran (\_zy_simnet_tvar_53[6][251] , \_zy_simnet_tvar_53[6].label[242] );
tran (\_zy_simnet_tvar_53[6][250] , \_zy_simnet_tvar_53[6].label[241] );
tran (\_zy_simnet_tvar_53[6][249] , \_zy_simnet_tvar_53[6].label[240] );
tran (\_zy_simnet_tvar_53[6][248] , \_zy_simnet_tvar_53[6].label[239] );
tran (\_zy_simnet_tvar_53[6][247] , \_zy_simnet_tvar_53[6].label[238] );
tran (\_zy_simnet_tvar_53[6][246] , \_zy_simnet_tvar_53[6].label[237] );
tran (\_zy_simnet_tvar_53[6][245] , \_zy_simnet_tvar_53[6].label[236] );
tran (\_zy_simnet_tvar_53[6][244] , \_zy_simnet_tvar_53[6].label[235] );
tran (\_zy_simnet_tvar_53[6][243] , \_zy_simnet_tvar_53[6].label[234] );
tran (\_zy_simnet_tvar_53[6][242] , \_zy_simnet_tvar_53[6].label[233] );
tran (\_zy_simnet_tvar_53[6][241] , \_zy_simnet_tvar_53[6].label[232] );
tran (\_zy_simnet_tvar_53[6][240] , \_zy_simnet_tvar_53[6].label[231] );
tran (\_zy_simnet_tvar_53[6][239] , \_zy_simnet_tvar_53[6].label[230] );
tran (\_zy_simnet_tvar_53[6][238] , \_zy_simnet_tvar_53[6].label[229] );
tran (\_zy_simnet_tvar_53[6][237] , \_zy_simnet_tvar_53[6].label[228] );
tran (\_zy_simnet_tvar_53[6][236] , \_zy_simnet_tvar_53[6].label[227] );
tran (\_zy_simnet_tvar_53[6][235] , \_zy_simnet_tvar_53[6].label[226] );
tran (\_zy_simnet_tvar_53[6][234] , \_zy_simnet_tvar_53[6].label[225] );
tran (\_zy_simnet_tvar_53[6][233] , \_zy_simnet_tvar_53[6].label[224] );
tran (\_zy_simnet_tvar_53[6][232] , \_zy_simnet_tvar_53[6].label[223] );
tran (\_zy_simnet_tvar_53[6][231] , \_zy_simnet_tvar_53[6].label[222] );
tran (\_zy_simnet_tvar_53[6][230] , \_zy_simnet_tvar_53[6].label[221] );
tran (\_zy_simnet_tvar_53[6][229] , \_zy_simnet_tvar_53[6].label[220] );
tran (\_zy_simnet_tvar_53[6][228] , \_zy_simnet_tvar_53[6].label[219] );
tran (\_zy_simnet_tvar_53[6][227] , \_zy_simnet_tvar_53[6].label[218] );
tran (\_zy_simnet_tvar_53[6][226] , \_zy_simnet_tvar_53[6].label[217] );
tran (\_zy_simnet_tvar_53[6][225] , \_zy_simnet_tvar_53[6].label[216] );
tran (\_zy_simnet_tvar_53[6][224] , \_zy_simnet_tvar_53[6].label[215] );
tran (\_zy_simnet_tvar_53[6][223] , \_zy_simnet_tvar_53[6].label[214] );
tran (\_zy_simnet_tvar_53[6][222] , \_zy_simnet_tvar_53[6].label[213] );
tran (\_zy_simnet_tvar_53[6][221] , \_zy_simnet_tvar_53[6].label[212] );
tran (\_zy_simnet_tvar_53[6][220] , \_zy_simnet_tvar_53[6].label[211] );
tran (\_zy_simnet_tvar_53[6][219] , \_zy_simnet_tvar_53[6].label[210] );
tran (\_zy_simnet_tvar_53[6][218] , \_zy_simnet_tvar_53[6].label[209] );
tran (\_zy_simnet_tvar_53[6][217] , \_zy_simnet_tvar_53[6].label[208] );
tran (\_zy_simnet_tvar_53[6][216] , \_zy_simnet_tvar_53[6].label[207] );
tran (\_zy_simnet_tvar_53[6][215] , \_zy_simnet_tvar_53[6].label[206] );
tran (\_zy_simnet_tvar_53[6][214] , \_zy_simnet_tvar_53[6].label[205] );
tran (\_zy_simnet_tvar_53[6][213] , \_zy_simnet_tvar_53[6].label[204] );
tran (\_zy_simnet_tvar_53[6][212] , \_zy_simnet_tvar_53[6].label[203] );
tran (\_zy_simnet_tvar_53[6][211] , \_zy_simnet_tvar_53[6].label[202] );
tran (\_zy_simnet_tvar_53[6][210] , \_zy_simnet_tvar_53[6].label[201] );
tran (\_zy_simnet_tvar_53[6][209] , \_zy_simnet_tvar_53[6].label[200] );
tran (\_zy_simnet_tvar_53[6][208] , \_zy_simnet_tvar_53[6].label[199] );
tran (\_zy_simnet_tvar_53[6][207] , \_zy_simnet_tvar_53[6].label[198] );
tran (\_zy_simnet_tvar_53[6][206] , \_zy_simnet_tvar_53[6].label[197] );
tran (\_zy_simnet_tvar_53[6][205] , \_zy_simnet_tvar_53[6].label[196] );
tran (\_zy_simnet_tvar_53[6][204] , \_zy_simnet_tvar_53[6].label[195] );
tran (\_zy_simnet_tvar_53[6][203] , \_zy_simnet_tvar_53[6].label[194] );
tran (\_zy_simnet_tvar_53[6][202] , \_zy_simnet_tvar_53[6].label[193] );
tran (\_zy_simnet_tvar_53[6][201] , \_zy_simnet_tvar_53[6].label[192] );
tran (\_zy_simnet_tvar_53[6][200] , \_zy_simnet_tvar_53[6].label[191] );
tran (\_zy_simnet_tvar_53[6][199] , \_zy_simnet_tvar_53[6].label[190] );
tran (\_zy_simnet_tvar_53[6][198] , \_zy_simnet_tvar_53[6].label[189] );
tran (\_zy_simnet_tvar_53[6][197] , \_zy_simnet_tvar_53[6].label[188] );
tran (\_zy_simnet_tvar_53[6][196] , \_zy_simnet_tvar_53[6].label[187] );
tran (\_zy_simnet_tvar_53[6][195] , \_zy_simnet_tvar_53[6].label[186] );
tran (\_zy_simnet_tvar_53[6][194] , \_zy_simnet_tvar_53[6].label[185] );
tran (\_zy_simnet_tvar_53[6][193] , \_zy_simnet_tvar_53[6].label[184] );
tran (\_zy_simnet_tvar_53[6][192] , \_zy_simnet_tvar_53[6].label[183] );
tran (\_zy_simnet_tvar_53[6][191] , \_zy_simnet_tvar_53[6].label[182] );
tran (\_zy_simnet_tvar_53[6][190] , \_zy_simnet_tvar_53[6].label[181] );
tran (\_zy_simnet_tvar_53[6][189] , \_zy_simnet_tvar_53[6].label[180] );
tran (\_zy_simnet_tvar_53[6][188] , \_zy_simnet_tvar_53[6].label[179] );
tran (\_zy_simnet_tvar_53[6][187] , \_zy_simnet_tvar_53[6].label[178] );
tran (\_zy_simnet_tvar_53[6][186] , \_zy_simnet_tvar_53[6].label[177] );
tran (\_zy_simnet_tvar_53[6][185] , \_zy_simnet_tvar_53[6].label[176] );
tran (\_zy_simnet_tvar_53[6][184] , \_zy_simnet_tvar_53[6].label[175] );
tran (\_zy_simnet_tvar_53[6][183] , \_zy_simnet_tvar_53[6].label[174] );
tran (\_zy_simnet_tvar_53[6][182] , \_zy_simnet_tvar_53[6].label[173] );
tran (\_zy_simnet_tvar_53[6][181] , \_zy_simnet_tvar_53[6].label[172] );
tran (\_zy_simnet_tvar_53[6][180] , \_zy_simnet_tvar_53[6].label[171] );
tran (\_zy_simnet_tvar_53[6][179] , \_zy_simnet_tvar_53[6].label[170] );
tran (\_zy_simnet_tvar_53[6][178] , \_zy_simnet_tvar_53[6].label[169] );
tran (\_zy_simnet_tvar_53[6][177] , \_zy_simnet_tvar_53[6].label[168] );
tran (\_zy_simnet_tvar_53[6][176] , \_zy_simnet_tvar_53[6].label[167] );
tran (\_zy_simnet_tvar_53[6][175] , \_zy_simnet_tvar_53[6].label[166] );
tran (\_zy_simnet_tvar_53[6][174] , \_zy_simnet_tvar_53[6].label[165] );
tran (\_zy_simnet_tvar_53[6][173] , \_zy_simnet_tvar_53[6].label[164] );
tran (\_zy_simnet_tvar_53[6][172] , \_zy_simnet_tvar_53[6].label[163] );
tran (\_zy_simnet_tvar_53[6][171] , \_zy_simnet_tvar_53[6].label[162] );
tran (\_zy_simnet_tvar_53[6][170] , \_zy_simnet_tvar_53[6].label[161] );
tran (\_zy_simnet_tvar_53[6][169] , \_zy_simnet_tvar_53[6].label[160] );
tran (\_zy_simnet_tvar_53[6][168] , \_zy_simnet_tvar_53[6].label[159] );
tran (\_zy_simnet_tvar_53[6][167] , \_zy_simnet_tvar_53[6].label[158] );
tran (\_zy_simnet_tvar_53[6][166] , \_zy_simnet_tvar_53[6].label[157] );
tran (\_zy_simnet_tvar_53[6][165] , \_zy_simnet_tvar_53[6].label[156] );
tran (\_zy_simnet_tvar_53[6][164] , \_zy_simnet_tvar_53[6].label[155] );
tran (\_zy_simnet_tvar_53[6][163] , \_zy_simnet_tvar_53[6].label[154] );
tran (\_zy_simnet_tvar_53[6][162] , \_zy_simnet_tvar_53[6].label[153] );
tran (\_zy_simnet_tvar_53[6][161] , \_zy_simnet_tvar_53[6].label[152] );
tran (\_zy_simnet_tvar_53[6][160] , \_zy_simnet_tvar_53[6].label[151] );
tran (\_zy_simnet_tvar_53[6][159] , \_zy_simnet_tvar_53[6].label[150] );
tran (\_zy_simnet_tvar_53[6][158] , \_zy_simnet_tvar_53[6].label[149] );
tran (\_zy_simnet_tvar_53[6][157] , \_zy_simnet_tvar_53[6].label[148] );
tran (\_zy_simnet_tvar_53[6][156] , \_zy_simnet_tvar_53[6].label[147] );
tran (\_zy_simnet_tvar_53[6][155] , \_zy_simnet_tvar_53[6].label[146] );
tran (\_zy_simnet_tvar_53[6][154] , \_zy_simnet_tvar_53[6].label[145] );
tran (\_zy_simnet_tvar_53[6][153] , \_zy_simnet_tvar_53[6].label[144] );
tran (\_zy_simnet_tvar_53[6][152] , \_zy_simnet_tvar_53[6].label[143] );
tran (\_zy_simnet_tvar_53[6][151] , \_zy_simnet_tvar_53[6].label[142] );
tran (\_zy_simnet_tvar_53[6][150] , \_zy_simnet_tvar_53[6].label[141] );
tran (\_zy_simnet_tvar_53[6][149] , \_zy_simnet_tvar_53[6].label[140] );
tran (\_zy_simnet_tvar_53[6][148] , \_zy_simnet_tvar_53[6].label[139] );
tran (\_zy_simnet_tvar_53[6][147] , \_zy_simnet_tvar_53[6].label[138] );
tran (\_zy_simnet_tvar_53[6][146] , \_zy_simnet_tvar_53[6].label[137] );
tran (\_zy_simnet_tvar_53[6][145] , \_zy_simnet_tvar_53[6].label[136] );
tran (\_zy_simnet_tvar_53[6][144] , \_zy_simnet_tvar_53[6].label[135] );
tran (\_zy_simnet_tvar_53[6][143] , \_zy_simnet_tvar_53[6].label[134] );
tran (\_zy_simnet_tvar_53[6][142] , \_zy_simnet_tvar_53[6].label[133] );
tran (\_zy_simnet_tvar_53[6][141] , \_zy_simnet_tvar_53[6].label[132] );
tran (\_zy_simnet_tvar_53[6][140] , \_zy_simnet_tvar_53[6].label[131] );
tran (\_zy_simnet_tvar_53[6][139] , \_zy_simnet_tvar_53[6].label[130] );
tran (\_zy_simnet_tvar_53[6][138] , \_zy_simnet_tvar_53[6].label[129] );
tran (\_zy_simnet_tvar_53[6][137] , \_zy_simnet_tvar_53[6].label[128] );
tran (\_zy_simnet_tvar_53[6][136] , \_zy_simnet_tvar_53[6].label[127] );
tran (\_zy_simnet_tvar_53[6][135] , \_zy_simnet_tvar_53[6].label[126] );
tran (\_zy_simnet_tvar_53[6][134] , \_zy_simnet_tvar_53[6].label[125] );
tran (\_zy_simnet_tvar_53[6][133] , \_zy_simnet_tvar_53[6].label[124] );
tran (\_zy_simnet_tvar_53[6][132] , \_zy_simnet_tvar_53[6].label[123] );
tran (\_zy_simnet_tvar_53[6][131] , \_zy_simnet_tvar_53[6].label[122] );
tran (\_zy_simnet_tvar_53[6][130] , \_zy_simnet_tvar_53[6].label[121] );
tran (\_zy_simnet_tvar_53[6][129] , \_zy_simnet_tvar_53[6].label[120] );
tran (\_zy_simnet_tvar_53[6][128] , \_zy_simnet_tvar_53[6].label[119] );
tran (\_zy_simnet_tvar_53[6][127] , \_zy_simnet_tvar_53[6].label[118] );
tran (\_zy_simnet_tvar_53[6][126] , \_zy_simnet_tvar_53[6].label[117] );
tran (\_zy_simnet_tvar_53[6][125] , \_zy_simnet_tvar_53[6].label[116] );
tran (\_zy_simnet_tvar_53[6][124] , \_zy_simnet_tvar_53[6].label[115] );
tran (\_zy_simnet_tvar_53[6][123] , \_zy_simnet_tvar_53[6].label[114] );
tran (\_zy_simnet_tvar_53[6][122] , \_zy_simnet_tvar_53[6].label[113] );
tran (\_zy_simnet_tvar_53[6][121] , \_zy_simnet_tvar_53[6].label[112] );
tran (\_zy_simnet_tvar_53[6][120] , \_zy_simnet_tvar_53[6].label[111] );
tran (\_zy_simnet_tvar_53[6][119] , \_zy_simnet_tvar_53[6].label[110] );
tran (\_zy_simnet_tvar_53[6][118] , \_zy_simnet_tvar_53[6].label[109] );
tran (\_zy_simnet_tvar_53[6][117] , \_zy_simnet_tvar_53[6].label[108] );
tran (\_zy_simnet_tvar_53[6][116] , \_zy_simnet_tvar_53[6].label[107] );
tran (\_zy_simnet_tvar_53[6][115] , \_zy_simnet_tvar_53[6].label[106] );
tran (\_zy_simnet_tvar_53[6][114] , \_zy_simnet_tvar_53[6].label[105] );
tran (\_zy_simnet_tvar_53[6][113] , \_zy_simnet_tvar_53[6].label[104] );
tran (\_zy_simnet_tvar_53[6][112] , \_zy_simnet_tvar_53[6].label[103] );
tran (\_zy_simnet_tvar_53[6][111] , \_zy_simnet_tvar_53[6].label[102] );
tran (\_zy_simnet_tvar_53[6][110] , \_zy_simnet_tvar_53[6].label[101] );
tran (\_zy_simnet_tvar_53[6][109] , \_zy_simnet_tvar_53[6].label[100] );
tran (\_zy_simnet_tvar_53[6][108] , \_zy_simnet_tvar_53[6].label[99] );
tran (\_zy_simnet_tvar_53[6][107] , \_zy_simnet_tvar_53[6].label[98] );
tran (\_zy_simnet_tvar_53[6][106] , \_zy_simnet_tvar_53[6].label[97] );
tran (\_zy_simnet_tvar_53[6][105] , \_zy_simnet_tvar_53[6].label[96] );
tran (\_zy_simnet_tvar_53[6][104] , \_zy_simnet_tvar_53[6].label[95] );
tran (\_zy_simnet_tvar_53[6][103] , \_zy_simnet_tvar_53[6].label[94] );
tran (\_zy_simnet_tvar_53[6][102] , \_zy_simnet_tvar_53[6].label[93] );
tran (\_zy_simnet_tvar_53[6][101] , \_zy_simnet_tvar_53[6].label[92] );
tran (\_zy_simnet_tvar_53[6][100] , \_zy_simnet_tvar_53[6].label[91] );
tran (\_zy_simnet_tvar_53[6][99] , \_zy_simnet_tvar_53[6].label[90] );
tran (\_zy_simnet_tvar_53[6][98] , \_zy_simnet_tvar_53[6].label[89] );
tran (\_zy_simnet_tvar_53[6][97] , \_zy_simnet_tvar_53[6].label[88] );
tran (\_zy_simnet_tvar_53[6][96] , \_zy_simnet_tvar_53[6].label[87] );
tran (\_zy_simnet_tvar_53[6][95] , \_zy_simnet_tvar_53[6].label[86] );
tran (\_zy_simnet_tvar_53[6][94] , \_zy_simnet_tvar_53[6].label[85] );
tran (\_zy_simnet_tvar_53[6][93] , \_zy_simnet_tvar_53[6].label[84] );
tran (\_zy_simnet_tvar_53[6][92] , \_zy_simnet_tvar_53[6].label[83] );
tran (\_zy_simnet_tvar_53[6][91] , \_zy_simnet_tvar_53[6].label[82] );
tran (\_zy_simnet_tvar_53[6][90] , \_zy_simnet_tvar_53[6].label[81] );
tran (\_zy_simnet_tvar_53[6][89] , \_zy_simnet_tvar_53[6].label[80] );
tran (\_zy_simnet_tvar_53[6][88] , \_zy_simnet_tvar_53[6].label[79] );
tran (\_zy_simnet_tvar_53[6][87] , \_zy_simnet_tvar_53[6].label[78] );
tran (\_zy_simnet_tvar_53[6][86] , \_zy_simnet_tvar_53[6].label[77] );
tran (\_zy_simnet_tvar_53[6][85] , \_zy_simnet_tvar_53[6].label[76] );
tran (\_zy_simnet_tvar_53[6][84] , \_zy_simnet_tvar_53[6].label[75] );
tran (\_zy_simnet_tvar_53[6][83] , \_zy_simnet_tvar_53[6].label[74] );
tran (\_zy_simnet_tvar_53[6][82] , \_zy_simnet_tvar_53[6].label[73] );
tran (\_zy_simnet_tvar_53[6][81] , \_zy_simnet_tvar_53[6].label[72] );
tran (\_zy_simnet_tvar_53[6][80] , \_zy_simnet_tvar_53[6].label[71] );
tran (\_zy_simnet_tvar_53[6][79] , \_zy_simnet_tvar_53[6].label[70] );
tran (\_zy_simnet_tvar_53[6][78] , \_zy_simnet_tvar_53[6].label[69] );
tran (\_zy_simnet_tvar_53[6][77] , \_zy_simnet_tvar_53[6].label[68] );
tran (\_zy_simnet_tvar_53[6][76] , \_zy_simnet_tvar_53[6].label[67] );
tran (\_zy_simnet_tvar_53[6][75] , \_zy_simnet_tvar_53[6].label[66] );
tran (\_zy_simnet_tvar_53[6][74] , \_zy_simnet_tvar_53[6].label[65] );
tran (\_zy_simnet_tvar_53[6][73] , \_zy_simnet_tvar_53[6].label[64] );
tran (\_zy_simnet_tvar_53[6][72] , \_zy_simnet_tvar_53[6].label[63] );
tran (\_zy_simnet_tvar_53[6][71] , \_zy_simnet_tvar_53[6].label[62] );
tran (\_zy_simnet_tvar_53[6][70] , \_zy_simnet_tvar_53[6].label[61] );
tran (\_zy_simnet_tvar_53[6][69] , \_zy_simnet_tvar_53[6].label[60] );
tran (\_zy_simnet_tvar_53[6][68] , \_zy_simnet_tvar_53[6].label[59] );
tran (\_zy_simnet_tvar_53[6][67] , \_zy_simnet_tvar_53[6].label[58] );
tran (\_zy_simnet_tvar_53[6][66] , \_zy_simnet_tvar_53[6].label[57] );
tran (\_zy_simnet_tvar_53[6][65] , \_zy_simnet_tvar_53[6].label[56] );
tran (\_zy_simnet_tvar_53[6][64] , \_zy_simnet_tvar_53[6].label[55] );
tran (\_zy_simnet_tvar_53[6][63] , \_zy_simnet_tvar_53[6].label[54] );
tran (\_zy_simnet_tvar_53[6][62] , \_zy_simnet_tvar_53[6].label[53] );
tran (\_zy_simnet_tvar_53[6][61] , \_zy_simnet_tvar_53[6].label[52] );
tran (\_zy_simnet_tvar_53[6][60] , \_zy_simnet_tvar_53[6].label[51] );
tran (\_zy_simnet_tvar_53[6][59] , \_zy_simnet_tvar_53[6].label[50] );
tran (\_zy_simnet_tvar_53[6][58] , \_zy_simnet_tvar_53[6].label[49] );
tran (\_zy_simnet_tvar_53[6][57] , \_zy_simnet_tvar_53[6].label[48] );
tran (\_zy_simnet_tvar_53[6][56] , \_zy_simnet_tvar_53[6].label[47] );
tran (\_zy_simnet_tvar_53[6][55] , \_zy_simnet_tvar_53[6].label[46] );
tran (\_zy_simnet_tvar_53[6][54] , \_zy_simnet_tvar_53[6].label[45] );
tran (\_zy_simnet_tvar_53[6][53] , \_zy_simnet_tvar_53[6].label[44] );
tran (\_zy_simnet_tvar_53[6][52] , \_zy_simnet_tvar_53[6].label[43] );
tran (\_zy_simnet_tvar_53[6][51] , \_zy_simnet_tvar_53[6].label[42] );
tran (\_zy_simnet_tvar_53[6][50] , \_zy_simnet_tvar_53[6].label[41] );
tran (\_zy_simnet_tvar_53[6][49] , \_zy_simnet_tvar_53[6].label[40] );
tran (\_zy_simnet_tvar_53[6][48] , \_zy_simnet_tvar_53[6].label[39] );
tran (\_zy_simnet_tvar_53[6][47] , \_zy_simnet_tvar_53[6].label[38] );
tran (\_zy_simnet_tvar_53[6][46] , \_zy_simnet_tvar_53[6].label[37] );
tran (\_zy_simnet_tvar_53[6][45] , \_zy_simnet_tvar_53[6].label[36] );
tran (\_zy_simnet_tvar_53[6][44] , \_zy_simnet_tvar_53[6].label[35] );
tran (\_zy_simnet_tvar_53[6][43] , \_zy_simnet_tvar_53[6].label[34] );
tran (\_zy_simnet_tvar_53[6][42] , \_zy_simnet_tvar_53[6].label[33] );
tran (\_zy_simnet_tvar_53[6][41] , \_zy_simnet_tvar_53[6].label[32] );
tran (\_zy_simnet_tvar_53[6][40] , \_zy_simnet_tvar_53[6].label[31] );
tran (\_zy_simnet_tvar_53[6][39] , \_zy_simnet_tvar_53[6].label[30] );
tran (\_zy_simnet_tvar_53[6][38] , \_zy_simnet_tvar_53[6].label[29] );
tran (\_zy_simnet_tvar_53[6][37] , \_zy_simnet_tvar_53[6].label[28] );
tran (\_zy_simnet_tvar_53[6][36] , \_zy_simnet_tvar_53[6].label[27] );
tran (\_zy_simnet_tvar_53[6][35] , \_zy_simnet_tvar_53[6].label[26] );
tran (\_zy_simnet_tvar_53[6][34] , \_zy_simnet_tvar_53[6].label[25] );
tran (\_zy_simnet_tvar_53[6][33] , \_zy_simnet_tvar_53[6].label[24] );
tran (\_zy_simnet_tvar_53[6][32] , \_zy_simnet_tvar_53[6].label[23] );
tran (\_zy_simnet_tvar_53[6][31] , \_zy_simnet_tvar_53[6].label[22] );
tran (\_zy_simnet_tvar_53[6][30] , \_zy_simnet_tvar_53[6].label[21] );
tran (\_zy_simnet_tvar_53[6][29] , \_zy_simnet_tvar_53[6].label[20] );
tran (\_zy_simnet_tvar_53[6][28] , \_zy_simnet_tvar_53[6].label[19] );
tran (\_zy_simnet_tvar_53[6][27] , \_zy_simnet_tvar_53[6].label[18] );
tran (\_zy_simnet_tvar_53[6][26] , \_zy_simnet_tvar_53[6].label[17] );
tran (\_zy_simnet_tvar_53[6][25] , \_zy_simnet_tvar_53[6].label[16] );
tran (\_zy_simnet_tvar_53[6][24] , \_zy_simnet_tvar_53[6].label[15] );
tran (\_zy_simnet_tvar_53[6][23] , \_zy_simnet_tvar_53[6].label[14] );
tran (\_zy_simnet_tvar_53[6][22] , \_zy_simnet_tvar_53[6].label[13] );
tran (\_zy_simnet_tvar_53[6][21] , \_zy_simnet_tvar_53[6].label[12] );
tran (\_zy_simnet_tvar_53[6][20] , \_zy_simnet_tvar_53[6].label[11] );
tran (\_zy_simnet_tvar_53[6][19] , \_zy_simnet_tvar_53[6].label[10] );
tran (\_zy_simnet_tvar_53[6][18] , \_zy_simnet_tvar_53[6].label[9] );
tran (\_zy_simnet_tvar_53[6][17] , \_zy_simnet_tvar_53[6].label[8] );
tran (\_zy_simnet_tvar_53[6][16] , \_zy_simnet_tvar_53[6].label[7] );
tran (\_zy_simnet_tvar_53[6][15] , \_zy_simnet_tvar_53[6].label[6] );
tran (\_zy_simnet_tvar_53[6][14] , \_zy_simnet_tvar_53[6].label[5] );
tran (\_zy_simnet_tvar_53[6][13] , \_zy_simnet_tvar_53[6].label[4] );
tran (\_zy_simnet_tvar_53[6][12] , \_zy_simnet_tvar_53[6].label[3] );
tran (\_zy_simnet_tvar_53[6][11] , \_zy_simnet_tvar_53[6].label[2] );
tran (\_zy_simnet_tvar_53[6][10] , \_zy_simnet_tvar_53[6].label[1] );
tran (\_zy_simnet_tvar_53[6][9] , \_zy_simnet_tvar_53[6].label[0] );
tran (\_zy_simnet_tvar_53[6][8] , \_zy_simnet_tvar_53[6].delimiter_valid[0] );
tran (\_zy_simnet_tvar_53[6][7] , \_zy_simnet_tvar_53[6].delimiter[7] );
tran (\_zy_simnet_tvar_53[6][6] , \_zy_simnet_tvar_53[6].delimiter[6] );
tran (\_zy_simnet_tvar_53[6][5] , \_zy_simnet_tvar_53[6].delimiter[5] );
tran (\_zy_simnet_tvar_53[6][4] , \_zy_simnet_tvar_53[6].delimiter[4] );
tran (\_zy_simnet_tvar_53[6][3] , \_zy_simnet_tvar_53[6].delimiter[3] );
tran (\_zy_simnet_tvar_53[6][2] , \_zy_simnet_tvar_53[6].delimiter[2] );
tran (\_zy_simnet_tvar_53[6][1] , \_zy_simnet_tvar_53[6].delimiter[1] );
tran (\_zy_simnet_tvar_53[6][0] , \_zy_simnet_tvar_53[6].delimiter[0] );
tran (\_zy_simnet_tvar_53[5][271] , \_zy_simnet_tvar_53[5].guid_size[0] );
tran (\_zy_simnet_tvar_53[5][270] , \_zy_simnet_tvar_53[5].label_size[5] );
tran (\_zy_simnet_tvar_53[5][269] , \_zy_simnet_tvar_53[5].label_size[4] );
tran (\_zy_simnet_tvar_53[5][268] , \_zy_simnet_tvar_53[5].label_size[3] );
tran (\_zy_simnet_tvar_53[5][267] , \_zy_simnet_tvar_53[5].label_size[2] );
tran (\_zy_simnet_tvar_53[5][266] , \_zy_simnet_tvar_53[5].label_size[1] );
tran (\_zy_simnet_tvar_53[5][265] , \_zy_simnet_tvar_53[5].label_size[0] );
tran (\_zy_simnet_tvar_53[5][264] , \_zy_simnet_tvar_53[5].label[255] );
tran (\_zy_simnet_tvar_53[5][263] , \_zy_simnet_tvar_53[5].label[254] );
tran (\_zy_simnet_tvar_53[5][262] , \_zy_simnet_tvar_53[5].label[253] );
tran (\_zy_simnet_tvar_53[5][261] , \_zy_simnet_tvar_53[5].label[252] );
tran (\_zy_simnet_tvar_53[5][260] , \_zy_simnet_tvar_53[5].label[251] );
tran (\_zy_simnet_tvar_53[5][259] , \_zy_simnet_tvar_53[5].label[250] );
tran (\_zy_simnet_tvar_53[5][258] , \_zy_simnet_tvar_53[5].label[249] );
tran (\_zy_simnet_tvar_53[5][257] , \_zy_simnet_tvar_53[5].label[248] );
tran (\_zy_simnet_tvar_53[5][256] , \_zy_simnet_tvar_53[5].label[247] );
tran (\_zy_simnet_tvar_53[5][255] , \_zy_simnet_tvar_53[5].label[246] );
tran (\_zy_simnet_tvar_53[5][254] , \_zy_simnet_tvar_53[5].label[245] );
tran (\_zy_simnet_tvar_53[5][253] , \_zy_simnet_tvar_53[5].label[244] );
tran (\_zy_simnet_tvar_53[5][252] , \_zy_simnet_tvar_53[5].label[243] );
tran (\_zy_simnet_tvar_53[5][251] , \_zy_simnet_tvar_53[5].label[242] );
tran (\_zy_simnet_tvar_53[5][250] , \_zy_simnet_tvar_53[5].label[241] );
tran (\_zy_simnet_tvar_53[5][249] , \_zy_simnet_tvar_53[5].label[240] );
tran (\_zy_simnet_tvar_53[5][248] , \_zy_simnet_tvar_53[5].label[239] );
tran (\_zy_simnet_tvar_53[5][247] , \_zy_simnet_tvar_53[5].label[238] );
tran (\_zy_simnet_tvar_53[5][246] , \_zy_simnet_tvar_53[5].label[237] );
tran (\_zy_simnet_tvar_53[5][245] , \_zy_simnet_tvar_53[5].label[236] );
tran (\_zy_simnet_tvar_53[5][244] , \_zy_simnet_tvar_53[5].label[235] );
tran (\_zy_simnet_tvar_53[5][243] , \_zy_simnet_tvar_53[5].label[234] );
tran (\_zy_simnet_tvar_53[5][242] , \_zy_simnet_tvar_53[5].label[233] );
tran (\_zy_simnet_tvar_53[5][241] , \_zy_simnet_tvar_53[5].label[232] );
tran (\_zy_simnet_tvar_53[5][240] , \_zy_simnet_tvar_53[5].label[231] );
tran (\_zy_simnet_tvar_53[5][239] , \_zy_simnet_tvar_53[5].label[230] );
tran (\_zy_simnet_tvar_53[5][238] , \_zy_simnet_tvar_53[5].label[229] );
tran (\_zy_simnet_tvar_53[5][237] , \_zy_simnet_tvar_53[5].label[228] );
tran (\_zy_simnet_tvar_53[5][236] , \_zy_simnet_tvar_53[5].label[227] );
tran (\_zy_simnet_tvar_53[5][235] , \_zy_simnet_tvar_53[5].label[226] );
tran (\_zy_simnet_tvar_53[5][234] , \_zy_simnet_tvar_53[5].label[225] );
tran (\_zy_simnet_tvar_53[5][233] , \_zy_simnet_tvar_53[5].label[224] );
tran (\_zy_simnet_tvar_53[5][232] , \_zy_simnet_tvar_53[5].label[223] );
tran (\_zy_simnet_tvar_53[5][231] , \_zy_simnet_tvar_53[5].label[222] );
tran (\_zy_simnet_tvar_53[5][230] , \_zy_simnet_tvar_53[5].label[221] );
tran (\_zy_simnet_tvar_53[5][229] , \_zy_simnet_tvar_53[5].label[220] );
tran (\_zy_simnet_tvar_53[5][228] , \_zy_simnet_tvar_53[5].label[219] );
tran (\_zy_simnet_tvar_53[5][227] , \_zy_simnet_tvar_53[5].label[218] );
tran (\_zy_simnet_tvar_53[5][226] , \_zy_simnet_tvar_53[5].label[217] );
tran (\_zy_simnet_tvar_53[5][225] , \_zy_simnet_tvar_53[5].label[216] );
tran (\_zy_simnet_tvar_53[5][224] , \_zy_simnet_tvar_53[5].label[215] );
tran (\_zy_simnet_tvar_53[5][223] , \_zy_simnet_tvar_53[5].label[214] );
tran (\_zy_simnet_tvar_53[5][222] , \_zy_simnet_tvar_53[5].label[213] );
tran (\_zy_simnet_tvar_53[5][221] , \_zy_simnet_tvar_53[5].label[212] );
tran (\_zy_simnet_tvar_53[5][220] , \_zy_simnet_tvar_53[5].label[211] );
tran (\_zy_simnet_tvar_53[5][219] , \_zy_simnet_tvar_53[5].label[210] );
tran (\_zy_simnet_tvar_53[5][218] , \_zy_simnet_tvar_53[5].label[209] );
tran (\_zy_simnet_tvar_53[5][217] , \_zy_simnet_tvar_53[5].label[208] );
tran (\_zy_simnet_tvar_53[5][216] , \_zy_simnet_tvar_53[5].label[207] );
tran (\_zy_simnet_tvar_53[5][215] , \_zy_simnet_tvar_53[5].label[206] );
tran (\_zy_simnet_tvar_53[5][214] , \_zy_simnet_tvar_53[5].label[205] );
tran (\_zy_simnet_tvar_53[5][213] , \_zy_simnet_tvar_53[5].label[204] );
tran (\_zy_simnet_tvar_53[5][212] , \_zy_simnet_tvar_53[5].label[203] );
tran (\_zy_simnet_tvar_53[5][211] , \_zy_simnet_tvar_53[5].label[202] );
tran (\_zy_simnet_tvar_53[5][210] , \_zy_simnet_tvar_53[5].label[201] );
tran (\_zy_simnet_tvar_53[5][209] , \_zy_simnet_tvar_53[5].label[200] );
tran (\_zy_simnet_tvar_53[5][208] , \_zy_simnet_tvar_53[5].label[199] );
tran (\_zy_simnet_tvar_53[5][207] , \_zy_simnet_tvar_53[5].label[198] );
tran (\_zy_simnet_tvar_53[5][206] , \_zy_simnet_tvar_53[5].label[197] );
tran (\_zy_simnet_tvar_53[5][205] , \_zy_simnet_tvar_53[5].label[196] );
tran (\_zy_simnet_tvar_53[5][204] , \_zy_simnet_tvar_53[5].label[195] );
tran (\_zy_simnet_tvar_53[5][203] , \_zy_simnet_tvar_53[5].label[194] );
tran (\_zy_simnet_tvar_53[5][202] , \_zy_simnet_tvar_53[5].label[193] );
tran (\_zy_simnet_tvar_53[5][201] , \_zy_simnet_tvar_53[5].label[192] );
tran (\_zy_simnet_tvar_53[5][200] , \_zy_simnet_tvar_53[5].label[191] );
tran (\_zy_simnet_tvar_53[5][199] , \_zy_simnet_tvar_53[5].label[190] );
tran (\_zy_simnet_tvar_53[5][198] , \_zy_simnet_tvar_53[5].label[189] );
tran (\_zy_simnet_tvar_53[5][197] , \_zy_simnet_tvar_53[5].label[188] );
tran (\_zy_simnet_tvar_53[5][196] , \_zy_simnet_tvar_53[5].label[187] );
tran (\_zy_simnet_tvar_53[5][195] , \_zy_simnet_tvar_53[5].label[186] );
tran (\_zy_simnet_tvar_53[5][194] , \_zy_simnet_tvar_53[5].label[185] );
tran (\_zy_simnet_tvar_53[5][193] , \_zy_simnet_tvar_53[5].label[184] );
tran (\_zy_simnet_tvar_53[5][192] , \_zy_simnet_tvar_53[5].label[183] );
tran (\_zy_simnet_tvar_53[5][191] , \_zy_simnet_tvar_53[5].label[182] );
tran (\_zy_simnet_tvar_53[5][190] , \_zy_simnet_tvar_53[5].label[181] );
tran (\_zy_simnet_tvar_53[5][189] , \_zy_simnet_tvar_53[5].label[180] );
tran (\_zy_simnet_tvar_53[5][188] , \_zy_simnet_tvar_53[5].label[179] );
tran (\_zy_simnet_tvar_53[5][187] , \_zy_simnet_tvar_53[5].label[178] );
tran (\_zy_simnet_tvar_53[5][186] , \_zy_simnet_tvar_53[5].label[177] );
tran (\_zy_simnet_tvar_53[5][185] , \_zy_simnet_tvar_53[5].label[176] );
tran (\_zy_simnet_tvar_53[5][184] , \_zy_simnet_tvar_53[5].label[175] );
tran (\_zy_simnet_tvar_53[5][183] , \_zy_simnet_tvar_53[5].label[174] );
tran (\_zy_simnet_tvar_53[5][182] , \_zy_simnet_tvar_53[5].label[173] );
tran (\_zy_simnet_tvar_53[5][181] , \_zy_simnet_tvar_53[5].label[172] );
tran (\_zy_simnet_tvar_53[5][180] , \_zy_simnet_tvar_53[5].label[171] );
tran (\_zy_simnet_tvar_53[5][179] , \_zy_simnet_tvar_53[5].label[170] );
tran (\_zy_simnet_tvar_53[5][178] , \_zy_simnet_tvar_53[5].label[169] );
tran (\_zy_simnet_tvar_53[5][177] , \_zy_simnet_tvar_53[5].label[168] );
tran (\_zy_simnet_tvar_53[5][176] , \_zy_simnet_tvar_53[5].label[167] );
tran (\_zy_simnet_tvar_53[5][175] , \_zy_simnet_tvar_53[5].label[166] );
tran (\_zy_simnet_tvar_53[5][174] , \_zy_simnet_tvar_53[5].label[165] );
tran (\_zy_simnet_tvar_53[5][173] , \_zy_simnet_tvar_53[5].label[164] );
tran (\_zy_simnet_tvar_53[5][172] , \_zy_simnet_tvar_53[5].label[163] );
tran (\_zy_simnet_tvar_53[5][171] , \_zy_simnet_tvar_53[5].label[162] );
tran (\_zy_simnet_tvar_53[5][170] , \_zy_simnet_tvar_53[5].label[161] );
tran (\_zy_simnet_tvar_53[5][169] , \_zy_simnet_tvar_53[5].label[160] );
tran (\_zy_simnet_tvar_53[5][168] , \_zy_simnet_tvar_53[5].label[159] );
tran (\_zy_simnet_tvar_53[5][167] , \_zy_simnet_tvar_53[5].label[158] );
tran (\_zy_simnet_tvar_53[5][166] , \_zy_simnet_tvar_53[5].label[157] );
tran (\_zy_simnet_tvar_53[5][165] , \_zy_simnet_tvar_53[5].label[156] );
tran (\_zy_simnet_tvar_53[5][164] , \_zy_simnet_tvar_53[5].label[155] );
tran (\_zy_simnet_tvar_53[5][163] , \_zy_simnet_tvar_53[5].label[154] );
tran (\_zy_simnet_tvar_53[5][162] , \_zy_simnet_tvar_53[5].label[153] );
tran (\_zy_simnet_tvar_53[5][161] , \_zy_simnet_tvar_53[5].label[152] );
tran (\_zy_simnet_tvar_53[5][160] , \_zy_simnet_tvar_53[5].label[151] );
tran (\_zy_simnet_tvar_53[5][159] , \_zy_simnet_tvar_53[5].label[150] );
tran (\_zy_simnet_tvar_53[5][158] , \_zy_simnet_tvar_53[5].label[149] );
tran (\_zy_simnet_tvar_53[5][157] , \_zy_simnet_tvar_53[5].label[148] );
tran (\_zy_simnet_tvar_53[5][156] , \_zy_simnet_tvar_53[5].label[147] );
tran (\_zy_simnet_tvar_53[5][155] , \_zy_simnet_tvar_53[5].label[146] );
tran (\_zy_simnet_tvar_53[5][154] , \_zy_simnet_tvar_53[5].label[145] );
tran (\_zy_simnet_tvar_53[5][153] , \_zy_simnet_tvar_53[5].label[144] );
tran (\_zy_simnet_tvar_53[5][152] , \_zy_simnet_tvar_53[5].label[143] );
tran (\_zy_simnet_tvar_53[5][151] , \_zy_simnet_tvar_53[5].label[142] );
tran (\_zy_simnet_tvar_53[5][150] , \_zy_simnet_tvar_53[5].label[141] );
tran (\_zy_simnet_tvar_53[5][149] , \_zy_simnet_tvar_53[5].label[140] );
tran (\_zy_simnet_tvar_53[5][148] , \_zy_simnet_tvar_53[5].label[139] );
tran (\_zy_simnet_tvar_53[5][147] , \_zy_simnet_tvar_53[5].label[138] );
tran (\_zy_simnet_tvar_53[5][146] , \_zy_simnet_tvar_53[5].label[137] );
tran (\_zy_simnet_tvar_53[5][145] , \_zy_simnet_tvar_53[5].label[136] );
tran (\_zy_simnet_tvar_53[5][144] , \_zy_simnet_tvar_53[5].label[135] );
tran (\_zy_simnet_tvar_53[5][143] , \_zy_simnet_tvar_53[5].label[134] );
tran (\_zy_simnet_tvar_53[5][142] , \_zy_simnet_tvar_53[5].label[133] );
tran (\_zy_simnet_tvar_53[5][141] , \_zy_simnet_tvar_53[5].label[132] );
tran (\_zy_simnet_tvar_53[5][140] , \_zy_simnet_tvar_53[5].label[131] );
tran (\_zy_simnet_tvar_53[5][139] , \_zy_simnet_tvar_53[5].label[130] );
tran (\_zy_simnet_tvar_53[5][138] , \_zy_simnet_tvar_53[5].label[129] );
tran (\_zy_simnet_tvar_53[5][137] , \_zy_simnet_tvar_53[5].label[128] );
tran (\_zy_simnet_tvar_53[5][136] , \_zy_simnet_tvar_53[5].label[127] );
tran (\_zy_simnet_tvar_53[5][135] , \_zy_simnet_tvar_53[5].label[126] );
tran (\_zy_simnet_tvar_53[5][134] , \_zy_simnet_tvar_53[5].label[125] );
tran (\_zy_simnet_tvar_53[5][133] , \_zy_simnet_tvar_53[5].label[124] );
tran (\_zy_simnet_tvar_53[5][132] , \_zy_simnet_tvar_53[5].label[123] );
tran (\_zy_simnet_tvar_53[5][131] , \_zy_simnet_tvar_53[5].label[122] );
tran (\_zy_simnet_tvar_53[5][130] , \_zy_simnet_tvar_53[5].label[121] );
tran (\_zy_simnet_tvar_53[5][129] , \_zy_simnet_tvar_53[5].label[120] );
tran (\_zy_simnet_tvar_53[5][128] , \_zy_simnet_tvar_53[5].label[119] );
tran (\_zy_simnet_tvar_53[5][127] , \_zy_simnet_tvar_53[5].label[118] );
tran (\_zy_simnet_tvar_53[5][126] , \_zy_simnet_tvar_53[5].label[117] );
tran (\_zy_simnet_tvar_53[5][125] , \_zy_simnet_tvar_53[5].label[116] );
tran (\_zy_simnet_tvar_53[5][124] , \_zy_simnet_tvar_53[5].label[115] );
tran (\_zy_simnet_tvar_53[5][123] , \_zy_simnet_tvar_53[5].label[114] );
tran (\_zy_simnet_tvar_53[5][122] , \_zy_simnet_tvar_53[5].label[113] );
tran (\_zy_simnet_tvar_53[5][121] , \_zy_simnet_tvar_53[5].label[112] );
tran (\_zy_simnet_tvar_53[5][120] , \_zy_simnet_tvar_53[5].label[111] );
tran (\_zy_simnet_tvar_53[5][119] , \_zy_simnet_tvar_53[5].label[110] );
tran (\_zy_simnet_tvar_53[5][118] , \_zy_simnet_tvar_53[5].label[109] );
tran (\_zy_simnet_tvar_53[5][117] , \_zy_simnet_tvar_53[5].label[108] );
tran (\_zy_simnet_tvar_53[5][116] , \_zy_simnet_tvar_53[5].label[107] );
tran (\_zy_simnet_tvar_53[5][115] , \_zy_simnet_tvar_53[5].label[106] );
tran (\_zy_simnet_tvar_53[5][114] , \_zy_simnet_tvar_53[5].label[105] );
tran (\_zy_simnet_tvar_53[5][113] , \_zy_simnet_tvar_53[5].label[104] );
tran (\_zy_simnet_tvar_53[5][112] , \_zy_simnet_tvar_53[5].label[103] );
tran (\_zy_simnet_tvar_53[5][111] , \_zy_simnet_tvar_53[5].label[102] );
tran (\_zy_simnet_tvar_53[5][110] , \_zy_simnet_tvar_53[5].label[101] );
tran (\_zy_simnet_tvar_53[5][109] , \_zy_simnet_tvar_53[5].label[100] );
tran (\_zy_simnet_tvar_53[5][108] , \_zy_simnet_tvar_53[5].label[99] );
tran (\_zy_simnet_tvar_53[5][107] , \_zy_simnet_tvar_53[5].label[98] );
tran (\_zy_simnet_tvar_53[5][106] , \_zy_simnet_tvar_53[5].label[97] );
tran (\_zy_simnet_tvar_53[5][105] , \_zy_simnet_tvar_53[5].label[96] );
tran (\_zy_simnet_tvar_53[5][104] , \_zy_simnet_tvar_53[5].label[95] );
tran (\_zy_simnet_tvar_53[5][103] , \_zy_simnet_tvar_53[5].label[94] );
tran (\_zy_simnet_tvar_53[5][102] , \_zy_simnet_tvar_53[5].label[93] );
tran (\_zy_simnet_tvar_53[5][101] , \_zy_simnet_tvar_53[5].label[92] );
tran (\_zy_simnet_tvar_53[5][100] , \_zy_simnet_tvar_53[5].label[91] );
tran (\_zy_simnet_tvar_53[5][99] , \_zy_simnet_tvar_53[5].label[90] );
tran (\_zy_simnet_tvar_53[5][98] , \_zy_simnet_tvar_53[5].label[89] );
tran (\_zy_simnet_tvar_53[5][97] , \_zy_simnet_tvar_53[5].label[88] );
tran (\_zy_simnet_tvar_53[5][96] , \_zy_simnet_tvar_53[5].label[87] );
tran (\_zy_simnet_tvar_53[5][95] , \_zy_simnet_tvar_53[5].label[86] );
tran (\_zy_simnet_tvar_53[5][94] , \_zy_simnet_tvar_53[5].label[85] );
tran (\_zy_simnet_tvar_53[5][93] , \_zy_simnet_tvar_53[5].label[84] );
tran (\_zy_simnet_tvar_53[5][92] , \_zy_simnet_tvar_53[5].label[83] );
tran (\_zy_simnet_tvar_53[5][91] , \_zy_simnet_tvar_53[5].label[82] );
tran (\_zy_simnet_tvar_53[5][90] , \_zy_simnet_tvar_53[5].label[81] );
tran (\_zy_simnet_tvar_53[5][89] , \_zy_simnet_tvar_53[5].label[80] );
tran (\_zy_simnet_tvar_53[5][88] , \_zy_simnet_tvar_53[5].label[79] );
tran (\_zy_simnet_tvar_53[5][87] , \_zy_simnet_tvar_53[5].label[78] );
tran (\_zy_simnet_tvar_53[5][86] , \_zy_simnet_tvar_53[5].label[77] );
tran (\_zy_simnet_tvar_53[5][85] , \_zy_simnet_tvar_53[5].label[76] );
tran (\_zy_simnet_tvar_53[5][84] , \_zy_simnet_tvar_53[5].label[75] );
tran (\_zy_simnet_tvar_53[5][83] , \_zy_simnet_tvar_53[5].label[74] );
tran (\_zy_simnet_tvar_53[5][82] , \_zy_simnet_tvar_53[5].label[73] );
tran (\_zy_simnet_tvar_53[5][81] , \_zy_simnet_tvar_53[5].label[72] );
tran (\_zy_simnet_tvar_53[5][80] , \_zy_simnet_tvar_53[5].label[71] );
tran (\_zy_simnet_tvar_53[5][79] , \_zy_simnet_tvar_53[5].label[70] );
tran (\_zy_simnet_tvar_53[5][78] , \_zy_simnet_tvar_53[5].label[69] );
tran (\_zy_simnet_tvar_53[5][77] , \_zy_simnet_tvar_53[5].label[68] );
tran (\_zy_simnet_tvar_53[5][76] , \_zy_simnet_tvar_53[5].label[67] );
tran (\_zy_simnet_tvar_53[5][75] , \_zy_simnet_tvar_53[5].label[66] );
tran (\_zy_simnet_tvar_53[5][74] , \_zy_simnet_tvar_53[5].label[65] );
tran (\_zy_simnet_tvar_53[5][73] , \_zy_simnet_tvar_53[5].label[64] );
tran (\_zy_simnet_tvar_53[5][72] , \_zy_simnet_tvar_53[5].label[63] );
tran (\_zy_simnet_tvar_53[5][71] , \_zy_simnet_tvar_53[5].label[62] );
tran (\_zy_simnet_tvar_53[5][70] , \_zy_simnet_tvar_53[5].label[61] );
tran (\_zy_simnet_tvar_53[5][69] , \_zy_simnet_tvar_53[5].label[60] );
tran (\_zy_simnet_tvar_53[5][68] , \_zy_simnet_tvar_53[5].label[59] );
tran (\_zy_simnet_tvar_53[5][67] , \_zy_simnet_tvar_53[5].label[58] );
tran (\_zy_simnet_tvar_53[5][66] , \_zy_simnet_tvar_53[5].label[57] );
tran (\_zy_simnet_tvar_53[5][65] , \_zy_simnet_tvar_53[5].label[56] );
tran (\_zy_simnet_tvar_53[5][64] , \_zy_simnet_tvar_53[5].label[55] );
tran (\_zy_simnet_tvar_53[5][63] , \_zy_simnet_tvar_53[5].label[54] );
tran (\_zy_simnet_tvar_53[5][62] , \_zy_simnet_tvar_53[5].label[53] );
tran (\_zy_simnet_tvar_53[5][61] , \_zy_simnet_tvar_53[5].label[52] );
tran (\_zy_simnet_tvar_53[5][60] , \_zy_simnet_tvar_53[5].label[51] );
tran (\_zy_simnet_tvar_53[5][59] , \_zy_simnet_tvar_53[5].label[50] );
tran (\_zy_simnet_tvar_53[5][58] , \_zy_simnet_tvar_53[5].label[49] );
tran (\_zy_simnet_tvar_53[5][57] , \_zy_simnet_tvar_53[5].label[48] );
tran (\_zy_simnet_tvar_53[5][56] , \_zy_simnet_tvar_53[5].label[47] );
tran (\_zy_simnet_tvar_53[5][55] , \_zy_simnet_tvar_53[5].label[46] );
tran (\_zy_simnet_tvar_53[5][54] , \_zy_simnet_tvar_53[5].label[45] );
tran (\_zy_simnet_tvar_53[5][53] , \_zy_simnet_tvar_53[5].label[44] );
tran (\_zy_simnet_tvar_53[5][52] , \_zy_simnet_tvar_53[5].label[43] );
tran (\_zy_simnet_tvar_53[5][51] , \_zy_simnet_tvar_53[5].label[42] );
tran (\_zy_simnet_tvar_53[5][50] , \_zy_simnet_tvar_53[5].label[41] );
tran (\_zy_simnet_tvar_53[5][49] , \_zy_simnet_tvar_53[5].label[40] );
tran (\_zy_simnet_tvar_53[5][48] , \_zy_simnet_tvar_53[5].label[39] );
tran (\_zy_simnet_tvar_53[5][47] , \_zy_simnet_tvar_53[5].label[38] );
tran (\_zy_simnet_tvar_53[5][46] , \_zy_simnet_tvar_53[5].label[37] );
tran (\_zy_simnet_tvar_53[5][45] , \_zy_simnet_tvar_53[5].label[36] );
tran (\_zy_simnet_tvar_53[5][44] , \_zy_simnet_tvar_53[5].label[35] );
tran (\_zy_simnet_tvar_53[5][43] , \_zy_simnet_tvar_53[5].label[34] );
tran (\_zy_simnet_tvar_53[5][42] , \_zy_simnet_tvar_53[5].label[33] );
tran (\_zy_simnet_tvar_53[5][41] , \_zy_simnet_tvar_53[5].label[32] );
tran (\_zy_simnet_tvar_53[5][40] , \_zy_simnet_tvar_53[5].label[31] );
tran (\_zy_simnet_tvar_53[5][39] , \_zy_simnet_tvar_53[5].label[30] );
tran (\_zy_simnet_tvar_53[5][38] , \_zy_simnet_tvar_53[5].label[29] );
tran (\_zy_simnet_tvar_53[5][37] , \_zy_simnet_tvar_53[5].label[28] );
tran (\_zy_simnet_tvar_53[5][36] , \_zy_simnet_tvar_53[5].label[27] );
tran (\_zy_simnet_tvar_53[5][35] , \_zy_simnet_tvar_53[5].label[26] );
tran (\_zy_simnet_tvar_53[5][34] , \_zy_simnet_tvar_53[5].label[25] );
tran (\_zy_simnet_tvar_53[5][33] , \_zy_simnet_tvar_53[5].label[24] );
tran (\_zy_simnet_tvar_53[5][32] , \_zy_simnet_tvar_53[5].label[23] );
tran (\_zy_simnet_tvar_53[5][31] , \_zy_simnet_tvar_53[5].label[22] );
tran (\_zy_simnet_tvar_53[5][30] , \_zy_simnet_tvar_53[5].label[21] );
tran (\_zy_simnet_tvar_53[5][29] , \_zy_simnet_tvar_53[5].label[20] );
tran (\_zy_simnet_tvar_53[5][28] , \_zy_simnet_tvar_53[5].label[19] );
tran (\_zy_simnet_tvar_53[5][27] , \_zy_simnet_tvar_53[5].label[18] );
tran (\_zy_simnet_tvar_53[5][26] , \_zy_simnet_tvar_53[5].label[17] );
tran (\_zy_simnet_tvar_53[5][25] , \_zy_simnet_tvar_53[5].label[16] );
tran (\_zy_simnet_tvar_53[5][24] , \_zy_simnet_tvar_53[5].label[15] );
tran (\_zy_simnet_tvar_53[5][23] , \_zy_simnet_tvar_53[5].label[14] );
tran (\_zy_simnet_tvar_53[5][22] , \_zy_simnet_tvar_53[5].label[13] );
tran (\_zy_simnet_tvar_53[5][21] , \_zy_simnet_tvar_53[5].label[12] );
tran (\_zy_simnet_tvar_53[5][20] , \_zy_simnet_tvar_53[5].label[11] );
tran (\_zy_simnet_tvar_53[5][19] , \_zy_simnet_tvar_53[5].label[10] );
tran (\_zy_simnet_tvar_53[5][18] , \_zy_simnet_tvar_53[5].label[9] );
tran (\_zy_simnet_tvar_53[5][17] , \_zy_simnet_tvar_53[5].label[8] );
tran (\_zy_simnet_tvar_53[5][16] , \_zy_simnet_tvar_53[5].label[7] );
tran (\_zy_simnet_tvar_53[5][15] , \_zy_simnet_tvar_53[5].label[6] );
tran (\_zy_simnet_tvar_53[5][14] , \_zy_simnet_tvar_53[5].label[5] );
tran (\_zy_simnet_tvar_53[5][13] , \_zy_simnet_tvar_53[5].label[4] );
tran (\_zy_simnet_tvar_53[5][12] , \_zy_simnet_tvar_53[5].label[3] );
tran (\_zy_simnet_tvar_53[5][11] , \_zy_simnet_tvar_53[5].label[2] );
tran (\_zy_simnet_tvar_53[5][10] , \_zy_simnet_tvar_53[5].label[1] );
tran (\_zy_simnet_tvar_53[5][9] , \_zy_simnet_tvar_53[5].label[0] );
tran (\_zy_simnet_tvar_53[5][8] , \_zy_simnet_tvar_53[5].delimiter_valid[0] );
tran (\_zy_simnet_tvar_53[5][7] , \_zy_simnet_tvar_53[5].delimiter[7] );
tran (\_zy_simnet_tvar_53[5][6] , \_zy_simnet_tvar_53[5].delimiter[6] );
tran (\_zy_simnet_tvar_53[5][5] , \_zy_simnet_tvar_53[5].delimiter[5] );
tran (\_zy_simnet_tvar_53[5][4] , \_zy_simnet_tvar_53[5].delimiter[4] );
tran (\_zy_simnet_tvar_53[5][3] , \_zy_simnet_tvar_53[5].delimiter[3] );
tran (\_zy_simnet_tvar_53[5][2] , \_zy_simnet_tvar_53[5].delimiter[2] );
tran (\_zy_simnet_tvar_53[5][1] , \_zy_simnet_tvar_53[5].delimiter[1] );
tran (\_zy_simnet_tvar_53[5][0] , \_zy_simnet_tvar_53[5].delimiter[0] );
tran (\_zy_simnet_tvar_53[4][271] , \_zy_simnet_tvar_53[4].guid_size[0] );
tran (\_zy_simnet_tvar_53[4][270] , \_zy_simnet_tvar_53[4].label_size[5] );
tran (\_zy_simnet_tvar_53[4][269] , \_zy_simnet_tvar_53[4].label_size[4] );
tran (\_zy_simnet_tvar_53[4][268] , \_zy_simnet_tvar_53[4].label_size[3] );
tran (\_zy_simnet_tvar_53[4][267] , \_zy_simnet_tvar_53[4].label_size[2] );
tran (\_zy_simnet_tvar_53[4][266] , \_zy_simnet_tvar_53[4].label_size[1] );
tran (\_zy_simnet_tvar_53[4][265] , \_zy_simnet_tvar_53[4].label_size[0] );
tran (\_zy_simnet_tvar_53[4][264] , \_zy_simnet_tvar_53[4].label[255] );
tran (\_zy_simnet_tvar_53[4][263] , \_zy_simnet_tvar_53[4].label[254] );
tran (\_zy_simnet_tvar_53[4][262] , \_zy_simnet_tvar_53[4].label[253] );
tran (\_zy_simnet_tvar_53[4][261] , \_zy_simnet_tvar_53[4].label[252] );
tran (\_zy_simnet_tvar_53[4][260] , \_zy_simnet_tvar_53[4].label[251] );
tran (\_zy_simnet_tvar_53[4][259] , \_zy_simnet_tvar_53[4].label[250] );
tran (\_zy_simnet_tvar_53[4][258] , \_zy_simnet_tvar_53[4].label[249] );
tran (\_zy_simnet_tvar_53[4][257] , \_zy_simnet_tvar_53[4].label[248] );
tran (\_zy_simnet_tvar_53[4][256] , \_zy_simnet_tvar_53[4].label[247] );
tran (\_zy_simnet_tvar_53[4][255] , \_zy_simnet_tvar_53[4].label[246] );
tran (\_zy_simnet_tvar_53[4][254] , \_zy_simnet_tvar_53[4].label[245] );
tran (\_zy_simnet_tvar_53[4][253] , \_zy_simnet_tvar_53[4].label[244] );
tran (\_zy_simnet_tvar_53[4][252] , \_zy_simnet_tvar_53[4].label[243] );
tran (\_zy_simnet_tvar_53[4][251] , \_zy_simnet_tvar_53[4].label[242] );
tran (\_zy_simnet_tvar_53[4][250] , \_zy_simnet_tvar_53[4].label[241] );
tran (\_zy_simnet_tvar_53[4][249] , \_zy_simnet_tvar_53[4].label[240] );
tran (\_zy_simnet_tvar_53[4][248] , \_zy_simnet_tvar_53[4].label[239] );
tran (\_zy_simnet_tvar_53[4][247] , \_zy_simnet_tvar_53[4].label[238] );
tran (\_zy_simnet_tvar_53[4][246] , \_zy_simnet_tvar_53[4].label[237] );
tran (\_zy_simnet_tvar_53[4][245] , \_zy_simnet_tvar_53[4].label[236] );
tran (\_zy_simnet_tvar_53[4][244] , \_zy_simnet_tvar_53[4].label[235] );
tran (\_zy_simnet_tvar_53[4][243] , \_zy_simnet_tvar_53[4].label[234] );
tran (\_zy_simnet_tvar_53[4][242] , \_zy_simnet_tvar_53[4].label[233] );
tran (\_zy_simnet_tvar_53[4][241] , \_zy_simnet_tvar_53[4].label[232] );
tran (\_zy_simnet_tvar_53[4][240] , \_zy_simnet_tvar_53[4].label[231] );
tran (\_zy_simnet_tvar_53[4][239] , \_zy_simnet_tvar_53[4].label[230] );
tran (\_zy_simnet_tvar_53[4][238] , \_zy_simnet_tvar_53[4].label[229] );
tran (\_zy_simnet_tvar_53[4][237] , \_zy_simnet_tvar_53[4].label[228] );
tran (\_zy_simnet_tvar_53[4][236] , \_zy_simnet_tvar_53[4].label[227] );
tran (\_zy_simnet_tvar_53[4][235] , \_zy_simnet_tvar_53[4].label[226] );
tran (\_zy_simnet_tvar_53[4][234] , \_zy_simnet_tvar_53[4].label[225] );
tran (\_zy_simnet_tvar_53[4][233] , \_zy_simnet_tvar_53[4].label[224] );
tran (\_zy_simnet_tvar_53[4][232] , \_zy_simnet_tvar_53[4].label[223] );
tran (\_zy_simnet_tvar_53[4][231] , \_zy_simnet_tvar_53[4].label[222] );
tran (\_zy_simnet_tvar_53[4][230] , \_zy_simnet_tvar_53[4].label[221] );
tran (\_zy_simnet_tvar_53[4][229] , \_zy_simnet_tvar_53[4].label[220] );
tran (\_zy_simnet_tvar_53[4][228] , \_zy_simnet_tvar_53[4].label[219] );
tran (\_zy_simnet_tvar_53[4][227] , \_zy_simnet_tvar_53[4].label[218] );
tran (\_zy_simnet_tvar_53[4][226] , \_zy_simnet_tvar_53[4].label[217] );
tran (\_zy_simnet_tvar_53[4][225] , \_zy_simnet_tvar_53[4].label[216] );
tran (\_zy_simnet_tvar_53[4][224] , \_zy_simnet_tvar_53[4].label[215] );
tran (\_zy_simnet_tvar_53[4][223] , \_zy_simnet_tvar_53[4].label[214] );
tran (\_zy_simnet_tvar_53[4][222] , \_zy_simnet_tvar_53[4].label[213] );
tran (\_zy_simnet_tvar_53[4][221] , \_zy_simnet_tvar_53[4].label[212] );
tran (\_zy_simnet_tvar_53[4][220] , \_zy_simnet_tvar_53[4].label[211] );
tran (\_zy_simnet_tvar_53[4][219] , \_zy_simnet_tvar_53[4].label[210] );
tran (\_zy_simnet_tvar_53[4][218] , \_zy_simnet_tvar_53[4].label[209] );
tran (\_zy_simnet_tvar_53[4][217] , \_zy_simnet_tvar_53[4].label[208] );
tran (\_zy_simnet_tvar_53[4][216] , \_zy_simnet_tvar_53[4].label[207] );
tran (\_zy_simnet_tvar_53[4][215] , \_zy_simnet_tvar_53[4].label[206] );
tran (\_zy_simnet_tvar_53[4][214] , \_zy_simnet_tvar_53[4].label[205] );
tran (\_zy_simnet_tvar_53[4][213] , \_zy_simnet_tvar_53[4].label[204] );
tran (\_zy_simnet_tvar_53[4][212] , \_zy_simnet_tvar_53[4].label[203] );
tran (\_zy_simnet_tvar_53[4][211] , \_zy_simnet_tvar_53[4].label[202] );
tran (\_zy_simnet_tvar_53[4][210] , \_zy_simnet_tvar_53[4].label[201] );
tran (\_zy_simnet_tvar_53[4][209] , \_zy_simnet_tvar_53[4].label[200] );
tran (\_zy_simnet_tvar_53[4][208] , \_zy_simnet_tvar_53[4].label[199] );
tran (\_zy_simnet_tvar_53[4][207] , \_zy_simnet_tvar_53[4].label[198] );
tran (\_zy_simnet_tvar_53[4][206] , \_zy_simnet_tvar_53[4].label[197] );
tran (\_zy_simnet_tvar_53[4][205] , \_zy_simnet_tvar_53[4].label[196] );
tran (\_zy_simnet_tvar_53[4][204] , \_zy_simnet_tvar_53[4].label[195] );
tran (\_zy_simnet_tvar_53[4][203] , \_zy_simnet_tvar_53[4].label[194] );
tran (\_zy_simnet_tvar_53[4][202] , \_zy_simnet_tvar_53[4].label[193] );
tran (\_zy_simnet_tvar_53[4][201] , \_zy_simnet_tvar_53[4].label[192] );
tran (\_zy_simnet_tvar_53[4][200] , \_zy_simnet_tvar_53[4].label[191] );
tran (\_zy_simnet_tvar_53[4][199] , \_zy_simnet_tvar_53[4].label[190] );
tran (\_zy_simnet_tvar_53[4][198] , \_zy_simnet_tvar_53[4].label[189] );
tran (\_zy_simnet_tvar_53[4][197] , \_zy_simnet_tvar_53[4].label[188] );
tran (\_zy_simnet_tvar_53[4][196] , \_zy_simnet_tvar_53[4].label[187] );
tran (\_zy_simnet_tvar_53[4][195] , \_zy_simnet_tvar_53[4].label[186] );
tran (\_zy_simnet_tvar_53[4][194] , \_zy_simnet_tvar_53[4].label[185] );
tran (\_zy_simnet_tvar_53[4][193] , \_zy_simnet_tvar_53[4].label[184] );
tran (\_zy_simnet_tvar_53[4][192] , \_zy_simnet_tvar_53[4].label[183] );
tran (\_zy_simnet_tvar_53[4][191] , \_zy_simnet_tvar_53[4].label[182] );
tran (\_zy_simnet_tvar_53[4][190] , \_zy_simnet_tvar_53[4].label[181] );
tran (\_zy_simnet_tvar_53[4][189] , \_zy_simnet_tvar_53[4].label[180] );
tran (\_zy_simnet_tvar_53[4][188] , \_zy_simnet_tvar_53[4].label[179] );
tran (\_zy_simnet_tvar_53[4][187] , \_zy_simnet_tvar_53[4].label[178] );
tran (\_zy_simnet_tvar_53[4][186] , \_zy_simnet_tvar_53[4].label[177] );
tran (\_zy_simnet_tvar_53[4][185] , \_zy_simnet_tvar_53[4].label[176] );
tran (\_zy_simnet_tvar_53[4][184] , \_zy_simnet_tvar_53[4].label[175] );
tran (\_zy_simnet_tvar_53[4][183] , \_zy_simnet_tvar_53[4].label[174] );
tran (\_zy_simnet_tvar_53[4][182] , \_zy_simnet_tvar_53[4].label[173] );
tran (\_zy_simnet_tvar_53[4][181] , \_zy_simnet_tvar_53[4].label[172] );
tran (\_zy_simnet_tvar_53[4][180] , \_zy_simnet_tvar_53[4].label[171] );
tran (\_zy_simnet_tvar_53[4][179] , \_zy_simnet_tvar_53[4].label[170] );
tran (\_zy_simnet_tvar_53[4][178] , \_zy_simnet_tvar_53[4].label[169] );
tran (\_zy_simnet_tvar_53[4][177] , \_zy_simnet_tvar_53[4].label[168] );
tran (\_zy_simnet_tvar_53[4][176] , \_zy_simnet_tvar_53[4].label[167] );
tran (\_zy_simnet_tvar_53[4][175] , \_zy_simnet_tvar_53[4].label[166] );
tran (\_zy_simnet_tvar_53[4][174] , \_zy_simnet_tvar_53[4].label[165] );
tran (\_zy_simnet_tvar_53[4][173] , \_zy_simnet_tvar_53[4].label[164] );
tran (\_zy_simnet_tvar_53[4][172] , \_zy_simnet_tvar_53[4].label[163] );
tran (\_zy_simnet_tvar_53[4][171] , \_zy_simnet_tvar_53[4].label[162] );
tran (\_zy_simnet_tvar_53[4][170] , \_zy_simnet_tvar_53[4].label[161] );
tran (\_zy_simnet_tvar_53[4][169] , \_zy_simnet_tvar_53[4].label[160] );
tran (\_zy_simnet_tvar_53[4][168] , \_zy_simnet_tvar_53[4].label[159] );
tran (\_zy_simnet_tvar_53[4][167] , \_zy_simnet_tvar_53[4].label[158] );
tran (\_zy_simnet_tvar_53[4][166] , \_zy_simnet_tvar_53[4].label[157] );
tran (\_zy_simnet_tvar_53[4][165] , \_zy_simnet_tvar_53[4].label[156] );
tran (\_zy_simnet_tvar_53[4][164] , \_zy_simnet_tvar_53[4].label[155] );
tran (\_zy_simnet_tvar_53[4][163] , \_zy_simnet_tvar_53[4].label[154] );
tran (\_zy_simnet_tvar_53[4][162] , \_zy_simnet_tvar_53[4].label[153] );
tran (\_zy_simnet_tvar_53[4][161] , \_zy_simnet_tvar_53[4].label[152] );
tran (\_zy_simnet_tvar_53[4][160] , \_zy_simnet_tvar_53[4].label[151] );
tran (\_zy_simnet_tvar_53[4][159] , \_zy_simnet_tvar_53[4].label[150] );
tran (\_zy_simnet_tvar_53[4][158] , \_zy_simnet_tvar_53[4].label[149] );
tran (\_zy_simnet_tvar_53[4][157] , \_zy_simnet_tvar_53[4].label[148] );
tran (\_zy_simnet_tvar_53[4][156] , \_zy_simnet_tvar_53[4].label[147] );
tran (\_zy_simnet_tvar_53[4][155] , \_zy_simnet_tvar_53[4].label[146] );
tran (\_zy_simnet_tvar_53[4][154] , \_zy_simnet_tvar_53[4].label[145] );
tran (\_zy_simnet_tvar_53[4][153] , \_zy_simnet_tvar_53[4].label[144] );
tran (\_zy_simnet_tvar_53[4][152] , \_zy_simnet_tvar_53[4].label[143] );
tran (\_zy_simnet_tvar_53[4][151] , \_zy_simnet_tvar_53[4].label[142] );
tran (\_zy_simnet_tvar_53[4][150] , \_zy_simnet_tvar_53[4].label[141] );
tran (\_zy_simnet_tvar_53[4][149] , \_zy_simnet_tvar_53[4].label[140] );
tran (\_zy_simnet_tvar_53[4][148] , \_zy_simnet_tvar_53[4].label[139] );
tran (\_zy_simnet_tvar_53[4][147] , \_zy_simnet_tvar_53[4].label[138] );
tran (\_zy_simnet_tvar_53[4][146] , \_zy_simnet_tvar_53[4].label[137] );
tran (\_zy_simnet_tvar_53[4][145] , \_zy_simnet_tvar_53[4].label[136] );
tran (\_zy_simnet_tvar_53[4][144] , \_zy_simnet_tvar_53[4].label[135] );
tran (\_zy_simnet_tvar_53[4][143] , \_zy_simnet_tvar_53[4].label[134] );
tran (\_zy_simnet_tvar_53[4][142] , \_zy_simnet_tvar_53[4].label[133] );
tran (\_zy_simnet_tvar_53[4][141] , \_zy_simnet_tvar_53[4].label[132] );
tran (\_zy_simnet_tvar_53[4][140] , \_zy_simnet_tvar_53[4].label[131] );
tran (\_zy_simnet_tvar_53[4][139] , \_zy_simnet_tvar_53[4].label[130] );
tran (\_zy_simnet_tvar_53[4][138] , \_zy_simnet_tvar_53[4].label[129] );
tran (\_zy_simnet_tvar_53[4][137] , \_zy_simnet_tvar_53[4].label[128] );
tran (\_zy_simnet_tvar_53[4][136] , \_zy_simnet_tvar_53[4].label[127] );
tran (\_zy_simnet_tvar_53[4][135] , \_zy_simnet_tvar_53[4].label[126] );
tran (\_zy_simnet_tvar_53[4][134] , \_zy_simnet_tvar_53[4].label[125] );
tran (\_zy_simnet_tvar_53[4][133] , \_zy_simnet_tvar_53[4].label[124] );
tran (\_zy_simnet_tvar_53[4][132] , \_zy_simnet_tvar_53[4].label[123] );
tran (\_zy_simnet_tvar_53[4][131] , \_zy_simnet_tvar_53[4].label[122] );
tran (\_zy_simnet_tvar_53[4][130] , \_zy_simnet_tvar_53[4].label[121] );
tran (\_zy_simnet_tvar_53[4][129] , \_zy_simnet_tvar_53[4].label[120] );
tran (\_zy_simnet_tvar_53[4][128] , \_zy_simnet_tvar_53[4].label[119] );
tran (\_zy_simnet_tvar_53[4][127] , \_zy_simnet_tvar_53[4].label[118] );
tran (\_zy_simnet_tvar_53[4][126] , \_zy_simnet_tvar_53[4].label[117] );
tran (\_zy_simnet_tvar_53[4][125] , \_zy_simnet_tvar_53[4].label[116] );
tran (\_zy_simnet_tvar_53[4][124] , \_zy_simnet_tvar_53[4].label[115] );
tran (\_zy_simnet_tvar_53[4][123] , \_zy_simnet_tvar_53[4].label[114] );
tran (\_zy_simnet_tvar_53[4][122] , \_zy_simnet_tvar_53[4].label[113] );
tran (\_zy_simnet_tvar_53[4][121] , \_zy_simnet_tvar_53[4].label[112] );
tran (\_zy_simnet_tvar_53[4][120] , \_zy_simnet_tvar_53[4].label[111] );
tran (\_zy_simnet_tvar_53[4][119] , \_zy_simnet_tvar_53[4].label[110] );
tran (\_zy_simnet_tvar_53[4][118] , \_zy_simnet_tvar_53[4].label[109] );
tran (\_zy_simnet_tvar_53[4][117] , \_zy_simnet_tvar_53[4].label[108] );
tran (\_zy_simnet_tvar_53[4][116] , \_zy_simnet_tvar_53[4].label[107] );
tran (\_zy_simnet_tvar_53[4][115] , \_zy_simnet_tvar_53[4].label[106] );
tran (\_zy_simnet_tvar_53[4][114] , \_zy_simnet_tvar_53[4].label[105] );
tran (\_zy_simnet_tvar_53[4][113] , \_zy_simnet_tvar_53[4].label[104] );
tran (\_zy_simnet_tvar_53[4][112] , \_zy_simnet_tvar_53[4].label[103] );
tran (\_zy_simnet_tvar_53[4][111] , \_zy_simnet_tvar_53[4].label[102] );
tran (\_zy_simnet_tvar_53[4][110] , \_zy_simnet_tvar_53[4].label[101] );
tran (\_zy_simnet_tvar_53[4][109] , \_zy_simnet_tvar_53[4].label[100] );
tran (\_zy_simnet_tvar_53[4][108] , \_zy_simnet_tvar_53[4].label[99] );
tran (\_zy_simnet_tvar_53[4][107] , \_zy_simnet_tvar_53[4].label[98] );
tran (\_zy_simnet_tvar_53[4][106] , \_zy_simnet_tvar_53[4].label[97] );
tran (\_zy_simnet_tvar_53[4][105] , \_zy_simnet_tvar_53[4].label[96] );
tran (\_zy_simnet_tvar_53[4][104] , \_zy_simnet_tvar_53[4].label[95] );
tran (\_zy_simnet_tvar_53[4][103] , \_zy_simnet_tvar_53[4].label[94] );
tran (\_zy_simnet_tvar_53[4][102] , \_zy_simnet_tvar_53[4].label[93] );
tran (\_zy_simnet_tvar_53[4][101] , \_zy_simnet_tvar_53[4].label[92] );
tran (\_zy_simnet_tvar_53[4][100] , \_zy_simnet_tvar_53[4].label[91] );
tran (\_zy_simnet_tvar_53[4][99] , \_zy_simnet_tvar_53[4].label[90] );
tran (\_zy_simnet_tvar_53[4][98] , \_zy_simnet_tvar_53[4].label[89] );
tran (\_zy_simnet_tvar_53[4][97] , \_zy_simnet_tvar_53[4].label[88] );
tran (\_zy_simnet_tvar_53[4][96] , \_zy_simnet_tvar_53[4].label[87] );
tran (\_zy_simnet_tvar_53[4][95] , \_zy_simnet_tvar_53[4].label[86] );
tran (\_zy_simnet_tvar_53[4][94] , \_zy_simnet_tvar_53[4].label[85] );
tran (\_zy_simnet_tvar_53[4][93] , \_zy_simnet_tvar_53[4].label[84] );
tran (\_zy_simnet_tvar_53[4][92] , \_zy_simnet_tvar_53[4].label[83] );
tran (\_zy_simnet_tvar_53[4][91] , \_zy_simnet_tvar_53[4].label[82] );
tran (\_zy_simnet_tvar_53[4][90] , \_zy_simnet_tvar_53[4].label[81] );
tran (\_zy_simnet_tvar_53[4][89] , \_zy_simnet_tvar_53[4].label[80] );
tran (\_zy_simnet_tvar_53[4][88] , \_zy_simnet_tvar_53[4].label[79] );
tran (\_zy_simnet_tvar_53[4][87] , \_zy_simnet_tvar_53[4].label[78] );
tran (\_zy_simnet_tvar_53[4][86] , \_zy_simnet_tvar_53[4].label[77] );
tran (\_zy_simnet_tvar_53[4][85] , \_zy_simnet_tvar_53[4].label[76] );
tran (\_zy_simnet_tvar_53[4][84] , \_zy_simnet_tvar_53[4].label[75] );
tran (\_zy_simnet_tvar_53[4][83] , \_zy_simnet_tvar_53[4].label[74] );
tran (\_zy_simnet_tvar_53[4][82] , \_zy_simnet_tvar_53[4].label[73] );
tran (\_zy_simnet_tvar_53[4][81] , \_zy_simnet_tvar_53[4].label[72] );
tran (\_zy_simnet_tvar_53[4][80] , \_zy_simnet_tvar_53[4].label[71] );
tran (\_zy_simnet_tvar_53[4][79] , \_zy_simnet_tvar_53[4].label[70] );
tran (\_zy_simnet_tvar_53[4][78] , \_zy_simnet_tvar_53[4].label[69] );
tran (\_zy_simnet_tvar_53[4][77] , \_zy_simnet_tvar_53[4].label[68] );
tran (\_zy_simnet_tvar_53[4][76] , \_zy_simnet_tvar_53[4].label[67] );
tran (\_zy_simnet_tvar_53[4][75] , \_zy_simnet_tvar_53[4].label[66] );
tran (\_zy_simnet_tvar_53[4][74] , \_zy_simnet_tvar_53[4].label[65] );
tran (\_zy_simnet_tvar_53[4][73] , \_zy_simnet_tvar_53[4].label[64] );
tran (\_zy_simnet_tvar_53[4][72] , \_zy_simnet_tvar_53[4].label[63] );
tran (\_zy_simnet_tvar_53[4][71] , \_zy_simnet_tvar_53[4].label[62] );
tran (\_zy_simnet_tvar_53[4][70] , \_zy_simnet_tvar_53[4].label[61] );
tran (\_zy_simnet_tvar_53[4][69] , \_zy_simnet_tvar_53[4].label[60] );
tran (\_zy_simnet_tvar_53[4][68] , \_zy_simnet_tvar_53[4].label[59] );
tran (\_zy_simnet_tvar_53[4][67] , \_zy_simnet_tvar_53[4].label[58] );
tran (\_zy_simnet_tvar_53[4][66] , \_zy_simnet_tvar_53[4].label[57] );
tran (\_zy_simnet_tvar_53[4][65] , \_zy_simnet_tvar_53[4].label[56] );
tran (\_zy_simnet_tvar_53[4][64] , \_zy_simnet_tvar_53[4].label[55] );
tran (\_zy_simnet_tvar_53[4][63] , \_zy_simnet_tvar_53[4].label[54] );
tran (\_zy_simnet_tvar_53[4][62] , \_zy_simnet_tvar_53[4].label[53] );
tran (\_zy_simnet_tvar_53[4][61] , \_zy_simnet_tvar_53[4].label[52] );
tran (\_zy_simnet_tvar_53[4][60] , \_zy_simnet_tvar_53[4].label[51] );
tran (\_zy_simnet_tvar_53[4][59] , \_zy_simnet_tvar_53[4].label[50] );
tran (\_zy_simnet_tvar_53[4][58] , \_zy_simnet_tvar_53[4].label[49] );
tran (\_zy_simnet_tvar_53[4][57] , \_zy_simnet_tvar_53[4].label[48] );
tran (\_zy_simnet_tvar_53[4][56] , \_zy_simnet_tvar_53[4].label[47] );
tran (\_zy_simnet_tvar_53[4][55] , \_zy_simnet_tvar_53[4].label[46] );
tran (\_zy_simnet_tvar_53[4][54] , \_zy_simnet_tvar_53[4].label[45] );
tran (\_zy_simnet_tvar_53[4][53] , \_zy_simnet_tvar_53[4].label[44] );
tran (\_zy_simnet_tvar_53[4][52] , \_zy_simnet_tvar_53[4].label[43] );
tran (\_zy_simnet_tvar_53[4][51] , \_zy_simnet_tvar_53[4].label[42] );
tran (\_zy_simnet_tvar_53[4][50] , \_zy_simnet_tvar_53[4].label[41] );
tran (\_zy_simnet_tvar_53[4][49] , \_zy_simnet_tvar_53[4].label[40] );
tran (\_zy_simnet_tvar_53[4][48] , \_zy_simnet_tvar_53[4].label[39] );
tran (\_zy_simnet_tvar_53[4][47] , \_zy_simnet_tvar_53[4].label[38] );
tran (\_zy_simnet_tvar_53[4][46] , \_zy_simnet_tvar_53[4].label[37] );
tran (\_zy_simnet_tvar_53[4][45] , \_zy_simnet_tvar_53[4].label[36] );
tran (\_zy_simnet_tvar_53[4][44] , \_zy_simnet_tvar_53[4].label[35] );
tran (\_zy_simnet_tvar_53[4][43] , \_zy_simnet_tvar_53[4].label[34] );
tran (\_zy_simnet_tvar_53[4][42] , \_zy_simnet_tvar_53[4].label[33] );
tran (\_zy_simnet_tvar_53[4][41] , \_zy_simnet_tvar_53[4].label[32] );
tran (\_zy_simnet_tvar_53[4][40] , \_zy_simnet_tvar_53[4].label[31] );
tran (\_zy_simnet_tvar_53[4][39] , \_zy_simnet_tvar_53[4].label[30] );
tran (\_zy_simnet_tvar_53[4][38] , \_zy_simnet_tvar_53[4].label[29] );
tran (\_zy_simnet_tvar_53[4][37] , \_zy_simnet_tvar_53[4].label[28] );
tran (\_zy_simnet_tvar_53[4][36] , \_zy_simnet_tvar_53[4].label[27] );
tran (\_zy_simnet_tvar_53[4][35] , \_zy_simnet_tvar_53[4].label[26] );
tran (\_zy_simnet_tvar_53[4][34] , \_zy_simnet_tvar_53[4].label[25] );
tran (\_zy_simnet_tvar_53[4][33] , \_zy_simnet_tvar_53[4].label[24] );
tran (\_zy_simnet_tvar_53[4][32] , \_zy_simnet_tvar_53[4].label[23] );
tran (\_zy_simnet_tvar_53[4][31] , \_zy_simnet_tvar_53[4].label[22] );
tran (\_zy_simnet_tvar_53[4][30] , \_zy_simnet_tvar_53[4].label[21] );
tran (\_zy_simnet_tvar_53[4][29] , \_zy_simnet_tvar_53[4].label[20] );
tran (\_zy_simnet_tvar_53[4][28] , \_zy_simnet_tvar_53[4].label[19] );
tran (\_zy_simnet_tvar_53[4][27] , \_zy_simnet_tvar_53[4].label[18] );
tran (\_zy_simnet_tvar_53[4][26] , \_zy_simnet_tvar_53[4].label[17] );
tran (\_zy_simnet_tvar_53[4][25] , \_zy_simnet_tvar_53[4].label[16] );
tran (\_zy_simnet_tvar_53[4][24] , \_zy_simnet_tvar_53[4].label[15] );
tran (\_zy_simnet_tvar_53[4][23] , \_zy_simnet_tvar_53[4].label[14] );
tran (\_zy_simnet_tvar_53[4][22] , \_zy_simnet_tvar_53[4].label[13] );
tran (\_zy_simnet_tvar_53[4][21] , \_zy_simnet_tvar_53[4].label[12] );
tran (\_zy_simnet_tvar_53[4][20] , \_zy_simnet_tvar_53[4].label[11] );
tran (\_zy_simnet_tvar_53[4][19] , \_zy_simnet_tvar_53[4].label[10] );
tran (\_zy_simnet_tvar_53[4][18] , \_zy_simnet_tvar_53[4].label[9] );
tran (\_zy_simnet_tvar_53[4][17] , \_zy_simnet_tvar_53[4].label[8] );
tran (\_zy_simnet_tvar_53[4][16] , \_zy_simnet_tvar_53[4].label[7] );
tran (\_zy_simnet_tvar_53[4][15] , \_zy_simnet_tvar_53[4].label[6] );
tran (\_zy_simnet_tvar_53[4][14] , \_zy_simnet_tvar_53[4].label[5] );
tran (\_zy_simnet_tvar_53[4][13] , \_zy_simnet_tvar_53[4].label[4] );
tran (\_zy_simnet_tvar_53[4][12] , \_zy_simnet_tvar_53[4].label[3] );
tran (\_zy_simnet_tvar_53[4][11] , \_zy_simnet_tvar_53[4].label[2] );
tran (\_zy_simnet_tvar_53[4][10] , \_zy_simnet_tvar_53[4].label[1] );
tran (\_zy_simnet_tvar_53[4][9] , \_zy_simnet_tvar_53[4].label[0] );
tran (\_zy_simnet_tvar_53[4][8] , \_zy_simnet_tvar_53[4].delimiter_valid[0] );
tran (\_zy_simnet_tvar_53[4][7] , \_zy_simnet_tvar_53[4].delimiter[7] );
tran (\_zy_simnet_tvar_53[4][6] , \_zy_simnet_tvar_53[4].delimiter[6] );
tran (\_zy_simnet_tvar_53[4][5] , \_zy_simnet_tvar_53[4].delimiter[5] );
tran (\_zy_simnet_tvar_53[4][4] , \_zy_simnet_tvar_53[4].delimiter[4] );
tran (\_zy_simnet_tvar_53[4][3] , \_zy_simnet_tvar_53[4].delimiter[3] );
tran (\_zy_simnet_tvar_53[4][2] , \_zy_simnet_tvar_53[4].delimiter[2] );
tran (\_zy_simnet_tvar_53[4][1] , \_zy_simnet_tvar_53[4].delimiter[1] );
tran (\_zy_simnet_tvar_53[4][0] , \_zy_simnet_tvar_53[4].delimiter[0] );
tran (\_zy_simnet_tvar_53[3][271] , \_zy_simnet_tvar_53[3].guid_size[0] );
tran (\_zy_simnet_tvar_53[3][270] , \_zy_simnet_tvar_53[3].label_size[5] );
tran (\_zy_simnet_tvar_53[3][269] , \_zy_simnet_tvar_53[3].label_size[4] );
tran (\_zy_simnet_tvar_53[3][268] , \_zy_simnet_tvar_53[3].label_size[3] );
tran (\_zy_simnet_tvar_53[3][267] , \_zy_simnet_tvar_53[3].label_size[2] );
tran (\_zy_simnet_tvar_53[3][266] , \_zy_simnet_tvar_53[3].label_size[1] );
tran (\_zy_simnet_tvar_53[3][265] , \_zy_simnet_tvar_53[3].label_size[0] );
tran (\_zy_simnet_tvar_53[3][264] , \_zy_simnet_tvar_53[3].label[255] );
tran (\_zy_simnet_tvar_53[3][263] , \_zy_simnet_tvar_53[3].label[254] );
tran (\_zy_simnet_tvar_53[3][262] , \_zy_simnet_tvar_53[3].label[253] );
tran (\_zy_simnet_tvar_53[3][261] , \_zy_simnet_tvar_53[3].label[252] );
tran (\_zy_simnet_tvar_53[3][260] , \_zy_simnet_tvar_53[3].label[251] );
tran (\_zy_simnet_tvar_53[3][259] , \_zy_simnet_tvar_53[3].label[250] );
tran (\_zy_simnet_tvar_53[3][258] , \_zy_simnet_tvar_53[3].label[249] );
tran (\_zy_simnet_tvar_53[3][257] , \_zy_simnet_tvar_53[3].label[248] );
tran (\_zy_simnet_tvar_53[3][256] , \_zy_simnet_tvar_53[3].label[247] );
tran (\_zy_simnet_tvar_53[3][255] , \_zy_simnet_tvar_53[3].label[246] );
tran (\_zy_simnet_tvar_53[3][254] , \_zy_simnet_tvar_53[3].label[245] );
tran (\_zy_simnet_tvar_53[3][253] , \_zy_simnet_tvar_53[3].label[244] );
tran (\_zy_simnet_tvar_53[3][252] , \_zy_simnet_tvar_53[3].label[243] );
tran (\_zy_simnet_tvar_53[3][251] , \_zy_simnet_tvar_53[3].label[242] );
tran (\_zy_simnet_tvar_53[3][250] , \_zy_simnet_tvar_53[3].label[241] );
tran (\_zy_simnet_tvar_53[3][249] , \_zy_simnet_tvar_53[3].label[240] );
tran (\_zy_simnet_tvar_53[3][248] , \_zy_simnet_tvar_53[3].label[239] );
tran (\_zy_simnet_tvar_53[3][247] , \_zy_simnet_tvar_53[3].label[238] );
tran (\_zy_simnet_tvar_53[3][246] , \_zy_simnet_tvar_53[3].label[237] );
tran (\_zy_simnet_tvar_53[3][245] , \_zy_simnet_tvar_53[3].label[236] );
tran (\_zy_simnet_tvar_53[3][244] , \_zy_simnet_tvar_53[3].label[235] );
tran (\_zy_simnet_tvar_53[3][243] , \_zy_simnet_tvar_53[3].label[234] );
tran (\_zy_simnet_tvar_53[3][242] , \_zy_simnet_tvar_53[3].label[233] );
tran (\_zy_simnet_tvar_53[3][241] , \_zy_simnet_tvar_53[3].label[232] );
tran (\_zy_simnet_tvar_53[3][240] , \_zy_simnet_tvar_53[3].label[231] );
tran (\_zy_simnet_tvar_53[3][239] , \_zy_simnet_tvar_53[3].label[230] );
tran (\_zy_simnet_tvar_53[3][238] , \_zy_simnet_tvar_53[3].label[229] );
tran (\_zy_simnet_tvar_53[3][237] , \_zy_simnet_tvar_53[3].label[228] );
tran (\_zy_simnet_tvar_53[3][236] , \_zy_simnet_tvar_53[3].label[227] );
tran (\_zy_simnet_tvar_53[3][235] , \_zy_simnet_tvar_53[3].label[226] );
tran (\_zy_simnet_tvar_53[3][234] , \_zy_simnet_tvar_53[3].label[225] );
tran (\_zy_simnet_tvar_53[3][233] , \_zy_simnet_tvar_53[3].label[224] );
tran (\_zy_simnet_tvar_53[3][232] , \_zy_simnet_tvar_53[3].label[223] );
tran (\_zy_simnet_tvar_53[3][231] , \_zy_simnet_tvar_53[3].label[222] );
tran (\_zy_simnet_tvar_53[3][230] , \_zy_simnet_tvar_53[3].label[221] );
tran (\_zy_simnet_tvar_53[3][229] , \_zy_simnet_tvar_53[3].label[220] );
tran (\_zy_simnet_tvar_53[3][228] , \_zy_simnet_tvar_53[3].label[219] );
tran (\_zy_simnet_tvar_53[3][227] , \_zy_simnet_tvar_53[3].label[218] );
tran (\_zy_simnet_tvar_53[3][226] , \_zy_simnet_tvar_53[3].label[217] );
tran (\_zy_simnet_tvar_53[3][225] , \_zy_simnet_tvar_53[3].label[216] );
tran (\_zy_simnet_tvar_53[3][224] , \_zy_simnet_tvar_53[3].label[215] );
tran (\_zy_simnet_tvar_53[3][223] , \_zy_simnet_tvar_53[3].label[214] );
tran (\_zy_simnet_tvar_53[3][222] , \_zy_simnet_tvar_53[3].label[213] );
tran (\_zy_simnet_tvar_53[3][221] , \_zy_simnet_tvar_53[3].label[212] );
tran (\_zy_simnet_tvar_53[3][220] , \_zy_simnet_tvar_53[3].label[211] );
tran (\_zy_simnet_tvar_53[3][219] , \_zy_simnet_tvar_53[3].label[210] );
tran (\_zy_simnet_tvar_53[3][218] , \_zy_simnet_tvar_53[3].label[209] );
tran (\_zy_simnet_tvar_53[3][217] , \_zy_simnet_tvar_53[3].label[208] );
tran (\_zy_simnet_tvar_53[3][216] , \_zy_simnet_tvar_53[3].label[207] );
tran (\_zy_simnet_tvar_53[3][215] , \_zy_simnet_tvar_53[3].label[206] );
tran (\_zy_simnet_tvar_53[3][214] , \_zy_simnet_tvar_53[3].label[205] );
tran (\_zy_simnet_tvar_53[3][213] , \_zy_simnet_tvar_53[3].label[204] );
tran (\_zy_simnet_tvar_53[3][212] , \_zy_simnet_tvar_53[3].label[203] );
tran (\_zy_simnet_tvar_53[3][211] , \_zy_simnet_tvar_53[3].label[202] );
tran (\_zy_simnet_tvar_53[3][210] , \_zy_simnet_tvar_53[3].label[201] );
tran (\_zy_simnet_tvar_53[3][209] , \_zy_simnet_tvar_53[3].label[200] );
tran (\_zy_simnet_tvar_53[3][208] , \_zy_simnet_tvar_53[3].label[199] );
tran (\_zy_simnet_tvar_53[3][207] , \_zy_simnet_tvar_53[3].label[198] );
tran (\_zy_simnet_tvar_53[3][206] , \_zy_simnet_tvar_53[3].label[197] );
tran (\_zy_simnet_tvar_53[3][205] , \_zy_simnet_tvar_53[3].label[196] );
tran (\_zy_simnet_tvar_53[3][204] , \_zy_simnet_tvar_53[3].label[195] );
tran (\_zy_simnet_tvar_53[3][203] , \_zy_simnet_tvar_53[3].label[194] );
tran (\_zy_simnet_tvar_53[3][202] , \_zy_simnet_tvar_53[3].label[193] );
tran (\_zy_simnet_tvar_53[3][201] , \_zy_simnet_tvar_53[3].label[192] );
tran (\_zy_simnet_tvar_53[3][200] , \_zy_simnet_tvar_53[3].label[191] );
tran (\_zy_simnet_tvar_53[3][199] , \_zy_simnet_tvar_53[3].label[190] );
tran (\_zy_simnet_tvar_53[3][198] , \_zy_simnet_tvar_53[3].label[189] );
tran (\_zy_simnet_tvar_53[3][197] , \_zy_simnet_tvar_53[3].label[188] );
tran (\_zy_simnet_tvar_53[3][196] , \_zy_simnet_tvar_53[3].label[187] );
tran (\_zy_simnet_tvar_53[3][195] , \_zy_simnet_tvar_53[3].label[186] );
tran (\_zy_simnet_tvar_53[3][194] , \_zy_simnet_tvar_53[3].label[185] );
tran (\_zy_simnet_tvar_53[3][193] , \_zy_simnet_tvar_53[3].label[184] );
tran (\_zy_simnet_tvar_53[3][192] , \_zy_simnet_tvar_53[3].label[183] );
tran (\_zy_simnet_tvar_53[3][191] , \_zy_simnet_tvar_53[3].label[182] );
tran (\_zy_simnet_tvar_53[3][190] , \_zy_simnet_tvar_53[3].label[181] );
tran (\_zy_simnet_tvar_53[3][189] , \_zy_simnet_tvar_53[3].label[180] );
tran (\_zy_simnet_tvar_53[3][188] , \_zy_simnet_tvar_53[3].label[179] );
tran (\_zy_simnet_tvar_53[3][187] , \_zy_simnet_tvar_53[3].label[178] );
tran (\_zy_simnet_tvar_53[3][186] , \_zy_simnet_tvar_53[3].label[177] );
tran (\_zy_simnet_tvar_53[3][185] , \_zy_simnet_tvar_53[3].label[176] );
tran (\_zy_simnet_tvar_53[3][184] , \_zy_simnet_tvar_53[3].label[175] );
tran (\_zy_simnet_tvar_53[3][183] , \_zy_simnet_tvar_53[3].label[174] );
tran (\_zy_simnet_tvar_53[3][182] , \_zy_simnet_tvar_53[3].label[173] );
tran (\_zy_simnet_tvar_53[3][181] , \_zy_simnet_tvar_53[3].label[172] );
tran (\_zy_simnet_tvar_53[3][180] , \_zy_simnet_tvar_53[3].label[171] );
tran (\_zy_simnet_tvar_53[3][179] , \_zy_simnet_tvar_53[3].label[170] );
tran (\_zy_simnet_tvar_53[3][178] , \_zy_simnet_tvar_53[3].label[169] );
tran (\_zy_simnet_tvar_53[3][177] , \_zy_simnet_tvar_53[3].label[168] );
tran (\_zy_simnet_tvar_53[3][176] , \_zy_simnet_tvar_53[3].label[167] );
tran (\_zy_simnet_tvar_53[3][175] , \_zy_simnet_tvar_53[3].label[166] );
tran (\_zy_simnet_tvar_53[3][174] , \_zy_simnet_tvar_53[3].label[165] );
tran (\_zy_simnet_tvar_53[3][173] , \_zy_simnet_tvar_53[3].label[164] );
tran (\_zy_simnet_tvar_53[3][172] , \_zy_simnet_tvar_53[3].label[163] );
tran (\_zy_simnet_tvar_53[3][171] , \_zy_simnet_tvar_53[3].label[162] );
tran (\_zy_simnet_tvar_53[3][170] , \_zy_simnet_tvar_53[3].label[161] );
tran (\_zy_simnet_tvar_53[3][169] , \_zy_simnet_tvar_53[3].label[160] );
tran (\_zy_simnet_tvar_53[3][168] , \_zy_simnet_tvar_53[3].label[159] );
tran (\_zy_simnet_tvar_53[3][167] , \_zy_simnet_tvar_53[3].label[158] );
tran (\_zy_simnet_tvar_53[3][166] , \_zy_simnet_tvar_53[3].label[157] );
tran (\_zy_simnet_tvar_53[3][165] , \_zy_simnet_tvar_53[3].label[156] );
tran (\_zy_simnet_tvar_53[3][164] , \_zy_simnet_tvar_53[3].label[155] );
tran (\_zy_simnet_tvar_53[3][163] , \_zy_simnet_tvar_53[3].label[154] );
tran (\_zy_simnet_tvar_53[3][162] , \_zy_simnet_tvar_53[3].label[153] );
tran (\_zy_simnet_tvar_53[3][161] , \_zy_simnet_tvar_53[3].label[152] );
tran (\_zy_simnet_tvar_53[3][160] , \_zy_simnet_tvar_53[3].label[151] );
tran (\_zy_simnet_tvar_53[3][159] , \_zy_simnet_tvar_53[3].label[150] );
tran (\_zy_simnet_tvar_53[3][158] , \_zy_simnet_tvar_53[3].label[149] );
tran (\_zy_simnet_tvar_53[3][157] , \_zy_simnet_tvar_53[3].label[148] );
tran (\_zy_simnet_tvar_53[3][156] , \_zy_simnet_tvar_53[3].label[147] );
tran (\_zy_simnet_tvar_53[3][155] , \_zy_simnet_tvar_53[3].label[146] );
tran (\_zy_simnet_tvar_53[3][154] , \_zy_simnet_tvar_53[3].label[145] );
tran (\_zy_simnet_tvar_53[3][153] , \_zy_simnet_tvar_53[3].label[144] );
tran (\_zy_simnet_tvar_53[3][152] , \_zy_simnet_tvar_53[3].label[143] );
tran (\_zy_simnet_tvar_53[3][151] , \_zy_simnet_tvar_53[3].label[142] );
tran (\_zy_simnet_tvar_53[3][150] , \_zy_simnet_tvar_53[3].label[141] );
tran (\_zy_simnet_tvar_53[3][149] , \_zy_simnet_tvar_53[3].label[140] );
tran (\_zy_simnet_tvar_53[3][148] , \_zy_simnet_tvar_53[3].label[139] );
tran (\_zy_simnet_tvar_53[3][147] , \_zy_simnet_tvar_53[3].label[138] );
tran (\_zy_simnet_tvar_53[3][146] , \_zy_simnet_tvar_53[3].label[137] );
tran (\_zy_simnet_tvar_53[3][145] , \_zy_simnet_tvar_53[3].label[136] );
tran (\_zy_simnet_tvar_53[3][144] , \_zy_simnet_tvar_53[3].label[135] );
tran (\_zy_simnet_tvar_53[3][143] , \_zy_simnet_tvar_53[3].label[134] );
tran (\_zy_simnet_tvar_53[3][142] , \_zy_simnet_tvar_53[3].label[133] );
tran (\_zy_simnet_tvar_53[3][141] , \_zy_simnet_tvar_53[3].label[132] );
tran (\_zy_simnet_tvar_53[3][140] , \_zy_simnet_tvar_53[3].label[131] );
tran (\_zy_simnet_tvar_53[3][139] , \_zy_simnet_tvar_53[3].label[130] );
tran (\_zy_simnet_tvar_53[3][138] , \_zy_simnet_tvar_53[3].label[129] );
tran (\_zy_simnet_tvar_53[3][137] , \_zy_simnet_tvar_53[3].label[128] );
tran (\_zy_simnet_tvar_53[3][136] , \_zy_simnet_tvar_53[3].label[127] );
tran (\_zy_simnet_tvar_53[3][135] , \_zy_simnet_tvar_53[3].label[126] );
tran (\_zy_simnet_tvar_53[3][134] , \_zy_simnet_tvar_53[3].label[125] );
tran (\_zy_simnet_tvar_53[3][133] , \_zy_simnet_tvar_53[3].label[124] );
tran (\_zy_simnet_tvar_53[3][132] , \_zy_simnet_tvar_53[3].label[123] );
tran (\_zy_simnet_tvar_53[3][131] , \_zy_simnet_tvar_53[3].label[122] );
tran (\_zy_simnet_tvar_53[3][130] , \_zy_simnet_tvar_53[3].label[121] );
tran (\_zy_simnet_tvar_53[3][129] , \_zy_simnet_tvar_53[3].label[120] );
tran (\_zy_simnet_tvar_53[3][128] , \_zy_simnet_tvar_53[3].label[119] );
tran (\_zy_simnet_tvar_53[3][127] , \_zy_simnet_tvar_53[3].label[118] );
tran (\_zy_simnet_tvar_53[3][126] , \_zy_simnet_tvar_53[3].label[117] );
tran (\_zy_simnet_tvar_53[3][125] , \_zy_simnet_tvar_53[3].label[116] );
tran (\_zy_simnet_tvar_53[3][124] , \_zy_simnet_tvar_53[3].label[115] );
tran (\_zy_simnet_tvar_53[3][123] , \_zy_simnet_tvar_53[3].label[114] );
tran (\_zy_simnet_tvar_53[3][122] , \_zy_simnet_tvar_53[3].label[113] );
tran (\_zy_simnet_tvar_53[3][121] , \_zy_simnet_tvar_53[3].label[112] );
tran (\_zy_simnet_tvar_53[3][120] , \_zy_simnet_tvar_53[3].label[111] );
tran (\_zy_simnet_tvar_53[3][119] , \_zy_simnet_tvar_53[3].label[110] );
tran (\_zy_simnet_tvar_53[3][118] , \_zy_simnet_tvar_53[3].label[109] );
tran (\_zy_simnet_tvar_53[3][117] , \_zy_simnet_tvar_53[3].label[108] );
tran (\_zy_simnet_tvar_53[3][116] , \_zy_simnet_tvar_53[3].label[107] );
tran (\_zy_simnet_tvar_53[3][115] , \_zy_simnet_tvar_53[3].label[106] );
tran (\_zy_simnet_tvar_53[3][114] , \_zy_simnet_tvar_53[3].label[105] );
tran (\_zy_simnet_tvar_53[3][113] , \_zy_simnet_tvar_53[3].label[104] );
tran (\_zy_simnet_tvar_53[3][112] , \_zy_simnet_tvar_53[3].label[103] );
tran (\_zy_simnet_tvar_53[3][111] , \_zy_simnet_tvar_53[3].label[102] );
tran (\_zy_simnet_tvar_53[3][110] , \_zy_simnet_tvar_53[3].label[101] );
tran (\_zy_simnet_tvar_53[3][109] , \_zy_simnet_tvar_53[3].label[100] );
tran (\_zy_simnet_tvar_53[3][108] , \_zy_simnet_tvar_53[3].label[99] );
tran (\_zy_simnet_tvar_53[3][107] , \_zy_simnet_tvar_53[3].label[98] );
tran (\_zy_simnet_tvar_53[3][106] , \_zy_simnet_tvar_53[3].label[97] );
tran (\_zy_simnet_tvar_53[3][105] , \_zy_simnet_tvar_53[3].label[96] );
tran (\_zy_simnet_tvar_53[3][104] , \_zy_simnet_tvar_53[3].label[95] );
tran (\_zy_simnet_tvar_53[3][103] , \_zy_simnet_tvar_53[3].label[94] );
tran (\_zy_simnet_tvar_53[3][102] , \_zy_simnet_tvar_53[3].label[93] );
tran (\_zy_simnet_tvar_53[3][101] , \_zy_simnet_tvar_53[3].label[92] );
tran (\_zy_simnet_tvar_53[3][100] , \_zy_simnet_tvar_53[3].label[91] );
tran (\_zy_simnet_tvar_53[3][99] , \_zy_simnet_tvar_53[3].label[90] );
tran (\_zy_simnet_tvar_53[3][98] , \_zy_simnet_tvar_53[3].label[89] );
tran (\_zy_simnet_tvar_53[3][97] , \_zy_simnet_tvar_53[3].label[88] );
tran (\_zy_simnet_tvar_53[3][96] , \_zy_simnet_tvar_53[3].label[87] );
tran (\_zy_simnet_tvar_53[3][95] , \_zy_simnet_tvar_53[3].label[86] );
tran (\_zy_simnet_tvar_53[3][94] , \_zy_simnet_tvar_53[3].label[85] );
tran (\_zy_simnet_tvar_53[3][93] , \_zy_simnet_tvar_53[3].label[84] );
tran (\_zy_simnet_tvar_53[3][92] , \_zy_simnet_tvar_53[3].label[83] );
tran (\_zy_simnet_tvar_53[3][91] , \_zy_simnet_tvar_53[3].label[82] );
tran (\_zy_simnet_tvar_53[3][90] , \_zy_simnet_tvar_53[3].label[81] );
tran (\_zy_simnet_tvar_53[3][89] , \_zy_simnet_tvar_53[3].label[80] );
tran (\_zy_simnet_tvar_53[3][88] , \_zy_simnet_tvar_53[3].label[79] );
tran (\_zy_simnet_tvar_53[3][87] , \_zy_simnet_tvar_53[3].label[78] );
tran (\_zy_simnet_tvar_53[3][86] , \_zy_simnet_tvar_53[3].label[77] );
tran (\_zy_simnet_tvar_53[3][85] , \_zy_simnet_tvar_53[3].label[76] );
tran (\_zy_simnet_tvar_53[3][84] , \_zy_simnet_tvar_53[3].label[75] );
tran (\_zy_simnet_tvar_53[3][83] , \_zy_simnet_tvar_53[3].label[74] );
tran (\_zy_simnet_tvar_53[3][82] , \_zy_simnet_tvar_53[3].label[73] );
tran (\_zy_simnet_tvar_53[3][81] , \_zy_simnet_tvar_53[3].label[72] );
tran (\_zy_simnet_tvar_53[3][80] , \_zy_simnet_tvar_53[3].label[71] );
tran (\_zy_simnet_tvar_53[3][79] , \_zy_simnet_tvar_53[3].label[70] );
tran (\_zy_simnet_tvar_53[3][78] , \_zy_simnet_tvar_53[3].label[69] );
tran (\_zy_simnet_tvar_53[3][77] , \_zy_simnet_tvar_53[3].label[68] );
tran (\_zy_simnet_tvar_53[3][76] , \_zy_simnet_tvar_53[3].label[67] );
tran (\_zy_simnet_tvar_53[3][75] , \_zy_simnet_tvar_53[3].label[66] );
tran (\_zy_simnet_tvar_53[3][74] , \_zy_simnet_tvar_53[3].label[65] );
tran (\_zy_simnet_tvar_53[3][73] , \_zy_simnet_tvar_53[3].label[64] );
tran (\_zy_simnet_tvar_53[3][72] , \_zy_simnet_tvar_53[3].label[63] );
tran (\_zy_simnet_tvar_53[3][71] , \_zy_simnet_tvar_53[3].label[62] );
tran (\_zy_simnet_tvar_53[3][70] , \_zy_simnet_tvar_53[3].label[61] );
tran (\_zy_simnet_tvar_53[3][69] , \_zy_simnet_tvar_53[3].label[60] );
tran (\_zy_simnet_tvar_53[3][68] , \_zy_simnet_tvar_53[3].label[59] );
tran (\_zy_simnet_tvar_53[3][67] , \_zy_simnet_tvar_53[3].label[58] );
tran (\_zy_simnet_tvar_53[3][66] , \_zy_simnet_tvar_53[3].label[57] );
tran (\_zy_simnet_tvar_53[3][65] , \_zy_simnet_tvar_53[3].label[56] );
tran (\_zy_simnet_tvar_53[3][64] , \_zy_simnet_tvar_53[3].label[55] );
tran (\_zy_simnet_tvar_53[3][63] , \_zy_simnet_tvar_53[3].label[54] );
tran (\_zy_simnet_tvar_53[3][62] , \_zy_simnet_tvar_53[3].label[53] );
tran (\_zy_simnet_tvar_53[3][61] , \_zy_simnet_tvar_53[3].label[52] );
tran (\_zy_simnet_tvar_53[3][60] , \_zy_simnet_tvar_53[3].label[51] );
tran (\_zy_simnet_tvar_53[3][59] , \_zy_simnet_tvar_53[3].label[50] );
tran (\_zy_simnet_tvar_53[3][58] , \_zy_simnet_tvar_53[3].label[49] );
tran (\_zy_simnet_tvar_53[3][57] , \_zy_simnet_tvar_53[3].label[48] );
tran (\_zy_simnet_tvar_53[3][56] , \_zy_simnet_tvar_53[3].label[47] );
tran (\_zy_simnet_tvar_53[3][55] , \_zy_simnet_tvar_53[3].label[46] );
tran (\_zy_simnet_tvar_53[3][54] , \_zy_simnet_tvar_53[3].label[45] );
tran (\_zy_simnet_tvar_53[3][53] , \_zy_simnet_tvar_53[3].label[44] );
tran (\_zy_simnet_tvar_53[3][52] , \_zy_simnet_tvar_53[3].label[43] );
tran (\_zy_simnet_tvar_53[3][51] , \_zy_simnet_tvar_53[3].label[42] );
tran (\_zy_simnet_tvar_53[3][50] , \_zy_simnet_tvar_53[3].label[41] );
tran (\_zy_simnet_tvar_53[3][49] , \_zy_simnet_tvar_53[3].label[40] );
tran (\_zy_simnet_tvar_53[3][48] , \_zy_simnet_tvar_53[3].label[39] );
tran (\_zy_simnet_tvar_53[3][47] , \_zy_simnet_tvar_53[3].label[38] );
tran (\_zy_simnet_tvar_53[3][46] , \_zy_simnet_tvar_53[3].label[37] );
tran (\_zy_simnet_tvar_53[3][45] , \_zy_simnet_tvar_53[3].label[36] );
tran (\_zy_simnet_tvar_53[3][44] , \_zy_simnet_tvar_53[3].label[35] );
tran (\_zy_simnet_tvar_53[3][43] , \_zy_simnet_tvar_53[3].label[34] );
tran (\_zy_simnet_tvar_53[3][42] , \_zy_simnet_tvar_53[3].label[33] );
tran (\_zy_simnet_tvar_53[3][41] , \_zy_simnet_tvar_53[3].label[32] );
tran (\_zy_simnet_tvar_53[3][40] , \_zy_simnet_tvar_53[3].label[31] );
tran (\_zy_simnet_tvar_53[3][39] , \_zy_simnet_tvar_53[3].label[30] );
tran (\_zy_simnet_tvar_53[3][38] , \_zy_simnet_tvar_53[3].label[29] );
tran (\_zy_simnet_tvar_53[3][37] , \_zy_simnet_tvar_53[3].label[28] );
tran (\_zy_simnet_tvar_53[3][36] , \_zy_simnet_tvar_53[3].label[27] );
tran (\_zy_simnet_tvar_53[3][35] , \_zy_simnet_tvar_53[3].label[26] );
tran (\_zy_simnet_tvar_53[3][34] , \_zy_simnet_tvar_53[3].label[25] );
tran (\_zy_simnet_tvar_53[3][33] , \_zy_simnet_tvar_53[3].label[24] );
tran (\_zy_simnet_tvar_53[3][32] , \_zy_simnet_tvar_53[3].label[23] );
tran (\_zy_simnet_tvar_53[3][31] , \_zy_simnet_tvar_53[3].label[22] );
tran (\_zy_simnet_tvar_53[3][30] , \_zy_simnet_tvar_53[3].label[21] );
tran (\_zy_simnet_tvar_53[3][29] , \_zy_simnet_tvar_53[3].label[20] );
tran (\_zy_simnet_tvar_53[3][28] , \_zy_simnet_tvar_53[3].label[19] );
tran (\_zy_simnet_tvar_53[3][27] , \_zy_simnet_tvar_53[3].label[18] );
tran (\_zy_simnet_tvar_53[3][26] , \_zy_simnet_tvar_53[3].label[17] );
tran (\_zy_simnet_tvar_53[3][25] , \_zy_simnet_tvar_53[3].label[16] );
tran (\_zy_simnet_tvar_53[3][24] , \_zy_simnet_tvar_53[3].label[15] );
tran (\_zy_simnet_tvar_53[3][23] , \_zy_simnet_tvar_53[3].label[14] );
tran (\_zy_simnet_tvar_53[3][22] , \_zy_simnet_tvar_53[3].label[13] );
tran (\_zy_simnet_tvar_53[3][21] , \_zy_simnet_tvar_53[3].label[12] );
tran (\_zy_simnet_tvar_53[3][20] , \_zy_simnet_tvar_53[3].label[11] );
tran (\_zy_simnet_tvar_53[3][19] , \_zy_simnet_tvar_53[3].label[10] );
tran (\_zy_simnet_tvar_53[3][18] , \_zy_simnet_tvar_53[3].label[9] );
tran (\_zy_simnet_tvar_53[3][17] , \_zy_simnet_tvar_53[3].label[8] );
tran (\_zy_simnet_tvar_53[3][16] , \_zy_simnet_tvar_53[3].label[7] );
tran (\_zy_simnet_tvar_53[3][15] , \_zy_simnet_tvar_53[3].label[6] );
tran (\_zy_simnet_tvar_53[3][14] , \_zy_simnet_tvar_53[3].label[5] );
tran (\_zy_simnet_tvar_53[3][13] , \_zy_simnet_tvar_53[3].label[4] );
tran (\_zy_simnet_tvar_53[3][12] , \_zy_simnet_tvar_53[3].label[3] );
tran (\_zy_simnet_tvar_53[3][11] , \_zy_simnet_tvar_53[3].label[2] );
tran (\_zy_simnet_tvar_53[3][10] , \_zy_simnet_tvar_53[3].label[1] );
tran (\_zy_simnet_tvar_53[3][9] , \_zy_simnet_tvar_53[3].label[0] );
tran (\_zy_simnet_tvar_53[3][8] , \_zy_simnet_tvar_53[3].delimiter_valid[0] );
tran (\_zy_simnet_tvar_53[3][7] , \_zy_simnet_tvar_53[3].delimiter[7] );
tran (\_zy_simnet_tvar_53[3][6] , \_zy_simnet_tvar_53[3].delimiter[6] );
tran (\_zy_simnet_tvar_53[3][5] , \_zy_simnet_tvar_53[3].delimiter[5] );
tran (\_zy_simnet_tvar_53[3][4] , \_zy_simnet_tvar_53[3].delimiter[4] );
tran (\_zy_simnet_tvar_53[3][3] , \_zy_simnet_tvar_53[3].delimiter[3] );
tran (\_zy_simnet_tvar_53[3][2] , \_zy_simnet_tvar_53[3].delimiter[2] );
tran (\_zy_simnet_tvar_53[3][1] , \_zy_simnet_tvar_53[3].delimiter[1] );
tran (\_zy_simnet_tvar_53[3][0] , \_zy_simnet_tvar_53[3].delimiter[0] );
tran (\_zy_simnet_tvar_53[2][271] , \_zy_simnet_tvar_53[2].guid_size[0] );
tran (\_zy_simnet_tvar_53[2][270] , \_zy_simnet_tvar_53[2].label_size[5] );
tran (\_zy_simnet_tvar_53[2][269] , \_zy_simnet_tvar_53[2].label_size[4] );
tran (\_zy_simnet_tvar_53[2][268] , \_zy_simnet_tvar_53[2].label_size[3] );
tran (\_zy_simnet_tvar_53[2][267] , \_zy_simnet_tvar_53[2].label_size[2] );
tran (\_zy_simnet_tvar_53[2][266] , \_zy_simnet_tvar_53[2].label_size[1] );
tran (\_zy_simnet_tvar_53[2][265] , \_zy_simnet_tvar_53[2].label_size[0] );
tran (\_zy_simnet_tvar_53[2][264] , \_zy_simnet_tvar_53[2].label[255] );
tran (\_zy_simnet_tvar_53[2][263] , \_zy_simnet_tvar_53[2].label[254] );
tran (\_zy_simnet_tvar_53[2][262] , \_zy_simnet_tvar_53[2].label[253] );
tran (\_zy_simnet_tvar_53[2][261] , \_zy_simnet_tvar_53[2].label[252] );
tran (\_zy_simnet_tvar_53[2][260] , \_zy_simnet_tvar_53[2].label[251] );
tran (\_zy_simnet_tvar_53[2][259] , \_zy_simnet_tvar_53[2].label[250] );
tran (\_zy_simnet_tvar_53[2][258] , \_zy_simnet_tvar_53[2].label[249] );
tran (\_zy_simnet_tvar_53[2][257] , \_zy_simnet_tvar_53[2].label[248] );
tran (\_zy_simnet_tvar_53[2][256] , \_zy_simnet_tvar_53[2].label[247] );
tran (\_zy_simnet_tvar_53[2][255] , \_zy_simnet_tvar_53[2].label[246] );
tran (\_zy_simnet_tvar_53[2][254] , \_zy_simnet_tvar_53[2].label[245] );
tran (\_zy_simnet_tvar_53[2][253] , \_zy_simnet_tvar_53[2].label[244] );
tran (\_zy_simnet_tvar_53[2][252] , \_zy_simnet_tvar_53[2].label[243] );
tran (\_zy_simnet_tvar_53[2][251] , \_zy_simnet_tvar_53[2].label[242] );
tran (\_zy_simnet_tvar_53[2][250] , \_zy_simnet_tvar_53[2].label[241] );
tran (\_zy_simnet_tvar_53[2][249] , \_zy_simnet_tvar_53[2].label[240] );
tran (\_zy_simnet_tvar_53[2][248] , \_zy_simnet_tvar_53[2].label[239] );
tran (\_zy_simnet_tvar_53[2][247] , \_zy_simnet_tvar_53[2].label[238] );
tran (\_zy_simnet_tvar_53[2][246] , \_zy_simnet_tvar_53[2].label[237] );
tran (\_zy_simnet_tvar_53[2][245] , \_zy_simnet_tvar_53[2].label[236] );
tran (\_zy_simnet_tvar_53[2][244] , \_zy_simnet_tvar_53[2].label[235] );
tran (\_zy_simnet_tvar_53[2][243] , \_zy_simnet_tvar_53[2].label[234] );
tran (\_zy_simnet_tvar_53[2][242] , \_zy_simnet_tvar_53[2].label[233] );
tran (\_zy_simnet_tvar_53[2][241] , \_zy_simnet_tvar_53[2].label[232] );
tran (\_zy_simnet_tvar_53[2][240] , \_zy_simnet_tvar_53[2].label[231] );
tran (\_zy_simnet_tvar_53[2][239] , \_zy_simnet_tvar_53[2].label[230] );
tran (\_zy_simnet_tvar_53[2][238] , \_zy_simnet_tvar_53[2].label[229] );
tran (\_zy_simnet_tvar_53[2][237] , \_zy_simnet_tvar_53[2].label[228] );
tran (\_zy_simnet_tvar_53[2][236] , \_zy_simnet_tvar_53[2].label[227] );
tran (\_zy_simnet_tvar_53[2][235] , \_zy_simnet_tvar_53[2].label[226] );
tran (\_zy_simnet_tvar_53[2][234] , \_zy_simnet_tvar_53[2].label[225] );
tran (\_zy_simnet_tvar_53[2][233] , \_zy_simnet_tvar_53[2].label[224] );
tran (\_zy_simnet_tvar_53[2][232] , \_zy_simnet_tvar_53[2].label[223] );
tran (\_zy_simnet_tvar_53[2][231] , \_zy_simnet_tvar_53[2].label[222] );
tran (\_zy_simnet_tvar_53[2][230] , \_zy_simnet_tvar_53[2].label[221] );
tran (\_zy_simnet_tvar_53[2][229] , \_zy_simnet_tvar_53[2].label[220] );
tran (\_zy_simnet_tvar_53[2][228] , \_zy_simnet_tvar_53[2].label[219] );
tran (\_zy_simnet_tvar_53[2][227] , \_zy_simnet_tvar_53[2].label[218] );
tran (\_zy_simnet_tvar_53[2][226] , \_zy_simnet_tvar_53[2].label[217] );
tran (\_zy_simnet_tvar_53[2][225] , \_zy_simnet_tvar_53[2].label[216] );
tran (\_zy_simnet_tvar_53[2][224] , \_zy_simnet_tvar_53[2].label[215] );
tran (\_zy_simnet_tvar_53[2][223] , \_zy_simnet_tvar_53[2].label[214] );
tran (\_zy_simnet_tvar_53[2][222] , \_zy_simnet_tvar_53[2].label[213] );
tran (\_zy_simnet_tvar_53[2][221] , \_zy_simnet_tvar_53[2].label[212] );
tran (\_zy_simnet_tvar_53[2][220] , \_zy_simnet_tvar_53[2].label[211] );
tran (\_zy_simnet_tvar_53[2][219] , \_zy_simnet_tvar_53[2].label[210] );
tran (\_zy_simnet_tvar_53[2][218] , \_zy_simnet_tvar_53[2].label[209] );
tran (\_zy_simnet_tvar_53[2][217] , \_zy_simnet_tvar_53[2].label[208] );
tran (\_zy_simnet_tvar_53[2][216] , \_zy_simnet_tvar_53[2].label[207] );
tran (\_zy_simnet_tvar_53[2][215] , \_zy_simnet_tvar_53[2].label[206] );
tran (\_zy_simnet_tvar_53[2][214] , \_zy_simnet_tvar_53[2].label[205] );
tran (\_zy_simnet_tvar_53[2][213] , \_zy_simnet_tvar_53[2].label[204] );
tran (\_zy_simnet_tvar_53[2][212] , \_zy_simnet_tvar_53[2].label[203] );
tran (\_zy_simnet_tvar_53[2][211] , \_zy_simnet_tvar_53[2].label[202] );
tran (\_zy_simnet_tvar_53[2][210] , \_zy_simnet_tvar_53[2].label[201] );
tran (\_zy_simnet_tvar_53[2][209] , \_zy_simnet_tvar_53[2].label[200] );
tran (\_zy_simnet_tvar_53[2][208] , \_zy_simnet_tvar_53[2].label[199] );
tran (\_zy_simnet_tvar_53[2][207] , \_zy_simnet_tvar_53[2].label[198] );
tran (\_zy_simnet_tvar_53[2][206] , \_zy_simnet_tvar_53[2].label[197] );
tran (\_zy_simnet_tvar_53[2][205] , \_zy_simnet_tvar_53[2].label[196] );
tran (\_zy_simnet_tvar_53[2][204] , \_zy_simnet_tvar_53[2].label[195] );
tran (\_zy_simnet_tvar_53[2][203] , \_zy_simnet_tvar_53[2].label[194] );
tran (\_zy_simnet_tvar_53[2][202] , \_zy_simnet_tvar_53[2].label[193] );
tran (\_zy_simnet_tvar_53[2][201] , \_zy_simnet_tvar_53[2].label[192] );
tran (\_zy_simnet_tvar_53[2][200] , \_zy_simnet_tvar_53[2].label[191] );
tran (\_zy_simnet_tvar_53[2][199] , \_zy_simnet_tvar_53[2].label[190] );
tran (\_zy_simnet_tvar_53[2][198] , \_zy_simnet_tvar_53[2].label[189] );
tran (\_zy_simnet_tvar_53[2][197] , \_zy_simnet_tvar_53[2].label[188] );
tran (\_zy_simnet_tvar_53[2][196] , \_zy_simnet_tvar_53[2].label[187] );
tran (\_zy_simnet_tvar_53[2][195] , \_zy_simnet_tvar_53[2].label[186] );
tran (\_zy_simnet_tvar_53[2][194] , \_zy_simnet_tvar_53[2].label[185] );
tran (\_zy_simnet_tvar_53[2][193] , \_zy_simnet_tvar_53[2].label[184] );
tran (\_zy_simnet_tvar_53[2][192] , \_zy_simnet_tvar_53[2].label[183] );
tran (\_zy_simnet_tvar_53[2][191] , \_zy_simnet_tvar_53[2].label[182] );
tran (\_zy_simnet_tvar_53[2][190] , \_zy_simnet_tvar_53[2].label[181] );
tran (\_zy_simnet_tvar_53[2][189] , \_zy_simnet_tvar_53[2].label[180] );
tran (\_zy_simnet_tvar_53[2][188] , \_zy_simnet_tvar_53[2].label[179] );
tran (\_zy_simnet_tvar_53[2][187] , \_zy_simnet_tvar_53[2].label[178] );
tran (\_zy_simnet_tvar_53[2][186] , \_zy_simnet_tvar_53[2].label[177] );
tran (\_zy_simnet_tvar_53[2][185] , \_zy_simnet_tvar_53[2].label[176] );
tran (\_zy_simnet_tvar_53[2][184] , \_zy_simnet_tvar_53[2].label[175] );
tran (\_zy_simnet_tvar_53[2][183] , \_zy_simnet_tvar_53[2].label[174] );
tran (\_zy_simnet_tvar_53[2][182] , \_zy_simnet_tvar_53[2].label[173] );
tran (\_zy_simnet_tvar_53[2][181] , \_zy_simnet_tvar_53[2].label[172] );
tran (\_zy_simnet_tvar_53[2][180] , \_zy_simnet_tvar_53[2].label[171] );
tran (\_zy_simnet_tvar_53[2][179] , \_zy_simnet_tvar_53[2].label[170] );
tran (\_zy_simnet_tvar_53[2][178] , \_zy_simnet_tvar_53[2].label[169] );
tran (\_zy_simnet_tvar_53[2][177] , \_zy_simnet_tvar_53[2].label[168] );
tran (\_zy_simnet_tvar_53[2][176] , \_zy_simnet_tvar_53[2].label[167] );
tran (\_zy_simnet_tvar_53[2][175] , \_zy_simnet_tvar_53[2].label[166] );
tran (\_zy_simnet_tvar_53[2][174] , \_zy_simnet_tvar_53[2].label[165] );
tran (\_zy_simnet_tvar_53[2][173] , \_zy_simnet_tvar_53[2].label[164] );
tran (\_zy_simnet_tvar_53[2][172] , \_zy_simnet_tvar_53[2].label[163] );
tran (\_zy_simnet_tvar_53[2][171] , \_zy_simnet_tvar_53[2].label[162] );
tran (\_zy_simnet_tvar_53[2][170] , \_zy_simnet_tvar_53[2].label[161] );
tran (\_zy_simnet_tvar_53[2][169] , \_zy_simnet_tvar_53[2].label[160] );
tran (\_zy_simnet_tvar_53[2][168] , \_zy_simnet_tvar_53[2].label[159] );
tran (\_zy_simnet_tvar_53[2][167] , \_zy_simnet_tvar_53[2].label[158] );
tran (\_zy_simnet_tvar_53[2][166] , \_zy_simnet_tvar_53[2].label[157] );
tran (\_zy_simnet_tvar_53[2][165] , \_zy_simnet_tvar_53[2].label[156] );
tran (\_zy_simnet_tvar_53[2][164] , \_zy_simnet_tvar_53[2].label[155] );
tran (\_zy_simnet_tvar_53[2][163] , \_zy_simnet_tvar_53[2].label[154] );
tran (\_zy_simnet_tvar_53[2][162] , \_zy_simnet_tvar_53[2].label[153] );
tran (\_zy_simnet_tvar_53[2][161] , \_zy_simnet_tvar_53[2].label[152] );
tran (\_zy_simnet_tvar_53[2][160] , \_zy_simnet_tvar_53[2].label[151] );
tran (\_zy_simnet_tvar_53[2][159] , \_zy_simnet_tvar_53[2].label[150] );
tran (\_zy_simnet_tvar_53[2][158] , \_zy_simnet_tvar_53[2].label[149] );
tran (\_zy_simnet_tvar_53[2][157] , \_zy_simnet_tvar_53[2].label[148] );
tran (\_zy_simnet_tvar_53[2][156] , \_zy_simnet_tvar_53[2].label[147] );
tran (\_zy_simnet_tvar_53[2][155] , \_zy_simnet_tvar_53[2].label[146] );
tran (\_zy_simnet_tvar_53[2][154] , \_zy_simnet_tvar_53[2].label[145] );
tran (\_zy_simnet_tvar_53[2][153] , \_zy_simnet_tvar_53[2].label[144] );
tran (\_zy_simnet_tvar_53[2][152] , \_zy_simnet_tvar_53[2].label[143] );
tran (\_zy_simnet_tvar_53[2][151] , \_zy_simnet_tvar_53[2].label[142] );
tran (\_zy_simnet_tvar_53[2][150] , \_zy_simnet_tvar_53[2].label[141] );
tran (\_zy_simnet_tvar_53[2][149] , \_zy_simnet_tvar_53[2].label[140] );
tran (\_zy_simnet_tvar_53[2][148] , \_zy_simnet_tvar_53[2].label[139] );
tran (\_zy_simnet_tvar_53[2][147] , \_zy_simnet_tvar_53[2].label[138] );
tran (\_zy_simnet_tvar_53[2][146] , \_zy_simnet_tvar_53[2].label[137] );
tran (\_zy_simnet_tvar_53[2][145] , \_zy_simnet_tvar_53[2].label[136] );
tran (\_zy_simnet_tvar_53[2][144] , \_zy_simnet_tvar_53[2].label[135] );
tran (\_zy_simnet_tvar_53[2][143] , \_zy_simnet_tvar_53[2].label[134] );
tran (\_zy_simnet_tvar_53[2][142] , \_zy_simnet_tvar_53[2].label[133] );
tran (\_zy_simnet_tvar_53[2][141] , \_zy_simnet_tvar_53[2].label[132] );
tran (\_zy_simnet_tvar_53[2][140] , \_zy_simnet_tvar_53[2].label[131] );
tran (\_zy_simnet_tvar_53[2][139] , \_zy_simnet_tvar_53[2].label[130] );
tran (\_zy_simnet_tvar_53[2][138] , \_zy_simnet_tvar_53[2].label[129] );
tran (\_zy_simnet_tvar_53[2][137] , \_zy_simnet_tvar_53[2].label[128] );
tran (\_zy_simnet_tvar_53[2][136] , \_zy_simnet_tvar_53[2].label[127] );
tran (\_zy_simnet_tvar_53[2][135] , \_zy_simnet_tvar_53[2].label[126] );
tran (\_zy_simnet_tvar_53[2][134] , \_zy_simnet_tvar_53[2].label[125] );
tran (\_zy_simnet_tvar_53[2][133] , \_zy_simnet_tvar_53[2].label[124] );
tran (\_zy_simnet_tvar_53[2][132] , \_zy_simnet_tvar_53[2].label[123] );
tran (\_zy_simnet_tvar_53[2][131] , \_zy_simnet_tvar_53[2].label[122] );
tran (\_zy_simnet_tvar_53[2][130] , \_zy_simnet_tvar_53[2].label[121] );
tran (\_zy_simnet_tvar_53[2][129] , \_zy_simnet_tvar_53[2].label[120] );
tran (\_zy_simnet_tvar_53[2][128] , \_zy_simnet_tvar_53[2].label[119] );
tran (\_zy_simnet_tvar_53[2][127] , \_zy_simnet_tvar_53[2].label[118] );
tran (\_zy_simnet_tvar_53[2][126] , \_zy_simnet_tvar_53[2].label[117] );
tran (\_zy_simnet_tvar_53[2][125] , \_zy_simnet_tvar_53[2].label[116] );
tran (\_zy_simnet_tvar_53[2][124] , \_zy_simnet_tvar_53[2].label[115] );
tran (\_zy_simnet_tvar_53[2][123] , \_zy_simnet_tvar_53[2].label[114] );
tran (\_zy_simnet_tvar_53[2][122] , \_zy_simnet_tvar_53[2].label[113] );
tran (\_zy_simnet_tvar_53[2][121] , \_zy_simnet_tvar_53[2].label[112] );
tran (\_zy_simnet_tvar_53[2][120] , \_zy_simnet_tvar_53[2].label[111] );
tran (\_zy_simnet_tvar_53[2][119] , \_zy_simnet_tvar_53[2].label[110] );
tran (\_zy_simnet_tvar_53[2][118] , \_zy_simnet_tvar_53[2].label[109] );
tran (\_zy_simnet_tvar_53[2][117] , \_zy_simnet_tvar_53[2].label[108] );
tran (\_zy_simnet_tvar_53[2][116] , \_zy_simnet_tvar_53[2].label[107] );
tran (\_zy_simnet_tvar_53[2][115] , \_zy_simnet_tvar_53[2].label[106] );
tran (\_zy_simnet_tvar_53[2][114] , \_zy_simnet_tvar_53[2].label[105] );
tran (\_zy_simnet_tvar_53[2][113] , \_zy_simnet_tvar_53[2].label[104] );
tran (\_zy_simnet_tvar_53[2][112] , \_zy_simnet_tvar_53[2].label[103] );
tran (\_zy_simnet_tvar_53[2][111] , \_zy_simnet_tvar_53[2].label[102] );
tran (\_zy_simnet_tvar_53[2][110] , \_zy_simnet_tvar_53[2].label[101] );
tran (\_zy_simnet_tvar_53[2][109] , \_zy_simnet_tvar_53[2].label[100] );
tran (\_zy_simnet_tvar_53[2][108] , \_zy_simnet_tvar_53[2].label[99] );
tran (\_zy_simnet_tvar_53[2][107] , \_zy_simnet_tvar_53[2].label[98] );
tran (\_zy_simnet_tvar_53[2][106] , \_zy_simnet_tvar_53[2].label[97] );
tran (\_zy_simnet_tvar_53[2][105] , \_zy_simnet_tvar_53[2].label[96] );
tran (\_zy_simnet_tvar_53[2][104] , \_zy_simnet_tvar_53[2].label[95] );
tran (\_zy_simnet_tvar_53[2][103] , \_zy_simnet_tvar_53[2].label[94] );
tran (\_zy_simnet_tvar_53[2][102] , \_zy_simnet_tvar_53[2].label[93] );
tran (\_zy_simnet_tvar_53[2][101] , \_zy_simnet_tvar_53[2].label[92] );
tran (\_zy_simnet_tvar_53[2][100] , \_zy_simnet_tvar_53[2].label[91] );
tran (\_zy_simnet_tvar_53[2][99] , \_zy_simnet_tvar_53[2].label[90] );
tran (\_zy_simnet_tvar_53[2][98] , \_zy_simnet_tvar_53[2].label[89] );
tran (\_zy_simnet_tvar_53[2][97] , \_zy_simnet_tvar_53[2].label[88] );
tran (\_zy_simnet_tvar_53[2][96] , \_zy_simnet_tvar_53[2].label[87] );
tran (\_zy_simnet_tvar_53[2][95] , \_zy_simnet_tvar_53[2].label[86] );
tran (\_zy_simnet_tvar_53[2][94] , \_zy_simnet_tvar_53[2].label[85] );
tran (\_zy_simnet_tvar_53[2][93] , \_zy_simnet_tvar_53[2].label[84] );
tran (\_zy_simnet_tvar_53[2][92] , \_zy_simnet_tvar_53[2].label[83] );
tran (\_zy_simnet_tvar_53[2][91] , \_zy_simnet_tvar_53[2].label[82] );
tran (\_zy_simnet_tvar_53[2][90] , \_zy_simnet_tvar_53[2].label[81] );
tran (\_zy_simnet_tvar_53[2][89] , \_zy_simnet_tvar_53[2].label[80] );
tran (\_zy_simnet_tvar_53[2][88] , \_zy_simnet_tvar_53[2].label[79] );
tran (\_zy_simnet_tvar_53[2][87] , \_zy_simnet_tvar_53[2].label[78] );
tran (\_zy_simnet_tvar_53[2][86] , \_zy_simnet_tvar_53[2].label[77] );
tran (\_zy_simnet_tvar_53[2][85] , \_zy_simnet_tvar_53[2].label[76] );
tran (\_zy_simnet_tvar_53[2][84] , \_zy_simnet_tvar_53[2].label[75] );
tran (\_zy_simnet_tvar_53[2][83] , \_zy_simnet_tvar_53[2].label[74] );
tran (\_zy_simnet_tvar_53[2][82] , \_zy_simnet_tvar_53[2].label[73] );
tran (\_zy_simnet_tvar_53[2][81] , \_zy_simnet_tvar_53[2].label[72] );
tran (\_zy_simnet_tvar_53[2][80] , \_zy_simnet_tvar_53[2].label[71] );
tran (\_zy_simnet_tvar_53[2][79] , \_zy_simnet_tvar_53[2].label[70] );
tran (\_zy_simnet_tvar_53[2][78] , \_zy_simnet_tvar_53[2].label[69] );
tran (\_zy_simnet_tvar_53[2][77] , \_zy_simnet_tvar_53[2].label[68] );
tran (\_zy_simnet_tvar_53[2][76] , \_zy_simnet_tvar_53[2].label[67] );
tran (\_zy_simnet_tvar_53[2][75] , \_zy_simnet_tvar_53[2].label[66] );
tran (\_zy_simnet_tvar_53[2][74] , \_zy_simnet_tvar_53[2].label[65] );
tran (\_zy_simnet_tvar_53[2][73] , \_zy_simnet_tvar_53[2].label[64] );
tran (\_zy_simnet_tvar_53[2][72] , \_zy_simnet_tvar_53[2].label[63] );
tran (\_zy_simnet_tvar_53[2][71] , \_zy_simnet_tvar_53[2].label[62] );
tran (\_zy_simnet_tvar_53[2][70] , \_zy_simnet_tvar_53[2].label[61] );
tran (\_zy_simnet_tvar_53[2][69] , \_zy_simnet_tvar_53[2].label[60] );
tran (\_zy_simnet_tvar_53[2][68] , \_zy_simnet_tvar_53[2].label[59] );
tran (\_zy_simnet_tvar_53[2][67] , \_zy_simnet_tvar_53[2].label[58] );
tran (\_zy_simnet_tvar_53[2][66] , \_zy_simnet_tvar_53[2].label[57] );
tran (\_zy_simnet_tvar_53[2][65] , \_zy_simnet_tvar_53[2].label[56] );
tran (\_zy_simnet_tvar_53[2][64] , \_zy_simnet_tvar_53[2].label[55] );
tran (\_zy_simnet_tvar_53[2][63] , \_zy_simnet_tvar_53[2].label[54] );
tran (\_zy_simnet_tvar_53[2][62] , \_zy_simnet_tvar_53[2].label[53] );
tran (\_zy_simnet_tvar_53[2][61] , \_zy_simnet_tvar_53[2].label[52] );
tran (\_zy_simnet_tvar_53[2][60] , \_zy_simnet_tvar_53[2].label[51] );
tran (\_zy_simnet_tvar_53[2][59] , \_zy_simnet_tvar_53[2].label[50] );
tran (\_zy_simnet_tvar_53[2][58] , \_zy_simnet_tvar_53[2].label[49] );
tran (\_zy_simnet_tvar_53[2][57] , \_zy_simnet_tvar_53[2].label[48] );
tran (\_zy_simnet_tvar_53[2][56] , \_zy_simnet_tvar_53[2].label[47] );
tran (\_zy_simnet_tvar_53[2][55] , \_zy_simnet_tvar_53[2].label[46] );
tran (\_zy_simnet_tvar_53[2][54] , \_zy_simnet_tvar_53[2].label[45] );
tran (\_zy_simnet_tvar_53[2][53] , \_zy_simnet_tvar_53[2].label[44] );
tran (\_zy_simnet_tvar_53[2][52] , \_zy_simnet_tvar_53[2].label[43] );
tran (\_zy_simnet_tvar_53[2][51] , \_zy_simnet_tvar_53[2].label[42] );
tran (\_zy_simnet_tvar_53[2][50] , \_zy_simnet_tvar_53[2].label[41] );
tran (\_zy_simnet_tvar_53[2][49] , \_zy_simnet_tvar_53[2].label[40] );
tran (\_zy_simnet_tvar_53[2][48] , \_zy_simnet_tvar_53[2].label[39] );
tran (\_zy_simnet_tvar_53[2][47] , \_zy_simnet_tvar_53[2].label[38] );
tran (\_zy_simnet_tvar_53[2][46] , \_zy_simnet_tvar_53[2].label[37] );
tran (\_zy_simnet_tvar_53[2][45] , \_zy_simnet_tvar_53[2].label[36] );
tran (\_zy_simnet_tvar_53[2][44] , \_zy_simnet_tvar_53[2].label[35] );
tran (\_zy_simnet_tvar_53[2][43] , \_zy_simnet_tvar_53[2].label[34] );
tran (\_zy_simnet_tvar_53[2][42] , \_zy_simnet_tvar_53[2].label[33] );
tran (\_zy_simnet_tvar_53[2][41] , \_zy_simnet_tvar_53[2].label[32] );
tran (\_zy_simnet_tvar_53[2][40] , \_zy_simnet_tvar_53[2].label[31] );
tran (\_zy_simnet_tvar_53[2][39] , \_zy_simnet_tvar_53[2].label[30] );
tran (\_zy_simnet_tvar_53[2][38] , \_zy_simnet_tvar_53[2].label[29] );
tran (\_zy_simnet_tvar_53[2][37] , \_zy_simnet_tvar_53[2].label[28] );
tran (\_zy_simnet_tvar_53[2][36] , \_zy_simnet_tvar_53[2].label[27] );
tran (\_zy_simnet_tvar_53[2][35] , \_zy_simnet_tvar_53[2].label[26] );
tran (\_zy_simnet_tvar_53[2][34] , \_zy_simnet_tvar_53[2].label[25] );
tran (\_zy_simnet_tvar_53[2][33] , \_zy_simnet_tvar_53[2].label[24] );
tran (\_zy_simnet_tvar_53[2][32] , \_zy_simnet_tvar_53[2].label[23] );
tran (\_zy_simnet_tvar_53[2][31] , \_zy_simnet_tvar_53[2].label[22] );
tran (\_zy_simnet_tvar_53[2][30] , \_zy_simnet_tvar_53[2].label[21] );
tran (\_zy_simnet_tvar_53[2][29] , \_zy_simnet_tvar_53[2].label[20] );
tran (\_zy_simnet_tvar_53[2][28] , \_zy_simnet_tvar_53[2].label[19] );
tran (\_zy_simnet_tvar_53[2][27] , \_zy_simnet_tvar_53[2].label[18] );
tran (\_zy_simnet_tvar_53[2][26] , \_zy_simnet_tvar_53[2].label[17] );
tran (\_zy_simnet_tvar_53[2][25] , \_zy_simnet_tvar_53[2].label[16] );
tran (\_zy_simnet_tvar_53[2][24] , \_zy_simnet_tvar_53[2].label[15] );
tran (\_zy_simnet_tvar_53[2][23] , \_zy_simnet_tvar_53[2].label[14] );
tran (\_zy_simnet_tvar_53[2][22] , \_zy_simnet_tvar_53[2].label[13] );
tran (\_zy_simnet_tvar_53[2][21] , \_zy_simnet_tvar_53[2].label[12] );
tran (\_zy_simnet_tvar_53[2][20] , \_zy_simnet_tvar_53[2].label[11] );
tran (\_zy_simnet_tvar_53[2][19] , \_zy_simnet_tvar_53[2].label[10] );
tran (\_zy_simnet_tvar_53[2][18] , \_zy_simnet_tvar_53[2].label[9] );
tran (\_zy_simnet_tvar_53[2][17] , \_zy_simnet_tvar_53[2].label[8] );
tran (\_zy_simnet_tvar_53[2][16] , \_zy_simnet_tvar_53[2].label[7] );
tran (\_zy_simnet_tvar_53[2][15] , \_zy_simnet_tvar_53[2].label[6] );
tran (\_zy_simnet_tvar_53[2][14] , \_zy_simnet_tvar_53[2].label[5] );
tran (\_zy_simnet_tvar_53[2][13] , \_zy_simnet_tvar_53[2].label[4] );
tran (\_zy_simnet_tvar_53[2][12] , \_zy_simnet_tvar_53[2].label[3] );
tran (\_zy_simnet_tvar_53[2][11] , \_zy_simnet_tvar_53[2].label[2] );
tran (\_zy_simnet_tvar_53[2][10] , \_zy_simnet_tvar_53[2].label[1] );
tran (\_zy_simnet_tvar_53[2][9] , \_zy_simnet_tvar_53[2].label[0] );
tran (\_zy_simnet_tvar_53[2][8] , \_zy_simnet_tvar_53[2].delimiter_valid[0] );
tran (\_zy_simnet_tvar_53[2][7] , \_zy_simnet_tvar_53[2].delimiter[7] );
tran (\_zy_simnet_tvar_53[2][6] , \_zy_simnet_tvar_53[2].delimiter[6] );
tran (\_zy_simnet_tvar_53[2][5] , \_zy_simnet_tvar_53[2].delimiter[5] );
tran (\_zy_simnet_tvar_53[2][4] , \_zy_simnet_tvar_53[2].delimiter[4] );
tran (\_zy_simnet_tvar_53[2][3] , \_zy_simnet_tvar_53[2].delimiter[3] );
tran (\_zy_simnet_tvar_53[2][2] , \_zy_simnet_tvar_53[2].delimiter[2] );
tran (\_zy_simnet_tvar_53[2][1] , \_zy_simnet_tvar_53[2].delimiter[1] );
tran (\_zy_simnet_tvar_53[2][0] , \_zy_simnet_tvar_53[2].delimiter[0] );
tran (\_zy_simnet_tvar_53[1][271] , \_zy_simnet_tvar_53[1].guid_size[0] );
tran (\_zy_simnet_tvar_53[1][270] , \_zy_simnet_tvar_53[1].label_size[5] );
tran (\_zy_simnet_tvar_53[1][269] , \_zy_simnet_tvar_53[1].label_size[4] );
tran (\_zy_simnet_tvar_53[1][268] , \_zy_simnet_tvar_53[1].label_size[3] );
tran (\_zy_simnet_tvar_53[1][267] , \_zy_simnet_tvar_53[1].label_size[2] );
tran (\_zy_simnet_tvar_53[1][266] , \_zy_simnet_tvar_53[1].label_size[1] );
tran (\_zy_simnet_tvar_53[1][265] , \_zy_simnet_tvar_53[1].label_size[0] );
tran (\_zy_simnet_tvar_53[1][264] , \_zy_simnet_tvar_53[1].label[255] );
tran (\_zy_simnet_tvar_53[1][263] , \_zy_simnet_tvar_53[1].label[254] );
tran (\_zy_simnet_tvar_53[1][262] , \_zy_simnet_tvar_53[1].label[253] );
tran (\_zy_simnet_tvar_53[1][261] , \_zy_simnet_tvar_53[1].label[252] );
tran (\_zy_simnet_tvar_53[1][260] , \_zy_simnet_tvar_53[1].label[251] );
tran (\_zy_simnet_tvar_53[1][259] , \_zy_simnet_tvar_53[1].label[250] );
tran (\_zy_simnet_tvar_53[1][258] , \_zy_simnet_tvar_53[1].label[249] );
tran (\_zy_simnet_tvar_53[1][257] , \_zy_simnet_tvar_53[1].label[248] );
tran (\_zy_simnet_tvar_53[1][256] , \_zy_simnet_tvar_53[1].label[247] );
tran (\_zy_simnet_tvar_53[1][255] , \_zy_simnet_tvar_53[1].label[246] );
tran (\_zy_simnet_tvar_53[1][254] , \_zy_simnet_tvar_53[1].label[245] );
tran (\_zy_simnet_tvar_53[1][253] , \_zy_simnet_tvar_53[1].label[244] );
tran (\_zy_simnet_tvar_53[1][252] , \_zy_simnet_tvar_53[1].label[243] );
tran (\_zy_simnet_tvar_53[1][251] , \_zy_simnet_tvar_53[1].label[242] );
tran (\_zy_simnet_tvar_53[1][250] , \_zy_simnet_tvar_53[1].label[241] );
tran (\_zy_simnet_tvar_53[1][249] , \_zy_simnet_tvar_53[1].label[240] );
tran (\_zy_simnet_tvar_53[1][248] , \_zy_simnet_tvar_53[1].label[239] );
tran (\_zy_simnet_tvar_53[1][247] , \_zy_simnet_tvar_53[1].label[238] );
tran (\_zy_simnet_tvar_53[1][246] , \_zy_simnet_tvar_53[1].label[237] );
tran (\_zy_simnet_tvar_53[1][245] , \_zy_simnet_tvar_53[1].label[236] );
tran (\_zy_simnet_tvar_53[1][244] , \_zy_simnet_tvar_53[1].label[235] );
tran (\_zy_simnet_tvar_53[1][243] , \_zy_simnet_tvar_53[1].label[234] );
tran (\_zy_simnet_tvar_53[1][242] , \_zy_simnet_tvar_53[1].label[233] );
tran (\_zy_simnet_tvar_53[1][241] , \_zy_simnet_tvar_53[1].label[232] );
tran (\_zy_simnet_tvar_53[1][240] , \_zy_simnet_tvar_53[1].label[231] );
tran (\_zy_simnet_tvar_53[1][239] , \_zy_simnet_tvar_53[1].label[230] );
tran (\_zy_simnet_tvar_53[1][238] , \_zy_simnet_tvar_53[1].label[229] );
tran (\_zy_simnet_tvar_53[1][237] , \_zy_simnet_tvar_53[1].label[228] );
tran (\_zy_simnet_tvar_53[1][236] , \_zy_simnet_tvar_53[1].label[227] );
tran (\_zy_simnet_tvar_53[1][235] , \_zy_simnet_tvar_53[1].label[226] );
tran (\_zy_simnet_tvar_53[1][234] , \_zy_simnet_tvar_53[1].label[225] );
tran (\_zy_simnet_tvar_53[1][233] , \_zy_simnet_tvar_53[1].label[224] );
tran (\_zy_simnet_tvar_53[1][232] , \_zy_simnet_tvar_53[1].label[223] );
tran (\_zy_simnet_tvar_53[1][231] , \_zy_simnet_tvar_53[1].label[222] );
tran (\_zy_simnet_tvar_53[1][230] , \_zy_simnet_tvar_53[1].label[221] );
tran (\_zy_simnet_tvar_53[1][229] , \_zy_simnet_tvar_53[1].label[220] );
tran (\_zy_simnet_tvar_53[1][228] , \_zy_simnet_tvar_53[1].label[219] );
tran (\_zy_simnet_tvar_53[1][227] , \_zy_simnet_tvar_53[1].label[218] );
tran (\_zy_simnet_tvar_53[1][226] , \_zy_simnet_tvar_53[1].label[217] );
tran (\_zy_simnet_tvar_53[1][225] , \_zy_simnet_tvar_53[1].label[216] );
tran (\_zy_simnet_tvar_53[1][224] , \_zy_simnet_tvar_53[1].label[215] );
tran (\_zy_simnet_tvar_53[1][223] , \_zy_simnet_tvar_53[1].label[214] );
tran (\_zy_simnet_tvar_53[1][222] , \_zy_simnet_tvar_53[1].label[213] );
tran (\_zy_simnet_tvar_53[1][221] , \_zy_simnet_tvar_53[1].label[212] );
tran (\_zy_simnet_tvar_53[1][220] , \_zy_simnet_tvar_53[1].label[211] );
tran (\_zy_simnet_tvar_53[1][219] , \_zy_simnet_tvar_53[1].label[210] );
tran (\_zy_simnet_tvar_53[1][218] , \_zy_simnet_tvar_53[1].label[209] );
tran (\_zy_simnet_tvar_53[1][217] , \_zy_simnet_tvar_53[1].label[208] );
tran (\_zy_simnet_tvar_53[1][216] , \_zy_simnet_tvar_53[1].label[207] );
tran (\_zy_simnet_tvar_53[1][215] , \_zy_simnet_tvar_53[1].label[206] );
tran (\_zy_simnet_tvar_53[1][214] , \_zy_simnet_tvar_53[1].label[205] );
tran (\_zy_simnet_tvar_53[1][213] , \_zy_simnet_tvar_53[1].label[204] );
tran (\_zy_simnet_tvar_53[1][212] , \_zy_simnet_tvar_53[1].label[203] );
tran (\_zy_simnet_tvar_53[1][211] , \_zy_simnet_tvar_53[1].label[202] );
tran (\_zy_simnet_tvar_53[1][210] , \_zy_simnet_tvar_53[1].label[201] );
tran (\_zy_simnet_tvar_53[1][209] , \_zy_simnet_tvar_53[1].label[200] );
tran (\_zy_simnet_tvar_53[1][208] , \_zy_simnet_tvar_53[1].label[199] );
tran (\_zy_simnet_tvar_53[1][207] , \_zy_simnet_tvar_53[1].label[198] );
tran (\_zy_simnet_tvar_53[1][206] , \_zy_simnet_tvar_53[1].label[197] );
tran (\_zy_simnet_tvar_53[1][205] , \_zy_simnet_tvar_53[1].label[196] );
tran (\_zy_simnet_tvar_53[1][204] , \_zy_simnet_tvar_53[1].label[195] );
tran (\_zy_simnet_tvar_53[1][203] , \_zy_simnet_tvar_53[1].label[194] );
tran (\_zy_simnet_tvar_53[1][202] , \_zy_simnet_tvar_53[1].label[193] );
tran (\_zy_simnet_tvar_53[1][201] , \_zy_simnet_tvar_53[1].label[192] );
tran (\_zy_simnet_tvar_53[1][200] , \_zy_simnet_tvar_53[1].label[191] );
tran (\_zy_simnet_tvar_53[1][199] , \_zy_simnet_tvar_53[1].label[190] );
tran (\_zy_simnet_tvar_53[1][198] , \_zy_simnet_tvar_53[1].label[189] );
tran (\_zy_simnet_tvar_53[1][197] , \_zy_simnet_tvar_53[1].label[188] );
tran (\_zy_simnet_tvar_53[1][196] , \_zy_simnet_tvar_53[1].label[187] );
tran (\_zy_simnet_tvar_53[1][195] , \_zy_simnet_tvar_53[1].label[186] );
tran (\_zy_simnet_tvar_53[1][194] , \_zy_simnet_tvar_53[1].label[185] );
tran (\_zy_simnet_tvar_53[1][193] , \_zy_simnet_tvar_53[1].label[184] );
tran (\_zy_simnet_tvar_53[1][192] , \_zy_simnet_tvar_53[1].label[183] );
tran (\_zy_simnet_tvar_53[1][191] , \_zy_simnet_tvar_53[1].label[182] );
tran (\_zy_simnet_tvar_53[1][190] , \_zy_simnet_tvar_53[1].label[181] );
tran (\_zy_simnet_tvar_53[1][189] , \_zy_simnet_tvar_53[1].label[180] );
tran (\_zy_simnet_tvar_53[1][188] , \_zy_simnet_tvar_53[1].label[179] );
tran (\_zy_simnet_tvar_53[1][187] , \_zy_simnet_tvar_53[1].label[178] );
tran (\_zy_simnet_tvar_53[1][186] , \_zy_simnet_tvar_53[1].label[177] );
tran (\_zy_simnet_tvar_53[1][185] , \_zy_simnet_tvar_53[1].label[176] );
tran (\_zy_simnet_tvar_53[1][184] , \_zy_simnet_tvar_53[1].label[175] );
tran (\_zy_simnet_tvar_53[1][183] , \_zy_simnet_tvar_53[1].label[174] );
tran (\_zy_simnet_tvar_53[1][182] , \_zy_simnet_tvar_53[1].label[173] );
tran (\_zy_simnet_tvar_53[1][181] , \_zy_simnet_tvar_53[1].label[172] );
tran (\_zy_simnet_tvar_53[1][180] , \_zy_simnet_tvar_53[1].label[171] );
tran (\_zy_simnet_tvar_53[1][179] , \_zy_simnet_tvar_53[1].label[170] );
tran (\_zy_simnet_tvar_53[1][178] , \_zy_simnet_tvar_53[1].label[169] );
tran (\_zy_simnet_tvar_53[1][177] , \_zy_simnet_tvar_53[1].label[168] );
tran (\_zy_simnet_tvar_53[1][176] , \_zy_simnet_tvar_53[1].label[167] );
tran (\_zy_simnet_tvar_53[1][175] , \_zy_simnet_tvar_53[1].label[166] );
tran (\_zy_simnet_tvar_53[1][174] , \_zy_simnet_tvar_53[1].label[165] );
tran (\_zy_simnet_tvar_53[1][173] , \_zy_simnet_tvar_53[1].label[164] );
tran (\_zy_simnet_tvar_53[1][172] , \_zy_simnet_tvar_53[1].label[163] );
tran (\_zy_simnet_tvar_53[1][171] , \_zy_simnet_tvar_53[1].label[162] );
tran (\_zy_simnet_tvar_53[1][170] , \_zy_simnet_tvar_53[1].label[161] );
tran (\_zy_simnet_tvar_53[1][169] , \_zy_simnet_tvar_53[1].label[160] );
tran (\_zy_simnet_tvar_53[1][168] , \_zy_simnet_tvar_53[1].label[159] );
tran (\_zy_simnet_tvar_53[1][167] , \_zy_simnet_tvar_53[1].label[158] );
tran (\_zy_simnet_tvar_53[1][166] , \_zy_simnet_tvar_53[1].label[157] );
tran (\_zy_simnet_tvar_53[1][165] , \_zy_simnet_tvar_53[1].label[156] );
tran (\_zy_simnet_tvar_53[1][164] , \_zy_simnet_tvar_53[1].label[155] );
tran (\_zy_simnet_tvar_53[1][163] , \_zy_simnet_tvar_53[1].label[154] );
tran (\_zy_simnet_tvar_53[1][162] , \_zy_simnet_tvar_53[1].label[153] );
tran (\_zy_simnet_tvar_53[1][161] , \_zy_simnet_tvar_53[1].label[152] );
tran (\_zy_simnet_tvar_53[1][160] , \_zy_simnet_tvar_53[1].label[151] );
tran (\_zy_simnet_tvar_53[1][159] , \_zy_simnet_tvar_53[1].label[150] );
tran (\_zy_simnet_tvar_53[1][158] , \_zy_simnet_tvar_53[1].label[149] );
tran (\_zy_simnet_tvar_53[1][157] , \_zy_simnet_tvar_53[1].label[148] );
tran (\_zy_simnet_tvar_53[1][156] , \_zy_simnet_tvar_53[1].label[147] );
tran (\_zy_simnet_tvar_53[1][155] , \_zy_simnet_tvar_53[1].label[146] );
tran (\_zy_simnet_tvar_53[1][154] , \_zy_simnet_tvar_53[1].label[145] );
tran (\_zy_simnet_tvar_53[1][153] , \_zy_simnet_tvar_53[1].label[144] );
tran (\_zy_simnet_tvar_53[1][152] , \_zy_simnet_tvar_53[1].label[143] );
tran (\_zy_simnet_tvar_53[1][151] , \_zy_simnet_tvar_53[1].label[142] );
tran (\_zy_simnet_tvar_53[1][150] , \_zy_simnet_tvar_53[1].label[141] );
tran (\_zy_simnet_tvar_53[1][149] , \_zy_simnet_tvar_53[1].label[140] );
tran (\_zy_simnet_tvar_53[1][148] , \_zy_simnet_tvar_53[1].label[139] );
tran (\_zy_simnet_tvar_53[1][147] , \_zy_simnet_tvar_53[1].label[138] );
tran (\_zy_simnet_tvar_53[1][146] , \_zy_simnet_tvar_53[1].label[137] );
tran (\_zy_simnet_tvar_53[1][145] , \_zy_simnet_tvar_53[1].label[136] );
tran (\_zy_simnet_tvar_53[1][144] , \_zy_simnet_tvar_53[1].label[135] );
tran (\_zy_simnet_tvar_53[1][143] , \_zy_simnet_tvar_53[1].label[134] );
tran (\_zy_simnet_tvar_53[1][142] , \_zy_simnet_tvar_53[1].label[133] );
tran (\_zy_simnet_tvar_53[1][141] , \_zy_simnet_tvar_53[1].label[132] );
tran (\_zy_simnet_tvar_53[1][140] , \_zy_simnet_tvar_53[1].label[131] );
tran (\_zy_simnet_tvar_53[1][139] , \_zy_simnet_tvar_53[1].label[130] );
tran (\_zy_simnet_tvar_53[1][138] , \_zy_simnet_tvar_53[1].label[129] );
tran (\_zy_simnet_tvar_53[1][137] , \_zy_simnet_tvar_53[1].label[128] );
tran (\_zy_simnet_tvar_53[1][136] , \_zy_simnet_tvar_53[1].label[127] );
tran (\_zy_simnet_tvar_53[1][135] , \_zy_simnet_tvar_53[1].label[126] );
tran (\_zy_simnet_tvar_53[1][134] , \_zy_simnet_tvar_53[1].label[125] );
tran (\_zy_simnet_tvar_53[1][133] , \_zy_simnet_tvar_53[1].label[124] );
tran (\_zy_simnet_tvar_53[1][132] , \_zy_simnet_tvar_53[1].label[123] );
tran (\_zy_simnet_tvar_53[1][131] , \_zy_simnet_tvar_53[1].label[122] );
tran (\_zy_simnet_tvar_53[1][130] , \_zy_simnet_tvar_53[1].label[121] );
tran (\_zy_simnet_tvar_53[1][129] , \_zy_simnet_tvar_53[1].label[120] );
tran (\_zy_simnet_tvar_53[1][128] , \_zy_simnet_tvar_53[1].label[119] );
tran (\_zy_simnet_tvar_53[1][127] , \_zy_simnet_tvar_53[1].label[118] );
tran (\_zy_simnet_tvar_53[1][126] , \_zy_simnet_tvar_53[1].label[117] );
tran (\_zy_simnet_tvar_53[1][125] , \_zy_simnet_tvar_53[1].label[116] );
tran (\_zy_simnet_tvar_53[1][124] , \_zy_simnet_tvar_53[1].label[115] );
tran (\_zy_simnet_tvar_53[1][123] , \_zy_simnet_tvar_53[1].label[114] );
tran (\_zy_simnet_tvar_53[1][122] , \_zy_simnet_tvar_53[1].label[113] );
tran (\_zy_simnet_tvar_53[1][121] , \_zy_simnet_tvar_53[1].label[112] );
tran (\_zy_simnet_tvar_53[1][120] , \_zy_simnet_tvar_53[1].label[111] );
tran (\_zy_simnet_tvar_53[1][119] , \_zy_simnet_tvar_53[1].label[110] );
tran (\_zy_simnet_tvar_53[1][118] , \_zy_simnet_tvar_53[1].label[109] );
tran (\_zy_simnet_tvar_53[1][117] , \_zy_simnet_tvar_53[1].label[108] );
tran (\_zy_simnet_tvar_53[1][116] , \_zy_simnet_tvar_53[1].label[107] );
tran (\_zy_simnet_tvar_53[1][115] , \_zy_simnet_tvar_53[1].label[106] );
tran (\_zy_simnet_tvar_53[1][114] , \_zy_simnet_tvar_53[1].label[105] );
tran (\_zy_simnet_tvar_53[1][113] , \_zy_simnet_tvar_53[1].label[104] );
tran (\_zy_simnet_tvar_53[1][112] , \_zy_simnet_tvar_53[1].label[103] );
tran (\_zy_simnet_tvar_53[1][111] , \_zy_simnet_tvar_53[1].label[102] );
tran (\_zy_simnet_tvar_53[1][110] , \_zy_simnet_tvar_53[1].label[101] );
tran (\_zy_simnet_tvar_53[1][109] , \_zy_simnet_tvar_53[1].label[100] );
tran (\_zy_simnet_tvar_53[1][108] , \_zy_simnet_tvar_53[1].label[99] );
tran (\_zy_simnet_tvar_53[1][107] , \_zy_simnet_tvar_53[1].label[98] );
tran (\_zy_simnet_tvar_53[1][106] , \_zy_simnet_tvar_53[1].label[97] );
tran (\_zy_simnet_tvar_53[1][105] , \_zy_simnet_tvar_53[1].label[96] );
tran (\_zy_simnet_tvar_53[1][104] , \_zy_simnet_tvar_53[1].label[95] );
tran (\_zy_simnet_tvar_53[1][103] , \_zy_simnet_tvar_53[1].label[94] );
tran (\_zy_simnet_tvar_53[1][102] , \_zy_simnet_tvar_53[1].label[93] );
tran (\_zy_simnet_tvar_53[1][101] , \_zy_simnet_tvar_53[1].label[92] );
tran (\_zy_simnet_tvar_53[1][100] , \_zy_simnet_tvar_53[1].label[91] );
tran (\_zy_simnet_tvar_53[1][99] , \_zy_simnet_tvar_53[1].label[90] );
tran (\_zy_simnet_tvar_53[1][98] , \_zy_simnet_tvar_53[1].label[89] );
tran (\_zy_simnet_tvar_53[1][97] , \_zy_simnet_tvar_53[1].label[88] );
tran (\_zy_simnet_tvar_53[1][96] , \_zy_simnet_tvar_53[1].label[87] );
tran (\_zy_simnet_tvar_53[1][95] , \_zy_simnet_tvar_53[1].label[86] );
tran (\_zy_simnet_tvar_53[1][94] , \_zy_simnet_tvar_53[1].label[85] );
tran (\_zy_simnet_tvar_53[1][93] , \_zy_simnet_tvar_53[1].label[84] );
tran (\_zy_simnet_tvar_53[1][92] , \_zy_simnet_tvar_53[1].label[83] );
tran (\_zy_simnet_tvar_53[1][91] , \_zy_simnet_tvar_53[1].label[82] );
tran (\_zy_simnet_tvar_53[1][90] , \_zy_simnet_tvar_53[1].label[81] );
tran (\_zy_simnet_tvar_53[1][89] , \_zy_simnet_tvar_53[1].label[80] );
tran (\_zy_simnet_tvar_53[1][88] , \_zy_simnet_tvar_53[1].label[79] );
tran (\_zy_simnet_tvar_53[1][87] , \_zy_simnet_tvar_53[1].label[78] );
tran (\_zy_simnet_tvar_53[1][86] , \_zy_simnet_tvar_53[1].label[77] );
tran (\_zy_simnet_tvar_53[1][85] , \_zy_simnet_tvar_53[1].label[76] );
tran (\_zy_simnet_tvar_53[1][84] , \_zy_simnet_tvar_53[1].label[75] );
tran (\_zy_simnet_tvar_53[1][83] , \_zy_simnet_tvar_53[1].label[74] );
tran (\_zy_simnet_tvar_53[1][82] , \_zy_simnet_tvar_53[1].label[73] );
tran (\_zy_simnet_tvar_53[1][81] , \_zy_simnet_tvar_53[1].label[72] );
tran (\_zy_simnet_tvar_53[1][80] , \_zy_simnet_tvar_53[1].label[71] );
tran (\_zy_simnet_tvar_53[1][79] , \_zy_simnet_tvar_53[1].label[70] );
tran (\_zy_simnet_tvar_53[1][78] , \_zy_simnet_tvar_53[1].label[69] );
tran (\_zy_simnet_tvar_53[1][77] , \_zy_simnet_tvar_53[1].label[68] );
tran (\_zy_simnet_tvar_53[1][76] , \_zy_simnet_tvar_53[1].label[67] );
tran (\_zy_simnet_tvar_53[1][75] , \_zy_simnet_tvar_53[1].label[66] );
tran (\_zy_simnet_tvar_53[1][74] , \_zy_simnet_tvar_53[1].label[65] );
tran (\_zy_simnet_tvar_53[1][73] , \_zy_simnet_tvar_53[1].label[64] );
tran (\_zy_simnet_tvar_53[1][72] , \_zy_simnet_tvar_53[1].label[63] );
tran (\_zy_simnet_tvar_53[1][71] , \_zy_simnet_tvar_53[1].label[62] );
tran (\_zy_simnet_tvar_53[1][70] , \_zy_simnet_tvar_53[1].label[61] );
tran (\_zy_simnet_tvar_53[1][69] , \_zy_simnet_tvar_53[1].label[60] );
tran (\_zy_simnet_tvar_53[1][68] , \_zy_simnet_tvar_53[1].label[59] );
tran (\_zy_simnet_tvar_53[1][67] , \_zy_simnet_tvar_53[1].label[58] );
tran (\_zy_simnet_tvar_53[1][66] , \_zy_simnet_tvar_53[1].label[57] );
tran (\_zy_simnet_tvar_53[1][65] , \_zy_simnet_tvar_53[1].label[56] );
tran (\_zy_simnet_tvar_53[1][64] , \_zy_simnet_tvar_53[1].label[55] );
tran (\_zy_simnet_tvar_53[1][63] , \_zy_simnet_tvar_53[1].label[54] );
tran (\_zy_simnet_tvar_53[1][62] , \_zy_simnet_tvar_53[1].label[53] );
tran (\_zy_simnet_tvar_53[1][61] , \_zy_simnet_tvar_53[1].label[52] );
tran (\_zy_simnet_tvar_53[1][60] , \_zy_simnet_tvar_53[1].label[51] );
tran (\_zy_simnet_tvar_53[1][59] , \_zy_simnet_tvar_53[1].label[50] );
tran (\_zy_simnet_tvar_53[1][58] , \_zy_simnet_tvar_53[1].label[49] );
tran (\_zy_simnet_tvar_53[1][57] , \_zy_simnet_tvar_53[1].label[48] );
tran (\_zy_simnet_tvar_53[1][56] , \_zy_simnet_tvar_53[1].label[47] );
tran (\_zy_simnet_tvar_53[1][55] , \_zy_simnet_tvar_53[1].label[46] );
tran (\_zy_simnet_tvar_53[1][54] , \_zy_simnet_tvar_53[1].label[45] );
tran (\_zy_simnet_tvar_53[1][53] , \_zy_simnet_tvar_53[1].label[44] );
tran (\_zy_simnet_tvar_53[1][52] , \_zy_simnet_tvar_53[1].label[43] );
tran (\_zy_simnet_tvar_53[1][51] , \_zy_simnet_tvar_53[1].label[42] );
tran (\_zy_simnet_tvar_53[1][50] , \_zy_simnet_tvar_53[1].label[41] );
tran (\_zy_simnet_tvar_53[1][49] , \_zy_simnet_tvar_53[1].label[40] );
tran (\_zy_simnet_tvar_53[1][48] , \_zy_simnet_tvar_53[1].label[39] );
tran (\_zy_simnet_tvar_53[1][47] , \_zy_simnet_tvar_53[1].label[38] );
tran (\_zy_simnet_tvar_53[1][46] , \_zy_simnet_tvar_53[1].label[37] );
tran (\_zy_simnet_tvar_53[1][45] , \_zy_simnet_tvar_53[1].label[36] );
tran (\_zy_simnet_tvar_53[1][44] , \_zy_simnet_tvar_53[1].label[35] );
tran (\_zy_simnet_tvar_53[1][43] , \_zy_simnet_tvar_53[1].label[34] );
tran (\_zy_simnet_tvar_53[1][42] , \_zy_simnet_tvar_53[1].label[33] );
tran (\_zy_simnet_tvar_53[1][41] , \_zy_simnet_tvar_53[1].label[32] );
tran (\_zy_simnet_tvar_53[1][40] , \_zy_simnet_tvar_53[1].label[31] );
tran (\_zy_simnet_tvar_53[1][39] , \_zy_simnet_tvar_53[1].label[30] );
tran (\_zy_simnet_tvar_53[1][38] , \_zy_simnet_tvar_53[1].label[29] );
tran (\_zy_simnet_tvar_53[1][37] , \_zy_simnet_tvar_53[1].label[28] );
tran (\_zy_simnet_tvar_53[1][36] , \_zy_simnet_tvar_53[1].label[27] );
tran (\_zy_simnet_tvar_53[1][35] , \_zy_simnet_tvar_53[1].label[26] );
tran (\_zy_simnet_tvar_53[1][34] , \_zy_simnet_tvar_53[1].label[25] );
tran (\_zy_simnet_tvar_53[1][33] , \_zy_simnet_tvar_53[1].label[24] );
tran (\_zy_simnet_tvar_53[1][32] , \_zy_simnet_tvar_53[1].label[23] );
tran (\_zy_simnet_tvar_53[1][31] , \_zy_simnet_tvar_53[1].label[22] );
tran (\_zy_simnet_tvar_53[1][30] , \_zy_simnet_tvar_53[1].label[21] );
tran (\_zy_simnet_tvar_53[1][29] , \_zy_simnet_tvar_53[1].label[20] );
tran (\_zy_simnet_tvar_53[1][28] , \_zy_simnet_tvar_53[1].label[19] );
tran (\_zy_simnet_tvar_53[1][27] , \_zy_simnet_tvar_53[1].label[18] );
tran (\_zy_simnet_tvar_53[1][26] , \_zy_simnet_tvar_53[1].label[17] );
tran (\_zy_simnet_tvar_53[1][25] , \_zy_simnet_tvar_53[1].label[16] );
tran (\_zy_simnet_tvar_53[1][24] , \_zy_simnet_tvar_53[1].label[15] );
tran (\_zy_simnet_tvar_53[1][23] , \_zy_simnet_tvar_53[1].label[14] );
tran (\_zy_simnet_tvar_53[1][22] , \_zy_simnet_tvar_53[1].label[13] );
tran (\_zy_simnet_tvar_53[1][21] , \_zy_simnet_tvar_53[1].label[12] );
tran (\_zy_simnet_tvar_53[1][20] , \_zy_simnet_tvar_53[1].label[11] );
tran (\_zy_simnet_tvar_53[1][19] , \_zy_simnet_tvar_53[1].label[10] );
tran (\_zy_simnet_tvar_53[1][18] , \_zy_simnet_tvar_53[1].label[9] );
tran (\_zy_simnet_tvar_53[1][17] , \_zy_simnet_tvar_53[1].label[8] );
tran (\_zy_simnet_tvar_53[1][16] , \_zy_simnet_tvar_53[1].label[7] );
tran (\_zy_simnet_tvar_53[1][15] , \_zy_simnet_tvar_53[1].label[6] );
tran (\_zy_simnet_tvar_53[1][14] , \_zy_simnet_tvar_53[1].label[5] );
tran (\_zy_simnet_tvar_53[1][13] , \_zy_simnet_tvar_53[1].label[4] );
tran (\_zy_simnet_tvar_53[1][12] , \_zy_simnet_tvar_53[1].label[3] );
tran (\_zy_simnet_tvar_53[1][11] , \_zy_simnet_tvar_53[1].label[2] );
tran (\_zy_simnet_tvar_53[1][10] , \_zy_simnet_tvar_53[1].label[1] );
tran (\_zy_simnet_tvar_53[1][9] , \_zy_simnet_tvar_53[1].label[0] );
tran (\_zy_simnet_tvar_53[1][8] , \_zy_simnet_tvar_53[1].delimiter_valid[0] );
tran (\_zy_simnet_tvar_53[1][7] , \_zy_simnet_tvar_53[1].delimiter[7] );
tran (\_zy_simnet_tvar_53[1][6] , \_zy_simnet_tvar_53[1].delimiter[6] );
tran (\_zy_simnet_tvar_53[1][5] , \_zy_simnet_tvar_53[1].delimiter[5] );
tran (\_zy_simnet_tvar_53[1][4] , \_zy_simnet_tvar_53[1].delimiter[4] );
tran (\_zy_simnet_tvar_53[1][3] , \_zy_simnet_tvar_53[1].delimiter[3] );
tran (\_zy_simnet_tvar_53[1][2] , \_zy_simnet_tvar_53[1].delimiter[2] );
tran (\_zy_simnet_tvar_53[1][1] , \_zy_simnet_tvar_53[1].delimiter[1] );
tran (\_zy_simnet_tvar_53[1][0] , \_zy_simnet_tvar_53[1].delimiter[0] );
tran (\_zy_simnet_tvar_53[0][271] , \_zy_simnet_tvar_53[0].guid_size[0] );
tran (\_zy_simnet_tvar_53[0][270] , \_zy_simnet_tvar_53[0].label_size[5] );
tran (\_zy_simnet_tvar_53[0][269] , \_zy_simnet_tvar_53[0].label_size[4] );
tran (\_zy_simnet_tvar_53[0][268] , \_zy_simnet_tvar_53[0].label_size[3] );
tran (\_zy_simnet_tvar_53[0][267] , \_zy_simnet_tvar_53[0].label_size[2] );
tran (\_zy_simnet_tvar_53[0][266] , \_zy_simnet_tvar_53[0].label_size[1] );
tran (\_zy_simnet_tvar_53[0][265] , \_zy_simnet_tvar_53[0].label_size[0] );
tran (\_zy_simnet_tvar_53[0][264] , \_zy_simnet_tvar_53[0].label[255] );
tran (\_zy_simnet_tvar_53[0][263] , \_zy_simnet_tvar_53[0].label[254] );
tran (\_zy_simnet_tvar_53[0][262] , \_zy_simnet_tvar_53[0].label[253] );
tran (\_zy_simnet_tvar_53[0][261] , \_zy_simnet_tvar_53[0].label[252] );
tran (\_zy_simnet_tvar_53[0][260] , \_zy_simnet_tvar_53[0].label[251] );
tran (\_zy_simnet_tvar_53[0][259] , \_zy_simnet_tvar_53[0].label[250] );
tran (\_zy_simnet_tvar_53[0][258] , \_zy_simnet_tvar_53[0].label[249] );
tran (\_zy_simnet_tvar_53[0][257] , \_zy_simnet_tvar_53[0].label[248] );
tran (\_zy_simnet_tvar_53[0][256] , \_zy_simnet_tvar_53[0].label[247] );
tran (\_zy_simnet_tvar_53[0][255] , \_zy_simnet_tvar_53[0].label[246] );
tran (\_zy_simnet_tvar_53[0][254] , \_zy_simnet_tvar_53[0].label[245] );
tran (\_zy_simnet_tvar_53[0][253] , \_zy_simnet_tvar_53[0].label[244] );
tran (\_zy_simnet_tvar_53[0][252] , \_zy_simnet_tvar_53[0].label[243] );
tran (\_zy_simnet_tvar_53[0][251] , \_zy_simnet_tvar_53[0].label[242] );
tran (\_zy_simnet_tvar_53[0][250] , \_zy_simnet_tvar_53[0].label[241] );
tran (\_zy_simnet_tvar_53[0][249] , \_zy_simnet_tvar_53[0].label[240] );
tran (\_zy_simnet_tvar_53[0][248] , \_zy_simnet_tvar_53[0].label[239] );
tran (\_zy_simnet_tvar_53[0][247] , \_zy_simnet_tvar_53[0].label[238] );
tran (\_zy_simnet_tvar_53[0][246] , \_zy_simnet_tvar_53[0].label[237] );
tran (\_zy_simnet_tvar_53[0][245] , \_zy_simnet_tvar_53[0].label[236] );
tran (\_zy_simnet_tvar_53[0][244] , \_zy_simnet_tvar_53[0].label[235] );
tran (\_zy_simnet_tvar_53[0][243] , \_zy_simnet_tvar_53[0].label[234] );
tran (\_zy_simnet_tvar_53[0][242] , \_zy_simnet_tvar_53[0].label[233] );
tran (\_zy_simnet_tvar_53[0][241] , \_zy_simnet_tvar_53[0].label[232] );
tran (\_zy_simnet_tvar_53[0][240] , \_zy_simnet_tvar_53[0].label[231] );
tran (\_zy_simnet_tvar_53[0][239] , \_zy_simnet_tvar_53[0].label[230] );
tran (\_zy_simnet_tvar_53[0][238] , \_zy_simnet_tvar_53[0].label[229] );
tran (\_zy_simnet_tvar_53[0][237] , \_zy_simnet_tvar_53[0].label[228] );
tran (\_zy_simnet_tvar_53[0][236] , \_zy_simnet_tvar_53[0].label[227] );
tran (\_zy_simnet_tvar_53[0][235] , \_zy_simnet_tvar_53[0].label[226] );
tran (\_zy_simnet_tvar_53[0][234] , \_zy_simnet_tvar_53[0].label[225] );
tran (\_zy_simnet_tvar_53[0][233] , \_zy_simnet_tvar_53[0].label[224] );
tran (\_zy_simnet_tvar_53[0][232] , \_zy_simnet_tvar_53[0].label[223] );
tran (\_zy_simnet_tvar_53[0][231] , \_zy_simnet_tvar_53[0].label[222] );
tran (\_zy_simnet_tvar_53[0][230] , \_zy_simnet_tvar_53[0].label[221] );
tran (\_zy_simnet_tvar_53[0][229] , \_zy_simnet_tvar_53[0].label[220] );
tran (\_zy_simnet_tvar_53[0][228] , \_zy_simnet_tvar_53[0].label[219] );
tran (\_zy_simnet_tvar_53[0][227] , \_zy_simnet_tvar_53[0].label[218] );
tran (\_zy_simnet_tvar_53[0][226] , \_zy_simnet_tvar_53[0].label[217] );
tran (\_zy_simnet_tvar_53[0][225] , \_zy_simnet_tvar_53[0].label[216] );
tran (\_zy_simnet_tvar_53[0][224] , \_zy_simnet_tvar_53[0].label[215] );
tran (\_zy_simnet_tvar_53[0][223] , \_zy_simnet_tvar_53[0].label[214] );
tran (\_zy_simnet_tvar_53[0][222] , \_zy_simnet_tvar_53[0].label[213] );
tran (\_zy_simnet_tvar_53[0][221] , \_zy_simnet_tvar_53[0].label[212] );
tran (\_zy_simnet_tvar_53[0][220] , \_zy_simnet_tvar_53[0].label[211] );
tran (\_zy_simnet_tvar_53[0][219] , \_zy_simnet_tvar_53[0].label[210] );
tran (\_zy_simnet_tvar_53[0][218] , \_zy_simnet_tvar_53[0].label[209] );
tran (\_zy_simnet_tvar_53[0][217] , \_zy_simnet_tvar_53[0].label[208] );
tran (\_zy_simnet_tvar_53[0][216] , \_zy_simnet_tvar_53[0].label[207] );
tran (\_zy_simnet_tvar_53[0][215] , \_zy_simnet_tvar_53[0].label[206] );
tran (\_zy_simnet_tvar_53[0][214] , \_zy_simnet_tvar_53[0].label[205] );
tran (\_zy_simnet_tvar_53[0][213] , \_zy_simnet_tvar_53[0].label[204] );
tran (\_zy_simnet_tvar_53[0][212] , \_zy_simnet_tvar_53[0].label[203] );
tran (\_zy_simnet_tvar_53[0][211] , \_zy_simnet_tvar_53[0].label[202] );
tran (\_zy_simnet_tvar_53[0][210] , \_zy_simnet_tvar_53[0].label[201] );
tran (\_zy_simnet_tvar_53[0][209] , \_zy_simnet_tvar_53[0].label[200] );
tran (\_zy_simnet_tvar_53[0][208] , \_zy_simnet_tvar_53[0].label[199] );
tran (\_zy_simnet_tvar_53[0][207] , \_zy_simnet_tvar_53[0].label[198] );
tran (\_zy_simnet_tvar_53[0][206] , \_zy_simnet_tvar_53[0].label[197] );
tran (\_zy_simnet_tvar_53[0][205] , \_zy_simnet_tvar_53[0].label[196] );
tran (\_zy_simnet_tvar_53[0][204] , \_zy_simnet_tvar_53[0].label[195] );
tran (\_zy_simnet_tvar_53[0][203] , \_zy_simnet_tvar_53[0].label[194] );
tran (\_zy_simnet_tvar_53[0][202] , \_zy_simnet_tvar_53[0].label[193] );
tran (\_zy_simnet_tvar_53[0][201] , \_zy_simnet_tvar_53[0].label[192] );
tran (\_zy_simnet_tvar_53[0][200] , \_zy_simnet_tvar_53[0].label[191] );
tran (\_zy_simnet_tvar_53[0][199] , \_zy_simnet_tvar_53[0].label[190] );
tran (\_zy_simnet_tvar_53[0][198] , \_zy_simnet_tvar_53[0].label[189] );
tran (\_zy_simnet_tvar_53[0][197] , \_zy_simnet_tvar_53[0].label[188] );
tran (\_zy_simnet_tvar_53[0][196] , \_zy_simnet_tvar_53[0].label[187] );
tran (\_zy_simnet_tvar_53[0][195] , \_zy_simnet_tvar_53[0].label[186] );
tran (\_zy_simnet_tvar_53[0][194] , \_zy_simnet_tvar_53[0].label[185] );
tran (\_zy_simnet_tvar_53[0][193] , \_zy_simnet_tvar_53[0].label[184] );
tran (\_zy_simnet_tvar_53[0][192] , \_zy_simnet_tvar_53[0].label[183] );
tran (\_zy_simnet_tvar_53[0][191] , \_zy_simnet_tvar_53[0].label[182] );
tran (\_zy_simnet_tvar_53[0][190] , \_zy_simnet_tvar_53[0].label[181] );
tran (\_zy_simnet_tvar_53[0][189] , \_zy_simnet_tvar_53[0].label[180] );
tran (\_zy_simnet_tvar_53[0][188] , \_zy_simnet_tvar_53[0].label[179] );
tran (\_zy_simnet_tvar_53[0][187] , \_zy_simnet_tvar_53[0].label[178] );
tran (\_zy_simnet_tvar_53[0][186] , \_zy_simnet_tvar_53[0].label[177] );
tran (\_zy_simnet_tvar_53[0][185] , \_zy_simnet_tvar_53[0].label[176] );
tran (\_zy_simnet_tvar_53[0][184] , \_zy_simnet_tvar_53[0].label[175] );
tran (\_zy_simnet_tvar_53[0][183] , \_zy_simnet_tvar_53[0].label[174] );
tran (\_zy_simnet_tvar_53[0][182] , \_zy_simnet_tvar_53[0].label[173] );
tran (\_zy_simnet_tvar_53[0][181] , \_zy_simnet_tvar_53[0].label[172] );
tran (\_zy_simnet_tvar_53[0][180] , \_zy_simnet_tvar_53[0].label[171] );
tran (\_zy_simnet_tvar_53[0][179] , \_zy_simnet_tvar_53[0].label[170] );
tran (\_zy_simnet_tvar_53[0][178] , \_zy_simnet_tvar_53[0].label[169] );
tran (\_zy_simnet_tvar_53[0][177] , \_zy_simnet_tvar_53[0].label[168] );
tran (\_zy_simnet_tvar_53[0][176] , \_zy_simnet_tvar_53[0].label[167] );
tran (\_zy_simnet_tvar_53[0][175] , \_zy_simnet_tvar_53[0].label[166] );
tran (\_zy_simnet_tvar_53[0][174] , \_zy_simnet_tvar_53[0].label[165] );
tran (\_zy_simnet_tvar_53[0][173] , \_zy_simnet_tvar_53[0].label[164] );
tran (\_zy_simnet_tvar_53[0][172] , \_zy_simnet_tvar_53[0].label[163] );
tran (\_zy_simnet_tvar_53[0][171] , \_zy_simnet_tvar_53[0].label[162] );
tran (\_zy_simnet_tvar_53[0][170] , \_zy_simnet_tvar_53[0].label[161] );
tran (\_zy_simnet_tvar_53[0][169] , \_zy_simnet_tvar_53[0].label[160] );
tran (\_zy_simnet_tvar_53[0][168] , \_zy_simnet_tvar_53[0].label[159] );
tran (\_zy_simnet_tvar_53[0][167] , \_zy_simnet_tvar_53[0].label[158] );
tran (\_zy_simnet_tvar_53[0][166] , \_zy_simnet_tvar_53[0].label[157] );
tran (\_zy_simnet_tvar_53[0][165] , \_zy_simnet_tvar_53[0].label[156] );
tran (\_zy_simnet_tvar_53[0][164] , \_zy_simnet_tvar_53[0].label[155] );
tran (\_zy_simnet_tvar_53[0][163] , \_zy_simnet_tvar_53[0].label[154] );
tran (\_zy_simnet_tvar_53[0][162] , \_zy_simnet_tvar_53[0].label[153] );
tran (\_zy_simnet_tvar_53[0][161] , \_zy_simnet_tvar_53[0].label[152] );
tran (\_zy_simnet_tvar_53[0][160] , \_zy_simnet_tvar_53[0].label[151] );
tran (\_zy_simnet_tvar_53[0][159] , \_zy_simnet_tvar_53[0].label[150] );
tran (\_zy_simnet_tvar_53[0][158] , \_zy_simnet_tvar_53[0].label[149] );
tran (\_zy_simnet_tvar_53[0][157] , \_zy_simnet_tvar_53[0].label[148] );
tran (\_zy_simnet_tvar_53[0][156] , \_zy_simnet_tvar_53[0].label[147] );
tran (\_zy_simnet_tvar_53[0][155] , \_zy_simnet_tvar_53[0].label[146] );
tran (\_zy_simnet_tvar_53[0][154] , \_zy_simnet_tvar_53[0].label[145] );
tran (\_zy_simnet_tvar_53[0][153] , \_zy_simnet_tvar_53[0].label[144] );
tran (\_zy_simnet_tvar_53[0][152] , \_zy_simnet_tvar_53[0].label[143] );
tran (\_zy_simnet_tvar_53[0][151] , \_zy_simnet_tvar_53[0].label[142] );
tran (\_zy_simnet_tvar_53[0][150] , \_zy_simnet_tvar_53[0].label[141] );
tran (\_zy_simnet_tvar_53[0][149] , \_zy_simnet_tvar_53[0].label[140] );
tran (\_zy_simnet_tvar_53[0][148] , \_zy_simnet_tvar_53[0].label[139] );
tran (\_zy_simnet_tvar_53[0][147] , \_zy_simnet_tvar_53[0].label[138] );
tran (\_zy_simnet_tvar_53[0][146] , \_zy_simnet_tvar_53[0].label[137] );
tran (\_zy_simnet_tvar_53[0][145] , \_zy_simnet_tvar_53[0].label[136] );
tran (\_zy_simnet_tvar_53[0][144] , \_zy_simnet_tvar_53[0].label[135] );
tran (\_zy_simnet_tvar_53[0][143] , \_zy_simnet_tvar_53[0].label[134] );
tran (\_zy_simnet_tvar_53[0][142] , \_zy_simnet_tvar_53[0].label[133] );
tran (\_zy_simnet_tvar_53[0][141] , \_zy_simnet_tvar_53[0].label[132] );
tran (\_zy_simnet_tvar_53[0][140] , \_zy_simnet_tvar_53[0].label[131] );
tran (\_zy_simnet_tvar_53[0][139] , \_zy_simnet_tvar_53[0].label[130] );
tran (\_zy_simnet_tvar_53[0][138] , \_zy_simnet_tvar_53[0].label[129] );
tran (\_zy_simnet_tvar_53[0][137] , \_zy_simnet_tvar_53[0].label[128] );
tran (\_zy_simnet_tvar_53[0][136] , \_zy_simnet_tvar_53[0].label[127] );
tran (\_zy_simnet_tvar_53[0][135] , \_zy_simnet_tvar_53[0].label[126] );
tran (\_zy_simnet_tvar_53[0][134] , \_zy_simnet_tvar_53[0].label[125] );
tran (\_zy_simnet_tvar_53[0][133] , \_zy_simnet_tvar_53[0].label[124] );
tran (\_zy_simnet_tvar_53[0][132] , \_zy_simnet_tvar_53[0].label[123] );
tran (\_zy_simnet_tvar_53[0][131] , \_zy_simnet_tvar_53[0].label[122] );
tran (\_zy_simnet_tvar_53[0][130] , \_zy_simnet_tvar_53[0].label[121] );
tran (\_zy_simnet_tvar_53[0][129] , \_zy_simnet_tvar_53[0].label[120] );
tran (\_zy_simnet_tvar_53[0][128] , \_zy_simnet_tvar_53[0].label[119] );
tran (\_zy_simnet_tvar_53[0][127] , \_zy_simnet_tvar_53[0].label[118] );
tran (\_zy_simnet_tvar_53[0][126] , \_zy_simnet_tvar_53[0].label[117] );
tran (\_zy_simnet_tvar_53[0][125] , \_zy_simnet_tvar_53[0].label[116] );
tran (\_zy_simnet_tvar_53[0][124] , \_zy_simnet_tvar_53[0].label[115] );
tran (\_zy_simnet_tvar_53[0][123] , \_zy_simnet_tvar_53[0].label[114] );
tran (\_zy_simnet_tvar_53[0][122] , \_zy_simnet_tvar_53[0].label[113] );
tran (\_zy_simnet_tvar_53[0][121] , \_zy_simnet_tvar_53[0].label[112] );
tran (\_zy_simnet_tvar_53[0][120] , \_zy_simnet_tvar_53[0].label[111] );
tran (\_zy_simnet_tvar_53[0][119] , \_zy_simnet_tvar_53[0].label[110] );
tran (\_zy_simnet_tvar_53[0][118] , \_zy_simnet_tvar_53[0].label[109] );
tran (\_zy_simnet_tvar_53[0][117] , \_zy_simnet_tvar_53[0].label[108] );
tran (\_zy_simnet_tvar_53[0][116] , \_zy_simnet_tvar_53[0].label[107] );
tran (\_zy_simnet_tvar_53[0][115] , \_zy_simnet_tvar_53[0].label[106] );
tran (\_zy_simnet_tvar_53[0][114] , \_zy_simnet_tvar_53[0].label[105] );
tran (\_zy_simnet_tvar_53[0][113] , \_zy_simnet_tvar_53[0].label[104] );
tran (\_zy_simnet_tvar_53[0][112] , \_zy_simnet_tvar_53[0].label[103] );
tran (\_zy_simnet_tvar_53[0][111] , \_zy_simnet_tvar_53[0].label[102] );
tran (\_zy_simnet_tvar_53[0][110] , \_zy_simnet_tvar_53[0].label[101] );
tran (\_zy_simnet_tvar_53[0][109] , \_zy_simnet_tvar_53[0].label[100] );
tran (\_zy_simnet_tvar_53[0][108] , \_zy_simnet_tvar_53[0].label[99] );
tran (\_zy_simnet_tvar_53[0][107] , \_zy_simnet_tvar_53[0].label[98] );
tran (\_zy_simnet_tvar_53[0][106] , \_zy_simnet_tvar_53[0].label[97] );
tran (\_zy_simnet_tvar_53[0][105] , \_zy_simnet_tvar_53[0].label[96] );
tran (\_zy_simnet_tvar_53[0][104] , \_zy_simnet_tvar_53[0].label[95] );
tran (\_zy_simnet_tvar_53[0][103] , \_zy_simnet_tvar_53[0].label[94] );
tran (\_zy_simnet_tvar_53[0][102] , \_zy_simnet_tvar_53[0].label[93] );
tran (\_zy_simnet_tvar_53[0][101] , \_zy_simnet_tvar_53[0].label[92] );
tran (\_zy_simnet_tvar_53[0][100] , \_zy_simnet_tvar_53[0].label[91] );
tran (\_zy_simnet_tvar_53[0][99] , \_zy_simnet_tvar_53[0].label[90] );
tran (\_zy_simnet_tvar_53[0][98] , \_zy_simnet_tvar_53[0].label[89] );
tran (\_zy_simnet_tvar_53[0][97] , \_zy_simnet_tvar_53[0].label[88] );
tran (\_zy_simnet_tvar_53[0][96] , \_zy_simnet_tvar_53[0].label[87] );
tran (\_zy_simnet_tvar_53[0][95] , \_zy_simnet_tvar_53[0].label[86] );
tran (\_zy_simnet_tvar_53[0][94] , \_zy_simnet_tvar_53[0].label[85] );
tran (\_zy_simnet_tvar_53[0][93] , \_zy_simnet_tvar_53[0].label[84] );
tran (\_zy_simnet_tvar_53[0][92] , \_zy_simnet_tvar_53[0].label[83] );
tran (\_zy_simnet_tvar_53[0][91] , \_zy_simnet_tvar_53[0].label[82] );
tran (\_zy_simnet_tvar_53[0][90] , \_zy_simnet_tvar_53[0].label[81] );
tran (\_zy_simnet_tvar_53[0][89] , \_zy_simnet_tvar_53[0].label[80] );
tran (\_zy_simnet_tvar_53[0][88] , \_zy_simnet_tvar_53[0].label[79] );
tran (\_zy_simnet_tvar_53[0][87] , \_zy_simnet_tvar_53[0].label[78] );
tran (\_zy_simnet_tvar_53[0][86] , \_zy_simnet_tvar_53[0].label[77] );
tran (\_zy_simnet_tvar_53[0][85] , \_zy_simnet_tvar_53[0].label[76] );
tran (\_zy_simnet_tvar_53[0][84] , \_zy_simnet_tvar_53[0].label[75] );
tran (\_zy_simnet_tvar_53[0][83] , \_zy_simnet_tvar_53[0].label[74] );
tran (\_zy_simnet_tvar_53[0][82] , \_zy_simnet_tvar_53[0].label[73] );
tran (\_zy_simnet_tvar_53[0][81] , \_zy_simnet_tvar_53[0].label[72] );
tran (\_zy_simnet_tvar_53[0][80] , \_zy_simnet_tvar_53[0].label[71] );
tran (\_zy_simnet_tvar_53[0][79] , \_zy_simnet_tvar_53[0].label[70] );
tran (\_zy_simnet_tvar_53[0][78] , \_zy_simnet_tvar_53[0].label[69] );
tran (\_zy_simnet_tvar_53[0][77] , \_zy_simnet_tvar_53[0].label[68] );
tran (\_zy_simnet_tvar_53[0][76] , \_zy_simnet_tvar_53[0].label[67] );
tran (\_zy_simnet_tvar_53[0][75] , \_zy_simnet_tvar_53[0].label[66] );
tran (\_zy_simnet_tvar_53[0][74] , \_zy_simnet_tvar_53[0].label[65] );
tran (\_zy_simnet_tvar_53[0][73] , \_zy_simnet_tvar_53[0].label[64] );
tran (\_zy_simnet_tvar_53[0][72] , \_zy_simnet_tvar_53[0].label[63] );
tran (\_zy_simnet_tvar_53[0][71] , \_zy_simnet_tvar_53[0].label[62] );
tran (\_zy_simnet_tvar_53[0][70] , \_zy_simnet_tvar_53[0].label[61] );
tran (\_zy_simnet_tvar_53[0][69] , \_zy_simnet_tvar_53[0].label[60] );
tran (\_zy_simnet_tvar_53[0][68] , \_zy_simnet_tvar_53[0].label[59] );
tran (\_zy_simnet_tvar_53[0][67] , \_zy_simnet_tvar_53[0].label[58] );
tran (\_zy_simnet_tvar_53[0][66] , \_zy_simnet_tvar_53[0].label[57] );
tran (\_zy_simnet_tvar_53[0][65] , \_zy_simnet_tvar_53[0].label[56] );
tran (\_zy_simnet_tvar_53[0][64] , \_zy_simnet_tvar_53[0].label[55] );
tran (\_zy_simnet_tvar_53[0][63] , \_zy_simnet_tvar_53[0].label[54] );
tran (\_zy_simnet_tvar_53[0][62] , \_zy_simnet_tvar_53[0].label[53] );
tran (\_zy_simnet_tvar_53[0][61] , \_zy_simnet_tvar_53[0].label[52] );
tran (\_zy_simnet_tvar_53[0][60] , \_zy_simnet_tvar_53[0].label[51] );
tran (\_zy_simnet_tvar_53[0][59] , \_zy_simnet_tvar_53[0].label[50] );
tran (\_zy_simnet_tvar_53[0][58] , \_zy_simnet_tvar_53[0].label[49] );
tran (\_zy_simnet_tvar_53[0][57] , \_zy_simnet_tvar_53[0].label[48] );
tran (\_zy_simnet_tvar_53[0][56] , \_zy_simnet_tvar_53[0].label[47] );
tran (\_zy_simnet_tvar_53[0][55] , \_zy_simnet_tvar_53[0].label[46] );
tran (\_zy_simnet_tvar_53[0][54] , \_zy_simnet_tvar_53[0].label[45] );
tran (\_zy_simnet_tvar_53[0][53] , \_zy_simnet_tvar_53[0].label[44] );
tran (\_zy_simnet_tvar_53[0][52] , \_zy_simnet_tvar_53[0].label[43] );
tran (\_zy_simnet_tvar_53[0][51] , \_zy_simnet_tvar_53[0].label[42] );
tran (\_zy_simnet_tvar_53[0][50] , \_zy_simnet_tvar_53[0].label[41] );
tran (\_zy_simnet_tvar_53[0][49] , \_zy_simnet_tvar_53[0].label[40] );
tran (\_zy_simnet_tvar_53[0][48] , \_zy_simnet_tvar_53[0].label[39] );
tran (\_zy_simnet_tvar_53[0][47] , \_zy_simnet_tvar_53[0].label[38] );
tran (\_zy_simnet_tvar_53[0][46] , \_zy_simnet_tvar_53[0].label[37] );
tran (\_zy_simnet_tvar_53[0][45] , \_zy_simnet_tvar_53[0].label[36] );
tran (\_zy_simnet_tvar_53[0][44] , \_zy_simnet_tvar_53[0].label[35] );
tran (\_zy_simnet_tvar_53[0][43] , \_zy_simnet_tvar_53[0].label[34] );
tran (\_zy_simnet_tvar_53[0][42] , \_zy_simnet_tvar_53[0].label[33] );
tran (\_zy_simnet_tvar_53[0][41] , \_zy_simnet_tvar_53[0].label[32] );
tran (\_zy_simnet_tvar_53[0][40] , \_zy_simnet_tvar_53[0].label[31] );
tran (\_zy_simnet_tvar_53[0][39] , \_zy_simnet_tvar_53[0].label[30] );
tran (\_zy_simnet_tvar_53[0][38] , \_zy_simnet_tvar_53[0].label[29] );
tran (\_zy_simnet_tvar_53[0][37] , \_zy_simnet_tvar_53[0].label[28] );
tran (\_zy_simnet_tvar_53[0][36] , \_zy_simnet_tvar_53[0].label[27] );
tran (\_zy_simnet_tvar_53[0][35] , \_zy_simnet_tvar_53[0].label[26] );
tran (\_zy_simnet_tvar_53[0][34] , \_zy_simnet_tvar_53[0].label[25] );
tran (\_zy_simnet_tvar_53[0][33] , \_zy_simnet_tvar_53[0].label[24] );
tran (\_zy_simnet_tvar_53[0][32] , \_zy_simnet_tvar_53[0].label[23] );
tran (\_zy_simnet_tvar_53[0][31] , \_zy_simnet_tvar_53[0].label[22] );
tran (\_zy_simnet_tvar_53[0][30] , \_zy_simnet_tvar_53[0].label[21] );
tran (\_zy_simnet_tvar_53[0][29] , \_zy_simnet_tvar_53[0].label[20] );
tran (\_zy_simnet_tvar_53[0][28] , \_zy_simnet_tvar_53[0].label[19] );
tran (\_zy_simnet_tvar_53[0][27] , \_zy_simnet_tvar_53[0].label[18] );
tran (\_zy_simnet_tvar_53[0][26] , \_zy_simnet_tvar_53[0].label[17] );
tran (\_zy_simnet_tvar_53[0][25] , \_zy_simnet_tvar_53[0].label[16] );
tran (\_zy_simnet_tvar_53[0][24] , \_zy_simnet_tvar_53[0].label[15] );
tran (\_zy_simnet_tvar_53[0][23] , \_zy_simnet_tvar_53[0].label[14] );
tran (\_zy_simnet_tvar_53[0][22] , \_zy_simnet_tvar_53[0].label[13] );
tran (\_zy_simnet_tvar_53[0][21] , \_zy_simnet_tvar_53[0].label[12] );
tran (\_zy_simnet_tvar_53[0][20] , \_zy_simnet_tvar_53[0].label[11] );
tran (\_zy_simnet_tvar_53[0][19] , \_zy_simnet_tvar_53[0].label[10] );
tran (\_zy_simnet_tvar_53[0][18] , \_zy_simnet_tvar_53[0].label[9] );
tran (\_zy_simnet_tvar_53[0][17] , \_zy_simnet_tvar_53[0].label[8] );
tran (\_zy_simnet_tvar_53[0][16] , \_zy_simnet_tvar_53[0].label[7] );
tran (\_zy_simnet_tvar_53[0][15] , \_zy_simnet_tvar_53[0].label[6] );
tran (\_zy_simnet_tvar_53[0][14] , \_zy_simnet_tvar_53[0].label[5] );
tran (\_zy_simnet_tvar_53[0][13] , \_zy_simnet_tvar_53[0].label[4] );
tran (\_zy_simnet_tvar_53[0][12] , \_zy_simnet_tvar_53[0].label[3] );
tran (\_zy_simnet_tvar_53[0][11] , \_zy_simnet_tvar_53[0].label[2] );
tran (\_zy_simnet_tvar_53[0][10] , \_zy_simnet_tvar_53[0].label[1] );
tran (\_zy_simnet_tvar_53[0][9] , \_zy_simnet_tvar_53[0].label[0] );
tran (\_zy_simnet_tvar_53[0][8] , \_zy_simnet_tvar_53[0].delimiter_valid[0] );
tran (\_zy_simnet_tvar_53[0][7] , \_zy_simnet_tvar_53[0].delimiter[7] );
tran (\_zy_simnet_tvar_53[0][6] , \_zy_simnet_tvar_53[0].delimiter[6] );
tran (\_zy_simnet_tvar_53[0][5] , \_zy_simnet_tvar_53[0].delimiter[5] );
tran (\_zy_simnet_tvar_53[0][4] , \_zy_simnet_tvar_53[0].delimiter[4] );
tran (\_zy_simnet_tvar_53[0][3] , \_zy_simnet_tvar_53[0].delimiter[3] );
tran (\_zy_simnet_tvar_53[0][2] , \_zy_simnet_tvar_53[0].delimiter[2] );
tran (\_zy_simnet_tvar_53[0][1] , \_zy_simnet_tvar_53[0].delimiter[1] );
tran (\_zy_simnet_tvar_53[0][0] , \_zy_simnet_tvar_53[0].delimiter[0] );
tran (\sa_ctrl[31][31] , \sa_ctrl[31].r.part0[31] );
tran (\sa_ctrl[31][31] , \sa_ctrl[31].f.spare[26] );
tran (\sa_ctrl[31][30] , \sa_ctrl[31].r.part0[30] );
tran (\sa_ctrl[31][30] , \sa_ctrl[31].f.spare[25] );
tran (\sa_ctrl[31][29] , \sa_ctrl[31].r.part0[29] );
tran (\sa_ctrl[31][29] , \sa_ctrl[31].f.spare[24] );
tran (\sa_ctrl[31][28] , \sa_ctrl[31].r.part0[28] );
tran (\sa_ctrl[31][28] , \sa_ctrl[31].f.spare[23] );
tran (\sa_ctrl[31][27] , \sa_ctrl[31].r.part0[27] );
tran (\sa_ctrl[31][27] , \sa_ctrl[31].f.spare[22] );
tran (\sa_ctrl[31][26] , \sa_ctrl[31].r.part0[26] );
tran (\sa_ctrl[31][26] , \sa_ctrl[31].f.spare[21] );
tran (\sa_ctrl[31][25] , \sa_ctrl[31].r.part0[25] );
tran (\sa_ctrl[31][25] , \sa_ctrl[31].f.spare[20] );
tran (\sa_ctrl[31][24] , \sa_ctrl[31].r.part0[24] );
tran (\sa_ctrl[31][24] , \sa_ctrl[31].f.spare[19] );
tran (\sa_ctrl[31][23] , \sa_ctrl[31].r.part0[23] );
tran (\sa_ctrl[31][23] , \sa_ctrl[31].f.spare[18] );
tran (\sa_ctrl[31][22] , \sa_ctrl[31].r.part0[22] );
tran (\sa_ctrl[31][22] , \sa_ctrl[31].f.spare[17] );
tran (\sa_ctrl[31][21] , \sa_ctrl[31].r.part0[21] );
tran (\sa_ctrl[31][21] , \sa_ctrl[31].f.spare[16] );
tran (\sa_ctrl[31][20] , \sa_ctrl[31].r.part0[20] );
tran (\sa_ctrl[31][20] , \sa_ctrl[31].f.spare[15] );
tran (\sa_ctrl[31][19] , \sa_ctrl[31].r.part0[19] );
tran (\sa_ctrl[31][19] , \sa_ctrl[31].f.spare[14] );
tran (\sa_ctrl[31][18] , \sa_ctrl[31].r.part0[18] );
tran (\sa_ctrl[31][18] , \sa_ctrl[31].f.spare[13] );
tran (\sa_ctrl[31][17] , \sa_ctrl[31].r.part0[17] );
tran (\sa_ctrl[31][17] , \sa_ctrl[31].f.spare[12] );
tran (\sa_ctrl[31][16] , \sa_ctrl[31].r.part0[16] );
tran (\sa_ctrl[31][16] , \sa_ctrl[31].f.spare[11] );
tran (\sa_ctrl[31][15] , \sa_ctrl[31].r.part0[15] );
tran (\sa_ctrl[31][15] , \sa_ctrl[31].f.spare[10] );
tran (\sa_ctrl[31][14] , \sa_ctrl[31].r.part0[14] );
tran (\sa_ctrl[31][14] , \sa_ctrl[31].f.spare[9] );
tran (\sa_ctrl[31][13] , \sa_ctrl[31].r.part0[13] );
tran (\sa_ctrl[31][13] , \sa_ctrl[31].f.spare[8] );
tran (\sa_ctrl[31][12] , \sa_ctrl[31].r.part0[12] );
tran (\sa_ctrl[31][12] , \sa_ctrl[31].f.spare[7] );
tran (\sa_ctrl[31][11] , \sa_ctrl[31].r.part0[11] );
tran (\sa_ctrl[31][11] , \sa_ctrl[31].f.spare[6] );
tran (\sa_ctrl[31][10] , \sa_ctrl[31].r.part0[10] );
tran (\sa_ctrl[31][10] , \sa_ctrl[31].f.spare[5] );
tran (\sa_ctrl[31][9] , \sa_ctrl[31].r.part0[9] );
tran (\sa_ctrl[31][9] , \sa_ctrl[31].f.spare[4] );
tran (\sa_ctrl[31][8] , \sa_ctrl[31].r.part0[8] );
tran (\sa_ctrl[31][8] , \sa_ctrl[31].f.spare[3] );
tran (\sa_ctrl[31][7] , \sa_ctrl[31].r.part0[7] );
tran (\sa_ctrl[31][7] , \sa_ctrl[31].f.spare[2] );
tran (\sa_ctrl[31][6] , \sa_ctrl[31].r.part0[6] );
tran (\sa_ctrl[31][6] , \sa_ctrl[31].f.spare[1] );
tran (\sa_ctrl[31][5] , \sa_ctrl[31].r.part0[5] );
tran (\sa_ctrl[31][5] , \sa_ctrl[31].f.spare[0] );
tran (\sa_ctrl[31][4] , \sa_ctrl[31].r.part0[4] );
tran (\sa_ctrl[31][4] , \sa_ctrl[31].f.sa_event_sel[4] );
tran (\sa_ctrl[31][3] , \sa_ctrl[31].r.part0[3] );
tran (\sa_ctrl[31][3] , \sa_ctrl[31].f.sa_event_sel[3] );
tran (\sa_ctrl[31][2] , \sa_ctrl[31].r.part0[2] );
tran (\sa_ctrl[31][2] , \sa_ctrl[31].f.sa_event_sel[2] );
tran (\sa_ctrl[31][1] , \sa_ctrl[31].r.part0[1] );
tran (\sa_ctrl[31][1] , \sa_ctrl[31].f.sa_event_sel[1] );
tran (\sa_ctrl[31][0] , \sa_ctrl[31].r.part0[0] );
tran (\sa_ctrl[31][0] , \sa_ctrl[31].f.sa_event_sel[0] );
tran (\sa_ctrl[30][31] , \sa_ctrl[30].r.part0[31] );
tran (\sa_ctrl[30][31] , \sa_ctrl[30].f.spare[26] );
tran (\sa_ctrl[30][30] , \sa_ctrl[30].r.part0[30] );
tran (\sa_ctrl[30][30] , \sa_ctrl[30].f.spare[25] );
tran (\sa_ctrl[30][29] , \sa_ctrl[30].r.part0[29] );
tran (\sa_ctrl[30][29] , \sa_ctrl[30].f.spare[24] );
tran (\sa_ctrl[30][28] , \sa_ctrl[30].r.part0[28] );
tran (\sa_ctrl[30][28] , \sa_ctrl[30].f.spare[23] );
tran (\sa_ctrl[30][27] , \sa_ctrl[30].r.part0[27] );
tran (\sa_ctrl[30][27] , \sa_ctrl[30].f.spare[22] );
tran (\sa_ctrl[30][26] , \sa_ctrl[30].r.part0[26] );
tran (\sa_ctrl[30][26] , \sa_ctrl[30].f.spare[21] );
tran (\sa_ctrl[30][25] , \sa_ctrl[30].r.part0[25] );
tran (\sa_ctrl[30][25] , \sa_ctrl[30].f.spare[20] );
tran (\sa_ctrl[30][24] , \sa_ctrl[30].r.part0[24] );
tran (\sa_ctrl[30][24] , \sa_ctrl[30].f.spare[19] );
tran (\sa_ctrl[30][23] , \sa_ctrl[30].r.part0[23] );
tran (\sa_ctrl[30][23] , \sa_ctrl[30].f.spare[18] );
tran (\sa_ctrl[30][22] , \sa_ctrl[30].r.part0[22] );
tran (\sa_ctrl[30][22] , \sa_ctrl[30].f.spare[17] );
tran (\sa_ctrl[30][21] , \sa_ctrl[30].r.part0[21] );
tran (\sa_ctrl[30][21] , \sa_ctrl[30].f.spare[16] );
tran (\sa_ctrl[30][20] , \sa_ctrl[30].r.part0[20] );
tran (\sa_ctrl[30][20] , \sa_ctrl[30].f.spare[15] );
tran (\sa_ctrl[30][19] , \sa_ctrl[30].r.part0[19] );
tran (\sa_ctrl[30][19] , \sa_ctrl[30].f.spare[14] );
tran (\sa_ctrl[30][18] , \sa_ctrl[30].r.part0[18] );
tran (\sa_ctrl[30][18] , \sa_ctrl[30].f.spare[13] );
tran (\sa_ctrl[30][17] , \sa_ctrl[30].r.part0[17] );
tran (\sa_ctrl[30][17] , \sa_ctrl[30].f.spare[12] );
tran (\sa_ctrl[30][16] , \sa_ctrl[30].r.part0[16] );
tran (\sa_ctrl[30][16] , \sa_ctrl[30].f.spare[11] );
tran (\sa_ctrl[30][15] , \sa_ctrl[30].r.part0[15] );
tran (\sa_ctrl[30][15] , \sa_ctrl[30].f.spare[10] );
tran (\sa_ctrl[30][14] , \sa_ctrl[30].r.part0[14] );
tran (\sa_ctrl[30][14] , \sa_ctrl[30].f.spare[9] );
tran (\sa_ctrl[30][13] , \sa_ctrl[30].r.part0[13] );
tran (\sa_ctrl[30][13] , \sa_ctrl[30].f.spare[8] );
tran (\sa_ctrl[30][12] , \sa_ctrl[30].r.part0[12] );
tran (\sa_ctrl[30][12] , \sa_ctrl[30].f.spare[7] );
tran (\sa_ctrl[30][11] , \sa_ctrl[30].r.part0[11] );
tran (\sa_ctrl[30][11] , \sa_ctrl[30].f.spare[6] );
tran (\sa_ctrl[30][10] , \sa_ctrl[30].r.part0[10] );
tran (\sa_ctrl[30][10] , \sa_ctrl[30].f.spare[5] );
tran (\sa_ctrl[30][9] , \sa_ctrl[30].r.part0[9] );
tran (\sa_ctrl[30][9] , \sa_ctrl[30].f.spare[4] );
tran (\sa_ctrl[30][8] , \sa_ctrl[30].r.part0[8] );
tran (\sa_ctrl[30][8] , \sa_ctrl[30].f.spare[3] );
tran (\sa_ctrl[30][7] , \sa_ctrl[30].r.part0[7] );
tran (\sa_ctrl[30][7] , \sa_ctrl[30].f.spare[2] );
tran (\sa_ctrl[30][6] , \sa_ctrl[30].r.part0[6] );
tran (\sa_ctrl[30][6] , \sa_ctrl[30].f.spare[1] );
tran (\sa_ctrl[30][5] , \sa_ctrl[30].r.part0[5] );
tran (\sa_ctrl[30][5] , \sa_ctrl[30].f.spare[0] );
tran (\sa_ctrl[30][4] , \sa_ctrl[30].r.part0[4] );
tran (\sa_ctrl[30][4] , \sa_ctrl[30].f.sa_event_sel[4] );
tran (\sa_ctrl[30][3] , \sa_ctrl[30].r.part0[3] );
tran (\sa_ctrl[30][3] , \sa_ctrl[30].f.sa_event_sel[3] );
tran (\sa_ctrl[30][2] , \sa_ctrl[30].r.part0[2] );
tran (\sa_ctrl[30][2] , \sa_ctrl[30].f.sa_event_sel[2] );
tran (\sa_ctrl[30][1] , \sa_ctrl[30].r.part0[1] );
tran (\sa_ctrl[30][1] , \sa_ctrl[30].f.sa_event_sel[1] );
tran (\sa_ctrl[30][0] , \sa_ctrl[30].r.part0[0] );
tran (\sa_ctrl[30][0] , \sa_ctrl[30].f.sa_event_sel[0] );
tran (\sa_ctrl[29][31] , \sa_ctrl[29].r.part0[31] );
tran (\sa_ctrl[29][31] , \sa_ctrl[29].f.spare[26] );
tran (\sa_ctrl[29][30] , \sa_ctrl[29].r.part0[30] );
tran (\sa_ctrl[29][30] , \sa_ctrl[29].f.spare[25] );
tran (\sa_ctrl[29][29] , \sa_ctrl[29].r.part0[29] );
tran (\sa_ctrl[29][29] , \sa_ctrl[29].f.spare[24] );
tran (\sa_ctrl[29][28] , \sa_ctrl[29].r.part0[28] );
tran (\sa_ctrl[29][28] , \sa_ctrl[29].f.spare[23] );
tran (\sa_ctrl[29][27] , \sa_ctrl[29].r.part0[27] );
tran (\sa_ctrl[29][27] , \sa_ctrl[29].f.spare[22] );
tran (\sa_ctrl[29][26] , \sa_ctrl[29].r.part0[26] );
tran (\sa_ctrl[29][26] , \sa_ctrl[29].f.spare[21] );
tran (\sa_ctrl[29][25] , \sa_ctrl[29].r.part0[25] );
tran (\sa_ctrl[29][25] , \sa_ctrl[29].f.spare[20] );
tran (\sa_ctrl[29][24] , \sa_ctrl[29].r.part0[24] );
tran (\sa_ctrl[29][24] , \sa_ctrl[29].f.spare[19] );
tran (\sa_ctrl[29][23] , \sa_ctrl[29].r.part0[23] );
tran (\sa_ctrl[29][23] , \sa_ctrl[29].f.spare[18] );
tran (\sa_ctrl[29][22] , \sa_ctrl[29].r.part0[22] );
tran (\sa_ctrl[29][22] , \sa_ctrl[29].f.spare[17] );
tran (\sa_ctrl[29][21] , \sa_ctrl[29].r.part0[21] );
tran (\sa_ctrl[29][21] , \sa_ctrl[29].f.spare[16] );
tran (\sa_ctrl[29][20] , \sa_ctrl[29].r.part0[20] );
tran (\sa_ctrl[29][20] , \sa_ctrl[29].f.spare[15] );
tran (\sa_ctrl[29][19] , \sa_ctrl[29].r.part0[19] );
tran (\sa_ctrl[29][19] , \sa_ctrl[29].f.spare[14] );
tran (\sa_ctrl[29][18] , \sa_ctrl[29].r.part0[18] );
tran (\sa_ctrl[29][18] , \sa_ctrl[29].f.spare[13] );
tran (\sa_ctrl[29][17] , \sa_ctrl[29].r.part0[17] );
tran (\sa_ctrl[29][17] , \sa_ctrl[29].f.spare[12] );
tran (\sa_ctrl[29][16] , \sa_ctrl[29].r.part0[16] );
tran (\sa_ctrl[29][16] , \sa_ctrl[29].f.spare[11] );
tran (\sa_ctrl[29][15] , \sa_ctrl[29].r.part0[15] );
tran (\sa_ctrl[29][15] , \sa_ctrl[29].f.spare[10] );
tran (\sa_ctrl[29][14] , \sa_ctrl[29].r.part0[14] );
tran (\sa_ctrl[29][14] , \sa_ctrl[29].f.spare[9] );
tran (\sa_ctrl[29][13] , \sa_ctrl[29].r.part0[13] );
tran (\sa_ctrl[29][13] , \sa_ctrl[29].f.spare[8] );
tran (\sa_ctrl[29][12] , \sa_ctrl[29].r.part0[12] );
tran (\sa_ctrl[29][12] , \sa_ctrl[29].f.spare[7] );
tran (\sa_ctrl[29][11] , \sa_ctrl[29].r.part0[11] );
tran (\sa_ctrl[29][11] , \sa_ctrl[29].f.spare[6] );
tran (\sa_ctrl[29][10] , \sa_ctrl[29].r.part0[10] );
tran (\sa_ctrl[29][10] , \sa_ctrl[29].f.spare[5] );
tran (\sa_ctrl[29][9] , \sa_ctrl[29].r.part0[9] );
tran (\sa_ctrl[29][9] , \sa_ctrl[29].f.spare[4] );
tran (\sa_ctrl[29][8] , \sa_ctrl[29].r.part0[8] );
tran (\sa_ctrl[29][8] , \sa_ctrl[29].f.spare[3] );
tran (\sa_ctrl[29][7] , \sa_ctrl[29].r.part0[7] );
tran (\sa_ctrl[29][7] , \sa_ctrl[29].f.spare[2] );
tran (\sa_ctrl[29][6] , \sa_ctrl[29].r.part0[6] );
tran (\sa_ctrl[29][6] , \sa_ctrl[29].f.spare[1] );
tran (\sa_ctrl[29][5] , \sa_ctrl[29].r.part0[5] );
tran (\sa_ctrl[29][5] , \sa_ctrl[29].f.spare[0] );
tran (\sa_ctrl[29][4] , \sa_ctrl[29].r.part0[4] );
tran (\sa_ctrl[29][4] , \sa_ctrl[29].f.sa_event_sel[4] );
tran (\sa_ctrl[29][3] , \sa_ctrl[29].r.part0[3] );
tran (\sa_ctrl[29][3] , \sa_ctrl[29].f.sa_event_sel[3] );
tran (\sa_ctrl[29][2] , \sa_ctrl[29].r.part0[2] );
tran (\sa_ctrl[29][2] , \sa_ctrl[29].f.sa_event_sel[2] );
tran (\sa_ctrl[29][1] , \sa_ctrl[29].r.part0[1] );
tran (\sa_ctrl[29][1] , \sa_ctrl[29].f.sa_event_sel[1] );
tran (\sa_ctrl[29][0] , \sa_ctrl[29].r.part0[0] );
tran (\sa_ctrl[29][0] , \sa_ctrl[29].f.sa_event_sel[0] );
tran (\sa_ctrl[28][31] , \sa_ctrl[28].r.part0[31] );
tran (\sa_ctrl[28][31] , \sa_ctrl[28].f.spare[26] );
tran (\sa_ctrl[28][30] , \sa_ctrl[28].r.part0[30] );
tran (\sa_ctrl[28][30] , \sa_ctrl[28].f.spare[25] );
tran (\sa_ctrl[28][29] , \sa_ctrl[28].r.part0[29] );
tran (\sa_ctrl[28][29] , \sa_ctrl[28].f.spare[24] );
tran (\sa_ctrl[28][28] , \sa_ctrl[28].r.part0[28] );
tran (\sa_ctrl[28][28] , \sa_ctrl[28].f.spare[23] );
tran (\sa_ctrl[28][27] , \sa_ctrl[28].r.part0[27] );
tran (\sa_ctrl[28][27] , \sa_ctrl[28].f.spare[22] );
tran (\sa_ctrl[28][26] , \sa_ctrl[28].r.part0[26] );
tran (\sa_ctrl[28][26] , \sa_ctrl[28].f.spare[21] );
tran (\sa_ctrl[28][25] , \sa_ctrl[28].r.part0[25] );
tran (\sa_ctrl[28][25] , \sa_ctrl[28].f.spare[20] );
tran (\sa_ctrl[28][24] , \sa_ctrl[28].r.part0[24] );
tran (\sa_ctrl[28][24] , \sa_ctrl[28].f.spare[19] );
tran (\sa_ctrl[28][23] , \sa_ctrl[28].r.part0[23] );
tran (\sa_ctrl[28][23] , \sa_ctrl[28].f.spare[18] );
tran (\sa_ctrl[28][22] , \sa_ctrl[28].r.part0[22] );
tran (\sa_ctrl[28][22] , \sa_ctrl[28].f.spare[17] );
tran (\sa_ctrl[28][21] , \sa_ctrl[28].r.part0[21] );
tran (\sa_ctrl[28][21] , \sa_ctrl[28].f.spare[16] );
tran (\sa_ctrl[28][20] , \sa_ctrl[28].r.part0[20] );
tran (\sa_ctrl[28][20] , \sa_ctrl[28].f.spare[15] );
tran (\sa_ctrl[28][19] , \sa_ctrl[28].r.part0[19] );
tran (\sa_ctrl[28][19] , \sa_ctrl[28].f.spare[14] );
tran (\sa_ctrl[28][18] , \sa_ctrl[28].r.part0[18] );
tran (\sa_ctrl[28][18] , \sa_ctrl[28].f.spare[13] );
tran (\sa_ctrl[28][17] , \sa_ctrl[28].r.part0[17] );
tran (\sa_ctrl[28][17] , \sa_ctrl[28].f.spare[12] );
tran (\sa_ctrl[28][16] , \sa_ctrl[28].r.part0[16] );
tran (\sa_ctrl[28][16] , \sa_ctrl[28].f.spare[11] );
tran (\sa_ctrl[28][15] , \sa_ctrl[28].r.part0[15] );
tran (\sa_ctrl[28][15] , \sa_ctrl[28].f.spare[10] );
tran (\sa_ctrl[28][14] , \sa_ctrl[28].r.part0[14] );
tran (\sa_ctrl[28][14] , \sa_ctrl[28].f.spare[9] );
tran (\sa_ctrl[28][13] , \sa_ctrl[28].r.part0[13] );
tran (\sa_ctrl[28][13] , \sa_ctrl[28].f.spare[8] );
tran (\sa_ctrl[28][12] , \sa_ctrl[28].r.part0[12] );
tran (\sa_ctrl[28][12] , \sa_ctrl[28].f.spare[7] );
tran (\sa_ctrl[28][11] , \sa_ctrl[28].r.part0[11] );
tran (\sa_ctrl[28][11] , \sa_ctrl[28].f.spare[6] );
tran (\sa_ctrl[28][10] , \sa_ctrl[28].r.part0[10] );
tran (\sa_ctrl[28][10] , \sa_ctrl[28].f.spare[5] );
tran (\sa_ctrl[28][9] , \sa_ctrl[28].r.part0[9] );
tran (\sa_ctrl[28][9] , \sa_ctrl[28].f.spare[4] );
tran (\sa_ctrl[28][8] , \sa_ctrl[28].r.part0[8] );
tran (\sa_ctrl[28][8] , \sa_ctrl[28].f.spare[3] );
tran (\sa_ctrl[28][7] , \sa_ctrl[28].r.part0[7] );
tran (\sa_ctrl[28][7] , \sa_ctrl[28].f.spare[2] );
tran (\sa_ctrl[28][6] , \sa_ctrl[28].r.part0[6] );
tran (\sa_ctrl[28][6] , \sa_ctrl[28].f.spare[1] );
tran (\sa_ctrl[28][5] , \sa_ctrl[28].r.part0[5] );
tran (\sa_ctrl[28][5] , \sa_ctrl[28].f.spare[0] );
tran (\sa_ctrl[28][4] , \sa_ctrl[28].r.part0[4] );
tran (\sa_ctrl[28][4] , \sa_ctrl[28].f.sa_event_sel[4] );
tran (\sa_ctrl[28][3] , \sa_ctrl[28].r.part0[3] );
tran (\sa_ctrl[28][3] , \sa_ctrl[28].f.sa_event_sel[3] );
tran (\sa_ctrl[28][2] , \sa_ctrl[28].r.part0[2] );
tran (\sa_ctrl[28][2] , \sa_ctrl[28].f.sa_event_sel[2] );
tran (\sa_ctrl[28][1] , \sa_ctrl[28].r.part0[1] );
tran (\sa_ctrl[28][1] , \sa_ctrl[28].f.sa_event_sel[1] );
tran (\sa_ctrl[28][0] , \sa_ctrl[28].r.part0[0] );
tran (\sa_ctrl[28][0] , \sa_ctrl[28].f.sa_event_sel[0] );
tran (\sa_ctrl[27][31] , \sa_ctrl[27].r.part0[31] );
tran (\sa_ctrl[27][31] , \sa_ctrl[27].f.spare[26] );
tran (\sa_ctrl[27][30] , \sa_ctrl[27].r.part0[30] );
tran (\sa_ctrl[27][30] , \sa_ctrl[27].f.spare[25] );
tran (\sa_ctrl[27][29] , \sa_ctrl[27].r.part0[29] );
tran (\sa_ctrl[27][29] , \sa_ctrl[27].f.spare[24] );
tran (\sa_ctrl[27][28] , \sa_ctrl[27].r.part0[28] );
tran (\sa_ctrl[27][28] , \sa_ctrl[27].f.spare[23] );
tran (\sa_ctrl[27][27] , \sa_ctrl[27].r.part0[27] );
tran (\sa_ctrl[27][27] , \sa_ctrl[27].f.spare[22] );
tran (\sa_ctrl[27][26] , \sa_ctrl[27].r.part0[26] );
tran (\sa_ctrl[27][26] , \sa_ctrl[27].f.spare[21] );
tran (\sa_ctrl[27][25] , \sa_ctrl[27].r.part0[25] );
tran (\sa_ctrl[27][25] , \sa_ctrl[27].f.spare[20] );
tran (\sa_ctrl[27][24] , \sa_ctrl[27].r.part0[24] );
tran (\sa_ctrl[27][24] , \sa_ctrl[27].f.spare[19] );
tran (\sa_ctrl[27][23] , \sa_ctrl[27].r.part0[23] );
tran (\sa_ctrl[27][23] , \sa_ctrl[27].f.spare[18] );
tran (\sa_ctrl[27][22] , \sa_ctrl[27].r.part0[22] );
tran (\sa_ctrl[27][22] , \sa_ctrl[27].f.spare[17] );
tran (\sa_ctrl[27][21] , \sa_ctrl[27].r.part0[21] );
tran (\sa_ctrl[27][21] , \sa_ctrl[27].f.spare[16] );
tran (\sa_ctrl[27][20] , \sa_ctrl[27].r.part0[20] );
tran (\sa_ctrl[27][20] , \sa_ctrl[27].f.spare[15] );
tran (\sa_ctrl[27][19] , \sa_ctrl[27].r.part0[19] );
tran (\sa_ctrl[27][19] , \sa_ctrl[27].f.spare[14] );
tran (\sa_ctrl[27][18] , \sa_ctrl[27].r.part0[18] );
tran (\sa_ctrl[27][18] , \sa_ctrl[27].f.spare[13] );
tran (\sa_ctrl[27][17] , \sa_ctrl[27].r.part0[17] );
tran (\sa_ctrl[27][17] , \sa_ctrl[27].f.spare[12] );
tran (\sa_ctrl[27][16] , \sa_ctrl[27].r.part0[16] );
tran (\sa_ctrl[27][16] , \sa_ctrl[27].f.spare[11] );
tran (\sa_ctrl[27][15] , \sa_ctrl[27].r.part0[15] );
tran (\sa_ctrl[27][15] , \sa_ctrl[27].f.spare[10] );
tran (\sa_ctrl[27][14] , \sa_ctrl[27].r.part0[14] );
tran (\sa_ctrl[27][14] , \sa_ctrl[27].f.spare[9] );
tran (\sa_ctrl[27][13] , \sa_ctrl[27].r.part0[13] );
tran (\sa_ctrl[27][13] , \sa_ctrl[27].f.spare[8] );
tran (\sa_ctrl[27][12] , \sa_ctrl[27].r.part0[12] );
tran (\sa_ctrl[27][12] , \sa_ctrl[27].f.spare[7] );
tran (\sa_ctrl[27][11] , \sa_ctrl[27].r.part0[11] );
tran (\sa_ctrl[27][11] , \sa_ctrl[27].f.spare[6] );
tran (\sa_ctrl[27][10] , \sa_ctrl[27].r.part0[10] );
tran (\sa_ctrl[27][10] , \sa_ctrl[27].f.spare[5] );
tran (\sa_ctrl[27][9] , \sa_ctrl[27].r.part0[9] );
tran (\sa_ctrl[27][9] , \sa_ctrl[27].f.spare[4] );
tran (\sa_ctrl[27][8] , \sa_ctrl[27].r.part0[8] );
tran (\sa_ctrl[27][8] , \sa_ctrl[27].f.spare[3] );
tran (\sa_ctrl[27][7] , \sa_ctrl[27].r.part0[7] );
tran (\sa_ctrl[27][7] , \sa_ctrl[27].f.spare[2] );
tran (\sa_ctrl[27][6] , \sa_ctrl[27].r.part0[6] );
tran (\sa_ctrl[27][6] , \sa_ctrl[27].f.spare[1] );
tran (\sa_ctrl[27][5] , \sa_ctrl[27].r.part0[5] );
tran (\sa_ctrl[27][5] , \sa_ctrl[27].f.spare[0] );
tran (\sa_ctrl[27][4] , \sa_ctrl[27].r.part0[4] );
tran (\sa_ctrl[27][4] , \sa_ctrl[27].f.sa_event_sel[4] );
tran (\sa_ctrl[27][3] , \sa_ctrl[27].r.part0[3] );
tran (\sa_ctrl[27][3] , \sa_ctrl[27].f.sa_event_sel[3] );
tran (\sa_ctrl[27][2] , \sa_ctrl[27].r.part0[2] );
tran (\sa_ctrl[27][2] , \sa_ctrl[27].f.sa_event_sel[2] );
tran (\sa_ctrl[27][1] , \sa_ctrl[27].r.part0[1] );
tran (\sa_ctrl[27][1] , \sa_ctrl[27].f.sa_event_sel[1] );
tran (\sa_ctrl[27][0] , \sa_ctrl[27].r.part0[0] );
tran (\sa_ctrl[27][0] , \sa_ctrl[27].f.sa_event_sel[0] );
tran (\sa_ctrl[26][31] , \sa_ctrl[26].r.part0[31] );
tran (\sa_ctrl[26][31] , \sa_ctrl[26].f.spare[26] );
tran (\sa_ctrl[26][30] , \sa_ctrl[26].r.part0[30] );
tran (\sa_ctrl[26][30] , \sa_ctrl[26].f.spare[25] );
tran (\sa_ctrl[26][29] , \sa_ctrl[26].r.part0[29] );
tran (\sa_ctrl[26][29] , \sa_ctrl[26].f.spare[24] );
tran (\sa_ctrl[26][28] , \sa_ctrl[26].r.part0[28] );
tran (\sa_ctrl[26][28] , \sa_ctrl[26].f.spare[23] );
tran (\sa_ctrl[26][27] , \sa_ctrl[26].r.part0[27] );
tran (\sa_ctrl[26][27] , \sa_ctrl[26].f.spare[22] );
tran (\sa_ctrl[26][26] , \sa_ctrl[26].r.part0[26] );
tran (\sa_ctrl[26][26] , \sa_ctrl[26].f.spare[21] );
tran (\sa_ctrl[26][25] , \sa_ctrl[26].r.part0[25] );
tran (\sa_ctrl[26][25] , \sa_ctrl[26].f.spare[20] );
tran (\sa_ctrl[26][24] , \sa_ctrl[26].r.part0[24] );
tran (\sa_ctrl[26][24] , \sa_ctrl[26].f.spare[19] );
tran (\sa_ctrl[26][23] , \sa_ctrl[26].r.part0[23] );
tran (\sa_ctrl[26][23] , \sa_ctrl[26].f.spare[18] );
tran (\sa_ctrl[26][22] , \sa_ctrl[26].r.part0[22] );
tran (\sa_ctrl[26][22] , \sa_ctrl[26].f.spare[17] );
tran (\sa_ctrl[26][21] , \sa_ctrl[26].r.part0[21] );
tran (\sa_ctrl[26][21] , \sa_ctrl[26].f.spare[16] );
tran (\sa_ctrl[26][20] , \sa_ctrl[26].r.part0[20] );
tran (\sa_ctrl[26][20] , \sa_ctrl[26].f.spare[15] );
tran (\sa_ctrl[26][19] , \sa_ctrl[26].r.part0[19] );
tran (\sa_ctrl[26][19] , \sa_ctrl[26].f.spare[14] );
tran (\sa_ctrl[26][18] , \sa_ctrl[26].r.part0[18] );
tran (\sa_ctrl[26][18] , \sa_ctrl[26].f.spare[13] );
tran (\sa_ctrl[26][17] , \sa_ctrl[26].r.part0[17] );
tran (\sa_ctrl[26][17] , \sa_ctrl[26].f.spare[12] );
tran (\sa_ctrl[26][16] , \sa_ctrl[26].r.part0[16] );
tran (\sa_ctrl[26][16] , \sa_ctrl[26].f.spare[11] );
tran (\sa_ctrl[26][15] , \sa_ctrl[26].r.part0[15] );
tran (\sa_ctrl[26][15] , \sa_ctrl[26].f.spare[10] );
tran (\sa_ctrl[26][14] , \sa_ctrl[26].r.part0[14] );
tran (\sa_ctrl[26][14] , \sa_ctrl[26].f.spare[9] );
tran (\sa_ctrl[26][13] , \sa_ctrl[26].r.part0[13] );
tran (\sa_ctrl[26][13] , \sa_ctrl[26].f.spare[8] );
tran (\sa_ctrl[26][12] , \sa_ctrl[26].r.part0[12] );
tran (\sa_ctrl[26][12] , \sa_ctrl[26].f.spare[7] );
tran (\sa_ctrl[26][11] , \sa_ctrl[26].r.part0[11] );
tran (\sa_ctrl[26][11] , \sa_ctrl[26].f.spare[6] );
tran (\sa_ctrl[26][10] , \sa_ctrl[26].r.part0[10] );
tran (\sa_ctrl[26][10] , \sa_ctrl[26].f.spare[5] );
tran (\sa_ctrl[26][9] , \sa_ctrl[26].r.part0[9] );
tran (\sa_ctrl[26][9] , \sa_ctrl[26].f.spare[4] );
tran (\sa_ctrl[26][8] , \sa_ctrl[26].r.part0[8] );
tran (\sa_ctrl[26][8] , \sa_ctrl[26].f.spare[3] );
tran (\sa_ctrl[26][7] , \sa_ctrl[26].r.part0[7] );
tran (\sa_ctrl[26][7] , \sa_ctrl[26].f.spare[2] );
tran (\sa_ctrl[26][6] , \sa_ctrl[26].r.part0[6] );
tran (\sa_ctrl[26][6] , \sa_ctrl[26].f.spare[1] );
tran (\sa_ctrl[26][5] , \sa_ctrl[26].r.part0[5] );
tran (\sa_ctrl[26][5] , \sa_ctrl[26].f.spare[0] );
tran (\sa_ctrl[26][4] , \sa_ctrl[26].r.part0[4] );
tran (\sa_ctrl[26][4] , \sa_ctrl[26].f.sa_event_sel[4] );
tran (\sa_ctrl[26][3] , \sa_ctrl[26].r.part0[3] );
tran (\sa_ctrl[26][3] , \sa_ctrl[26].f.sa_event_sel[3] );
tran (\sa_ctrl[26][2] , \sa_ctrl[26].r.part0[2] );
tran (\sa_ctrl[26][2] , \sa_ctrl[26].f.sa_event_sel[2] );
tran (\sa_ctrl[26][1] , \sa_ctrl[26].r.part0[1] );
tran (\sa_ctrl[26][1] , \sa_ctrl[26].f.sa_event_sel[1] );
tran (\sa_ctrl[26][0] , \sa_ctrl[26].r.part0[0] );
tran (\sa_ctrl[26][0] , \sa_ctrl[26].f.sa_event_sel[0] );
tran (\sa_ctrl[25][31] , \sa_ctrl[25].r.part0[31] );
tran (\sa_ctrl[25][31] , \sa_ctrl[25].f.spare[26] );
tran (\sa_ctrl[25][30] , \sa_ctrl[25].r.part0[30] );
tran (\sa_ctrl[25][30] , \sa_ctrl[25].f.spare[25] );
tran (\sa_ctrl[25][29] , \sa_ctrl[25].r.part0[29] );
tran (\sa_ctrl[25][29] , \sa_ctrl[25].f.spare[24] );
tran (\sa_ctrl[25][28] , \sa_ctrl[25].r.part0[28] );
tran (\sa_ctrl[25][28] , \sa_ctrl[25].f.spare[23] );
tran (\sa_ctrl[25][27] , \sa_ctrl[25].r.part0[27] );
tran (\sa_ctrl[25][27] , \sa_ctrl[25].f.spare[22] );
tran (\sa_ctrl[25][26] , \sa_ctrl[25].r.part0[26] );
tran (\sa_ctrl[25][26] , \sa_ctrl[25].f.spare[21] );
tran (\sa_ctrl[25][25] , \sa_ctrl[25].r.part0[25] );
tran (\sa_ctrl[25][25] , \sa_ctrl[25].f.spare[20] );
tran (\sa_ctrl[25][24] , \sa_ctrl[25].r.part0[24] );
tran (\sa_ctrl[25][24] , \sa_ctrl[25].f.spare[19] );
tran (\sa_ctrl[25][23] , \sa_ctrl[25].r.part0[23] );
tran (\sa_ctrl[25][23] , \sa_ctrl[25].f.spare[18] );
tran (\sa_ctrl[25][22] , \sa_ctrl[25].r.part0[22] );
tran (\sa_ctrl[25][22] , \sa_ctrl[25].f.spare[17] );
tran (\sa_ctrl[25][21] , \sa_ctrl[25].r.part0[21] );
tran (\sa_ctrl[25][21] , \sa_ctrl[25].f.spare[16] );
tran (\sa_ctrl[25][20] , \sa_ctrl[25].r.part0[20] );
tran (\sa_ctrl[25][20] , \sa_ctrl[25].f.spare[15] );
tran (\sa_ctrl[25][19] , \sa_ctrl[25].r.part0[19] );
tran (\sa_ctrl[25][19] , \sa_ctrl[25].f.spare[14] );
tran (\sa_ctrl[25][18] , \sa_ctrl[25].r.part0[18] );
tran (\sa_ctrl[25][18] , \sa_ctrl[25].f.spare[13] );
tran (\sa_ctrl[25][17] , \sa_ctrl[25].r.part0[17] );
tran (\sa_ctrl[25][17] , \sa_ctrl[25].f.spare[12] );
tran (\sa_ctrl[25][16] , \sa_ctrl[25].r.part0[16] );
tran (\sa_ctrl[25][16] , \sa_ctrl[25].f.spare[11] );
tran (\sa_ctrl[25][15] , \sa_ctrl[25].r.part0[15] );
tran (\sa_ctrl[25][15] , \sa_ctrl[25].f.spare[10] );
tran (\sa_ctrl[25][14] , \sa_ctrl[25].r.part0[14] );
tran (\sa_ctrl[25][14] , \sa_ctrl[25].f.spare[9] );
tran (\sa_ctrl[25][13] , \sa_ctrl[25].r.part0[13] );
tran (\sa_ctrl[25][13] , \sa_ctrl[25].f.spare[8] );
tran (\sa_ctrl[25][12] , \sa_ctrl[25].r.part0[12] );
tran (\sa_ctrl[25][12] , \sa_ctrl[25].f.spare[7] );
tran (\sa_ctrl[25][11] , \sa_ctrl[25].r.part0[11] );
tran (\sa_ctrl[25][11] , \sa_ctrl[25].f.spare[6] );
tran (\sa_ctrl[25][10] , \sa_ctrl[25].r.part0[10] );
tran (\sa_ctrl[25][10] , \sa_ctrl[25].f.spare[5] );
tran (\sa_ctrl[25][9] , \sa_ctrl[25].r.part0[9] );
tran (\sa_ctrl[25][9] , \sa_ctrl[25].f.spare[4] );
tran (\sa_ctrl[25][8] , \sa_ctrl[25].r.part0[8] );
tran (\sa_ctrl[25][8] , \sa_ctrl[25].f.spare[3] );
tran (\sa_ctrl[25][7] , \sa_ctrl[25].r.part0[7] );
tran (\sa_ctrl[25][7] , \sa_ctrl[25].f.spare[2] );
tran (\sa_ctrl[25][6] , \sa_ctrl[25].r.part0[6] );
tran (\sa_ctrl[25][6] , \sa_ctrl[25].f.spare[1] );
tran (\sa_ctrl[25][5] , \sa_ctrl[25].r.part0[5] );
tran (\sa_ctrl[25][5] , \sa_ctrl[25].f.spare[0] );
tran (\sa_ctrl[25][4] , \sa_ctrl[25].r.part0[4] );
tran (\sa_ctrl[25][4] , \sa_ctrl[25].f.sa_event_sel[4] );
tran (\sa_ctrl[25][3] , \sa_ctrl[25].r.part0[3] );
tran (\sa_ctrl[25][3] , \sa_ctrl[25].f.sa_event_sel[3] );
tran (\sa_ctrl[25][2] , \sa_ctrl[25].r.part0[2] );
tran (\sa_ctrl[25][2] , \sa_ctrl[25].f.sa_event_sel[2] );
tran (\sa_ctrl[25][1] , \sa_ctrl[25].r.part0[1] );
tran (\sa_ctrl[25][1] , \sa_ctrl[25].f.sa_event_sel[1] );
tran (\sa_ctrl[25][0] , \sa_ctrl[25].r.part0[0] );
tran (\sa_ctrl[25][0] , \sa_ctrl[25].f.sa_event_sel[0] );
tran (\sa_ctrl[24][31] , \sa_ctrl[24].r.part0[31] );
tran (\sa_ctrl[24][31] , \sa_ctrl[24].f.spare[26] );
tran (\sa_ctrl[24][30] , \sa_ctrl[24].r.part0[30] );
tran (\sa_ctrl[24][30] , \sa_ctrl[24].f.spare[25] );
tran (\sa_ctrl[24][29] , \sa_ctrl[24].r.part0[29] );
tran (\sa_ctrl[24][29] , \sa_ctrl[24].f.spare[24] );
tran (\sa_ctrl[24][28] , \sa_ctrl[24].r.part0[28] );
tran (\sa_ctrl[24][28] , \sa_ctrl[24].f.spare[23] );
tran (\sa_ctrl[24][27] , \sa_ctrl[24].r.part0[27] );
tran (\sa_ctrl[24][27] , \sa_ctrl[24].f.spare[22] );
tran (\sa_ctrl[24][26] , \sa_ctrl[24].r.part0[26] );
tran (\sa_ctrl[24][26] , \sa_ctrl[24].f.spare[21] );
tran (\sa_ctrl[24][25] , \sa_ctrl[24].r.part0[25] );
tran (\sa_ctrl[24][25] , \sa_ctrl[24].f.spare[20] );
tran (\sa_ctrl[24][24] , \sa_ctrl[24].r.part0[24] );
tran (\sa_ctrl[24][24] , \sa_ctrl[24].f.spare[19] );
tran (\sa_ctrl[24][23] , \sa_ctrl[24].r.part0[23] );
tran (\sa_ctrl[24][23] , \sa_ctrl[24].f.spare[18] );
tran (\sa_ctrl[24][22] , \sa_ctrl[24].r.part0[22] );
tran (\sa_ctrl[24][22] , \sa_ctrl[24].f.spare[17] );
tran (\sa_ctrl[24][21] , \sa_ctrl[24].r.part0[21] );
tran (\sa_ctrl[24][21] , \sa_ctrl[24].f.spare[16] );
tran (\sa_ctrl[24][20] , \sa_ctrl[24].r.part0[20] );
tran (\sa_ctrl[24][20] , \sa_ctrl[24].f.spare[15] );
tran (\sa_ctrl[24][19] , \sa_ctrl[24].r.part0[19] );
tran (\sa_ctrl[24][19] , \sa_ctrl[24].f.spare[14] );
tran (\sa_ctrl[24][18] , \sa_ctrl[24].r.part0[18] );
tran (\sa_ctrl[24][18] , \sa_ctrl[24].f.spare[13] );
tran (\sa_ctrl[24][17] , \sa_ctrl[24].r.part0[17] );
tran (\sa_ctrl[24][17] , \sa_ctrl[24].f.spare[12] );
tran (\sa_ctrl[24][16] , \sa_ctrl[24].r.part0[16] );
tran (\sa_ctrl[24][16] , \sa_ctrl[24].f.spare[11] );
tran (\sa_ctrl[24][15] , \sa_ctrl[24].r.part0[15] );
tran (\sa_ctrl[24][15] , \sa_ctrl[24].f.spare[10] );
tran (\sa_ctrl[24][14] , \sa_ctrl[24].r.part0[14] );
tran (\sa_ctrl[24][14] , \sa_ctrl[24].f.spare[9] );
tran (\sa_ctrl[24][13] , \sa_ctrl[24].r.part0[13] );
tran (\sa_ctrl[24][13] , \sa_ctrl[24].f.spare[8] );
tran (\sa_ctrl[24][12] , \sa_ctrl[24].r.part0[12] );
tran (\sa_ctrl[24][12] , \sa_ctrl[24].f.spare[7] );
tran (\sa_ctrl[24][11] , \sa_ctrl[24].r.part0[11] );
tran (\sa_ctrl[24][11] , \sa_ctrl[24].f.spare[6] );
tran (\sa_ctrl[24][10] , \sa_ctrl[24].r.part0[10] );
tran (\sa_ctrl[24][10] , \sa_ctrl[24].f.spare[5] );
tran (\sa_ctrl[24][9] , \sa_ctrl[24].r.part0[9] );
tran (\sa_ctrl[24][9] , \sa_ctrl[24].f.spare[4] );
tran (\sa_ctrl[24][8] , \sa_ctrl[24].r.part0[8] );
tran (\sa_ctrl[24][8] , \sa_ctrl[24].f.spare[3] );
tran (\sa_ctrl[24][7] , \sa_ctrl[24].r.part0[7] );
tran (\sa_ctrl[24][7] , \sa_ctrl[24].f.spare[2] );
tran (\sa_ctrl[24][6] , \sa_ctrl[24].r.part0[6] );
tran (\sa_ctrl[24][6] , \sa_ctrl[24].f.spare[1] );
tran (\sa_ctrl[24][5] , \sa_ctrl[24].r.part0[5] );
tran (\sa_ctrl[24][5] , \sa_ctrl[24].f.spare[0] );
tran (\sa_ctrl[24][4] , \sa_ctrl[24].r.part0[4] );
tran (\sa_ctrl[24][4] , \sa_ctrl[24].f.sa_event_sel[4] );
tran (\sa_ctrl[24][3] , \sa_ctrl[24].r.part0[3] );
tran (\sa_ctrl[24][3] , \sa_ctrl[24].f.sa_event_sel[3] );
tran (\sa_ctrl[24][2] , \sa_ctrl[24].r.part0[2] );
tran (\sa_ctrl[24][2] , \sa_ctrl[24].f.sa_event_sel[2] );
tran (\sa_ctrl[24][1] , \sa_ctrl[24].r.part0[1] );
tran (\sa_ctrl[24][1] , \sa_ctrl[24].f.sa_event_sel[1] );
tran (\sa_ctrl[24][0] , \sa_ctrl[24].r.part0[0] );
tran (\sa_ctrl[24][0] , \sa_ctrl[24].f.sa_event_sel[0] );
tran (\sa_ctrl[23][31] , \sa_ctrl[23].r.part0[31] );
tran (\sa_ctrl[23][31] , \sa_ctrl[23].f.spare[26] );
tran (\sa_ctrl[23][30] , \sa_ctrl[23].r.part0[30] );
tran (\sa_ctrl[23][30] , \sa_ctrl[23].f.spare[25] );
tran (\sa_ctrl[23][29] , \sa_ctrl[23].r.part0[29] );
tran (\sa_ctrl[23][29] , \sa_ctrl[23].f.spare[24] );
tran (\sa_ctrl[23][28] , \sa_ctrl[23].r.part0[28] );
tran (\sa_ctrl[23][28] , \sa_ctrl[23].f.spare[23] );
tran (\sa_ctrl[23][27] , \sa_ctrl[23].r.part0[27] );
tran (\sa_ctrl[23][27] , \sa_ctrl[23].f.spare[22] );
tran (\sa_ctrl[23][26] , \sa_ctrl[23].r.part0[26] );
tran (\sa_ctrl[23][26] , \sa_ctrl[23].f.spare[21] );
tran (\sa_ctrl[23][25] , \sa_ctrl[23].r.part0[25] );
tran (\sa_ctrl[23][25] , \sa_ctrl[23].f.spare[20] );
tran (\sa_ctrl[23][24] , \sa_ctrl[23].r.part0[24] );
tran (\sa_ctrl[23][24] , \sa_ctrl[23].f.spare[19] );
tran (\sa_ctrl[23][23] , \sa_ctrl[23].r.part0[23] );
tran (\sa_ctrl[23][23] , \sa_ctrl[23].f.spare[18] );
tran (\sa_ctrl[23][22] , \sa_ctrl[23].r.part0[22] );
tran (\sa_ctrl[23][22] , \sa_ctrl[23].f.spare[17] );
tran (\sa_ctrl[23][21] , \sa_ctrl[23].r.part0[21] );
tran (\sa_ctrl[23][21] , \sa_ctrl[23].f.spare[16] );
tran (\sa_ctrl[23][20] , \sa_ctrl[23].r.part0[20] );
tran (\sa_ctrl[23][20] , \sa_ctrl[23].f.spare[15] );
tran (\sa_ctrl[23][19] , \sa_ctrl[23].r.part0[19] );
tran (\sa_ctrl[23][19] , \sa_ctrl[23].f.spare[14] );
tran (\sa_ctrl[23][18] , \sa_ctrl[23].r.part0[18] );
tran (\sa_ctrl[23][18] , \sa_ctrl[23].f.spare[13] );
tran (\sa_ctrl[23][17] , \sa_ctrl[23].r.part0[17] );
tran (\sa_ctrl[23][17] , \sa_ctrl[23].f.spare[12] );
tran (\sa_ctrl[23][16] , \sa_ctrl[23].r.part0[16] );
tran (\sa_ctrl[23][16] , \sa_ctrl[23].f.spare[11] );
tran (\sa_ctrl[23][15] , \sa_ctrl[23].r.part0[15] );
tran (\sa_ctrl[23][15] , \sa_ctrl[23].f.spare[10] );
tran (\sa_ctrl[23][14] , \sa_ctrl[23].r.part0[14] );
tran (\sa_ctrl[23][14] , \sa_ctrl[23].f.spare[9] );
tran (\sa_ctrl[23][13] , \sa_ctrl[23].r.part0[13] );
tran (\sa_ctrl[23][13] , \sa_ctrl[23].f.spare[8] );
tran (\sa_ctrl[23][12] , \sa_ctrl[23].r.part0[12] );
tran (\sa_ctrl[23][12] , \sa_ctrl[23].f.spare[7] );
tran (\sa_ctrl[23][11] , \sa_ctrl[23].r.part0[11] );
tran (\sa_ctrl[23][11] , \sa_ctrl[23].f.spare[6] );
tran (\sa_ctrl[23][10] , \sa_ctrl[23].r.part0[10] );
tran (\sa_ctrl[23][10] , \sa_ctrl[23].f.spare[5] );
tran (\sa_ctrl[23][9] , \sa_ctrl[23].r.part0[9] );
tran (\sa_ctrl[23][9] , \sa_ctrl[23].f.spare[4] );
tran (\sa_ctrl[23][8] , \sa_ctrl[23].r.part0[8] );
tran (\sa_ctrl[23][8] , \sa_ctrl[23].f.spare[3] );
tran (\sa_ctrl[23][7] , \sa_ctrl[23].r.part0[7] );
tran (\sa_ctrl[23][7] , \sa_ctrl[23].f.spare[2] );
tran (\sa_ctrl[23][6] , \sa_ctrl[23].r.part0[6] );
tran (\sa_ctrl[23][6] , \sa_ctrl[23].f.spare[1] );
tran (\sa_ctrl[23][5] , \sa_ctrl[23].r.part0[5] );
tran (\sa_ctrl[23][5] , \sa_ctrl[23].f.spare[0] );
tran (\sa_ctrl[23][4] , \sa_ctrl[23].r.part0[4] );
tran (\sa_ctrl[23][4] , \sa_ctrl[23].f.sa_event_sel[4] );
tran (\sa_ctrl[23][3] , \sa_ctrl[23].r.part0[3] );
tran (\sa_ctrl[23][3] , \sa_ctrl[23].f.sa_event_sel[3] );
tran (\sa_ctrl[23][2] , \sa_ctrl[23].r.part0[2] );
tran (\sa_ctrl[23][2] , \sa_ctrl[23].f.sa_event_sel[2] );
tran (\sa_ctrl[23][1] , \sa_ctrl[23].r.part0[1] );
tran (\sa_ctrl[23][1] , \sa_ctrl[23].f.sa_event_sel[1] );
tran (\sa_ctrl[23][0] , \sa_ctrl[23].r.part0[0] );
tran (\sa_ctrl[23][0] , \sa_ctrl[23].f.sa_event_sel[0] );
tran (\sa_ctrl[22][31] , \sa_ctrl[22].r.part0[31] );
tran (\sa_ctrl[22][31] , \sa_ctrl[22].f.spare[26] );
tran (\sa_ctrl[22][30] , \sa_ctrl[22].r.part0[30] );
tran (\sa_ctrl[22][30] , \sa_ctrl[22].f.spare[25] );
tran (\sa_ctrl[22][29] , \sa_ctrl[22].r.part0[29] );
tran (\sa_ctrl[22][29] , \sa_ctrl[22].f.spare[24] );
tran (\sa_ctrl[22][28] , \sa_ctrl[22].r.part0[28] );
tran (\sa_ctrl[22][28] , \sa_ctrl[22].f.spare[23] );
tran (\sa_ctrl[22][27] , \sa_ctrl[22].r.part0[27] );
tran (\sa_ctrl[22][27] , \sa_ctrl[22].f.spare[22] );
tran (\sa_ctrl[22][26] , \sa_ctrl[22].r.part0[26] );
tran (\sa_ctrl[22][26] , \sa_ctrl[22].f.spare[21] );
tran (\sa_ctrl[22][25] , \sa_ctrl[22].r.part0[25] );
tran (\sa_ctrl[22][25] , \sa_ctrl[22].f.spare[20] );
tran (\sa_ctrl[22][24] , \sa_ctrl[22].r.part0[24] );
tran (\sa_ctrl[22][24] , \sa_ctrl[22].f.spare[19] );
tran (\sa_ctrl[22][23] , \sa_ctrl[22].r.part0[23] );
tran (\sa_ctrl[22][23] , \sa_ctrl[22].f.spare[18] );
tran (\sa_ctrl[22][22] , \sa_ctrl[22].r.part0[22] );
tran (\sa_ctrl[22][22] , \sa_ctrl[22].f.spare[17] );
tran (\sa_ctrl[22][21] , \sa_ctrl[22].r.part0[21] );
tran (\sa_ctrl[22][21] , \sa_ctrl[22].f.spare[16] );
tran (\sa_ctrl[22][20] , \sa_ctrl[22].r.part0[20] );
tran (\sa_ctrl[22][20] , \sa_ctrl[22].f.spare[15] );
tran (\sa_ctrl[22][19] , \sa_ctrl[22].r.part0[19] );
tran (\sa_ctrl[22][19] , \sa_ctrl[22].f.spare[14] );
tran (\sa_ctrl[22][18] , \sa_ctrl[22].r.part0[18] );
tran (\sa_ctrl[22][18] , \sa_ctrl[22].f.spare[13] );
tran (\sa_ctrl[22][17] , \sa_ctrl[22].r.part0[17] );
tran (\sa_ctrl[22][17] , \sa_ctrl[22].f.spare[12] );
tran (\sa_ctrl[22][16] , \sa_ctrl[22].r.part0[16] );
tran (\sa_ctrl[22][16] , \sa_ctrl[22].f.spare[11] );
tran (\sa_ctrl[22][15] , \sa_ctrl[22].r.part0[15] );
tran (\sa_ctrl[22][15] , \sa_ctrl[22].f.spare[10] );
tran (\sa_ctrl[22][14] , \sa_ctrl[22].r.part0[14] );
tran (\sa_ctrl[22][14] , \sa_ctrl[22].f.spare[9] );
tran (\sa_ctrl[22][13] , \sa_ctrl[22].r.part0[13] );
tran (\sa_ctrl[22][13] , \sa_ctrl[22].f.spare[8] );
tran (\sa_ctrl[22][12] , \sa_ctrl[22].r.part0[12] );
tran (\sa_ctrl[22][12] , \sa_ctrl[22].f.spare[7] );
tran (\sa_ctrl[22][11] , \sa_ctrl[22].r.part0[11] );
tran (\sa_ctrl[22][11] , \sa_ctrl[22].f.spare[6] );
tran (\sa_ctrl[22][10] , \sa_ctrl[22].r.part0[10] );
tran (\sa_ctrl[22][10] , \sa_ctrl[22].f.spare[5] );
tran (\sa_ctrl[22][9] , \sa_ctrl[22].r.part0[9] );
tran (\sa_ctrl[22][9] , \sa_ctrl[22].f.spare[4] );
tran (\sa_ctrl[22][8] , \sa_ctrl[22].r.part0[8] );
tran (\sa_ctrl[22][8] , \sa_ctrl[22].f.spare[3] );
tran (\sa_ctrl[22][7] , \sa_ctrl[22].r.part0[7] );
tran (\sa_ctrl[22][7] , \sa_ctrl[22].f.spare[2] );
tran (\sa_ctrl[22][6] , \sa_ctrl[22].r.part0[6] );
tran (\sa_ctrl[22][6] , \sa_ctrl[22].f.spare[1] );
tran (\sa_ctrl[22][5] , \sa_ctrl[22].r.part0[5] );
tran (\sa_ctrl[22][5] , \sa_ctrl[22].f.spare[0] );
tran (\sa_ctrl[22][4] , \sa_ctrl[22].r.part0[4] );
tran (\sa_ctrl[22][4] , \sa_ctrl[22].f.sa_event_sel[4] );
tran (\sa_ctrl[22][3] , \sa_ctrl[22].r.part0[3] );
tran (\sa_ctrl[22][3] , \sa_ctrl[22].f.sa_event_sel[3] );
tran (\sa_ctrl[22][2] , \sa_ctrl[22].r.part0[2] );
tran (\sa_ctrl[22][2] , \sa_ctrl[22].f.sa_event_sel[2] );
tran (\sa_ctrl[22][1] , \sa_ctrl[22].r.part0[1] );
tran (\sa_ctrl[22][1] , \sa_ctrl[22].f.sa_event_sel[1] );
tran (\sa_ctrl[22][0] , \sa_ctrl[22].r.part0[0] );
tran (\sa_ctrl[22][0] , \sa_ctrl[22].f.sa_event_sel[0] );
tran (\sa_ctrl[21][31] , \sa_ctrl[21].r.part0[31] );
tran (\sa_ctrl[21][31] , \sa_ctrl[21].f.spare[26] );
tran (\sa_ctrl[21][30] , \sa_ctrl[21].r.part0[30] );
tran (\sa_ctrl[21][30] , \sa_ctrl[21].f.spare[25] );
tran (\sa_ctrl[21][29] , \sa_ctrl[21].r.part0[29] );
tran (\sa_ctrl[21][29] , \sa_ctrl[21].f.spare[24] );
tran (\sa_ctrl[21][28] , \sa_ctrl[21].r.part0[28] );
tran (\sa_ctrl[21][28] , \sa_ctrl[21].f.spare[23] );
tran (\sa_ctrl[21][27] , \sa_ctrl[21].r.part0[27] );
tran (\sa_ctrl[21][27] , \sa_ctrl[21].f.spare[22] );
tran (\sa_ctrl[21][26] , \sa_ctrl[21].r.part0[26] );
tran (\sa_ctrl[21][26] , \sa_ctrl[21].f.spare[21] );
tran (\sa_ctrl[21][25] , \sa_ctrl[21].r.part0[25] );
tran (\sa_ctrl[21][25] , \sa_ctrl[21].f.spare[20] );
tran (\sa_ctrl[21][24] , \sa_ctrl[21].r.part0[24] );
tran (\sa_ctrl[21][24] , \sa_ctrl[21].f.spare[19] );
tran (\sa_ctrl[21][23] , \sa_ctrl[21].r.part0[23] );
tran (\sa_ctrl[21][23] , \sa_ctrl[21].f.spare[18] );
tran (\sa_ctrl[21][22] , \sa_ctrl[21].r.part0[22] );
tran (\sa_ctrl[21][22] , \sa_ctrl[21].f.spare[17] );
tran (\sa_ctrl[21][21] , \sa_ctrl[21].r.part0[21] );
tran (\sa_ctrl[21][21] , \sa_ctrl[21].f.spare[16] );
tran (\sa_ctrl[21][20] , \sa_ctrl[21].r.part0[20] );
tran (\sa_ctrl[21][20] , \sa_ctrl[21].f.spare[15] );
tran (\sa_ctrl[21][19] , \sa_ctrl[21].r.part0[19] );
tran (\sa_ctrl[21][19] , \sa_ctrl[21].f.spare[14] );
tran (\sa_ctrl[21][18] , \sa_ctrl[21].r.part0[18] );
tran (\sa_ctrl[21][18] , \sa_ctrl[21].f.spare[13] );
tran (\sa_ctrl[21][17] , \sa_ctrl[21].r.part0[17] );
tran (\sa_ctrl[21][17] , \sa_ctrl[21].f.spare[12] );
tran (\sa_ctrl[21][16] , \sa_ctrl[21].r.part0[16] );
tran (\sa_ctrl[21][16] , \sa_ctrl[21].f.spare[11] );
tran (\sa_ctrl[21][15] , \sa_ctrl[21].r.part0[15] );
tran (\sa_ctrl[21][15] , \sa_ctrl[21].f.spare[10] );
tran (\sa_ctrl[21][14] , \sa_ctrl[21].r.part0[14] );
tran (\sa_ctrl[21][14] , \sa_ctrl[21].f.spare[9] );
tran (\sa_ctrl[21][13] , \sa_ctrl[21].r.part0[13] );
tran (\sa_ctrl[21][13] , \sa_ctrl[21].f.spare[8] );
tran (\sa_ctrl[21][12] , \sa_ctrl[21].r.part0[12] );
tran (\sa_ctrl[21][12] , \sa_ctrl[21].f.spare[7] );
tran (\sa_ctrl[21][11] , \sa_ctrl[21].r.part0[11] );
tran (\sa_ctrl[21][11] , \sa_ctrl[21].f.spare[6] );
tran (\sa_ctrl[21][10] , \sa_ctrl[21].r.part0[10] );
tran (\sa_ctrl[21][10] , \sa_ctrl[21].f.spare[5] );
tran (\sa_ctrl[21][9] , \sa_ctrl[21].r.part0[9] );
tran (\sa_ctrl[21][9] , \sa_ctrl[21].f.spare[4] );
tran (\sa_ctrl[21][8] , \sa_ctrl[21].r.part0[8] );
tran (\sa_ctrl[21][8] , \sa_ctrl[21].f.spare[3] );
tran (\sa_ctrl[21][7] , \sa_ctrl[21].r.part0[7] );
tran (\sa_ctrl[21][7] , \sa_ctrl[21].f.spare[2] );
tran (\sa_ctrl[21][6] , \sa_ctrl[21].r.part0[6] );
tran (\sa_ctrl[21][6] , \sa_ctrl[21].f.spare[1] );
tran (\sa_ctrl[21][5] , \sa_ctrl[21].r.part0[5] );
tran (\sa_ctrl[21][5] , \sa_ctrl[21].f.spare[0] );
tran (\sa_ctrl[21][4] , \sa_ctrl[21].r.part0[4] );
tran (\sa_ctrl[21][4] , \sa_ctrl[21].f.sa_event_sel[4] );
tran (\sa_ctrl[21][3] , \sa_ctrl[21].r.part0[3] );
tran (\sa_ctrl[21][3] , \sa_ctrl[21].f.sa_event_sel[3] );
tran (\sa_ctrl[21][2] , \sa_ctrl[21].r.part0[2] );
tran (\sa_ctrl[21][2] , \sa_ctrl[21].f.sa_event_sel[2] );
tran (\sa_ctrl[21][1] , \sa_ctrl[21].r.part0[1] );
tran (\sa_ctrl[21][1] , \sa_ctrl[21].f.sa_event_sel[1] );
tran (\sa_ctrl[21][0] , \sa_ctrl[21].r.part0[0] );
tran (\sa_ctrl[21][0] , \sa_ctrl[21].f.sa_event_sel[0] );
tran (\sa_ctrl[20][31] , \sa_ctrl[20].r.part0[31] );
tran (\sa_ctrl[20][31] , \sa_ctrl[20].f.spare[26] );
tran (\sa_ctrl[20][30] , \sa_ctrl[20].r.part0[30] );
tran (\sa_ctrl[20][30] , \sa_ctrl[20].f.spare[25] );
tran (\sa_ctrl[20][29] , \sa_ctrl[20].r.part0[29] );
tran (\sa_ctrl[20][29] , \sa_ctrl[20].f.spare[24] );
tran (\sa_ctrl[20][28] , \sa_ctrl[20].r.part0[28] );
tran (\sa_ctrl[20][28] , \sa_ctrl[20].f.spare[23] );
tran (\sa_ctrl[20][27] , \sa_ctrl[20].r.part0[27] );
tran (\sa_ctrl[20][27] , \sa_ctrl[20].f.spare[22] );
tran (\sa_ctrl[20][26] , \sa_ctrl[20].r.part0[26] );
tran (\sa_ctrl[20][26] , \sa_ctrl[20].f.spare[21] );
tran (\sa_ctrl[20][25] , \sa_ctrl[20].r.part0[25] );
tran (\sa_ctrl[20][25] , \sa_ctrl[20].f.spare[20] );
tran (\sa_ctrl[20][24] , \sa_ctrl[20].r.part0[24] );
tran (\sa_ctrl[20][24] , \sa_ctrl[20].f.spare[19] );
tran (\sa_ctrl[20][23] , \sa_ctrl[20].r.part0[23] );
tran (\sa_ctrl[20][23] , \sa_ctrl[20].f.spare[18] );
tran (\sa_ctrl[20][22] , \sa_ctrl[20].r.part0[22] );
tran (\sa_ctrl[20][22] , \sa_ctrl[20].f.spare[17] );
tran (\sa_ctrl[20][21] , \sa_ctrl[20].r.part0[21] );
tran (\sa_ctrl[20][21] , \sa_ctrl[20].f.spare[16] );
tran (\sa_ctrl[20][20] , \sa_ctrl[20].r.part0[20] );
tran (\sa_ctrl[20][20] , \sa_ctrl[20].f.spare[15] );
tran (\sa_ctrl[20][19] , \sa_ctrl[20].r.part0[19] );
tran (\sa_ctrl[20][19] , \sa_ctrl[20].f.spare[14] );
tran (\sa_ctrl[20][18] , \sa_ctrl[20].r.part0[18] );
tran (\sa_ctrl[20][18] , \sa_ctrl[20].f.spare[13] );
tran (\sa_ctrl[20][17] , \sa_ctrl[20].r.part0[17] );
tran (\sa_ctrl[20][17] , \sa_ctrl[20].f.spare[12] );
tran (\sa_ctrl[20][16] , \sa_ctrl[20].r.part0[16] );
tran (\sa_ctrl[20][16] , \sa_ctrl[20].f.spare[11] );
tran (\sa_ctrl[20][15] , \sa_ctrl[20].r.part0[15] );
tran (\sa_ctrl[20][15] , \sa_ctrl[20].f.spare[10] );
tran (\sa_ctrl[20][14] , \sa_ctrl[20].r.part0[14] );
tran (\sa_ctrl[20][14] , \sa_ctrl[20].f.spare[9] );
tran (\sa_ctrl[20][13] , \sa_ctrl[20].r.part0[13] );
tran (\sa_ctrl[20][13] , \sa_ctrl[20].f.spare[8] );
tran (\sa_ctrl[20][12] , \sa_ctrl[20].r.part0[12] );
tran (\sa_ctrl[20][12] , \sa_ctrl[20].f.spare[7] );
tran (\sa_ctrl[20][11] , \sa_ctrl[20].r.part0[11] );
tran (\sa_ctrl[20][11] , \sa_ctrl[20].f.spare[6] );
tran (\sa_ctrl[20][10] , \sa_ctrl[20].r.part0[10] );
tran (\sa_ctrl[20][10] , \sa_ctrl[20].f.spare[5] );
tran (\sa_ctrl[20][9] , \sa_ctrl[20].r.part0[9] );
tran (\sa_ctrl[20][9] , \sa_ctrl[20].f.spare[4] );
tran (\sa_ctrl[20][8] , \sa_ctrl[20].r.part0[8] );
tran (\sa_ctrl[20][8] , \sa_ctrl[20].f.spare[3] );
tran (\sa_ctrl[20][7] , \sa_ctrl[20].r.part0[7] );
tran (\sa_ctrl[20][7] , \sa_ctrl[20].f.spare[2] );
tran (\sa_ctrl[20][6] , \sa_ctrl[20].r.part0[6] );
tran (\sa_ctrl[20][6] , \sa_ctrl[20].f.spare[1] );
tran (\sa_ctrl[20][5] , \sa_ctrl[20].r.part0[5] );
tran (\sa_ctrl[20][5] , \sa_ctrl[20].f.spare[0] );
tran (\sa_ctrl[20][4] , \sa_ctrl[20].r.part0[4] );
tran (\sa_ctrl[20][4] , \sa_ctrl[20].f.sa_event_sel[4] );
tran (\sa_ctrl[20][3] , \sa_ctrl[20].r.part0[3] );
tran (\sa_ctrl[20][3] , \sa_ctrl[20].f.sa_event_sel[3] );
tran (\sa_ctrl[20][2] , \sa_ctrl[20].r.part0[2] );
tran (\sa_ctrl[20][2] , \sa_ctrl[20].f.sa_event_sel[2] );
tran (\sa_ctrl[20][1] , \sa_ctrl[20].r.part0[1] );
tran (\sa_ctrl[20][1] , \sa_ctrl[20].f.sa_event_sel[1] );
tran (\sa_ctrl[20][0] , \sa_ctrl[20].r.part0[0] );
tran (\sa_ctrl[20][0] , \sa_ctrl[20].f.sa_event_sel[0] );
tran (\sa_ctrl[19][31] , \sa_ctrl[19].r.part0[31] );
tran (\sa_ctrl[19][31] , \sa_ctrl[19].f.spare[26] );
tran (\sa_ctrl[19][30] , \sa_ctrl[19].r.part0[30] );
tran (\sa_ctrl[19][30] , \sa_ctrl[19].f.spare[25] );
tran (\sa_ctrl[19][29] , \sa_ctrl[19].r.part0[29] );
tran (\sa_ctrl[19][29] , \sa_ctrl[19].f.spare[24] );
tran (\sa_ctrl[19][28] , \sa_ctrl[19].r.part0[28] );
tran (\sa_ctrl[19][28] , \sa_ctrl[19].f.spare[23] );
tran (\sa_ctrl[19][27] , \sa_ctrl[19].r.part0[27] );
tran (\sa_ctrl[19][27] , \sa_ctrl[19].f.spare[22] );
tran (\sa_ctrl[19][26] , \sa_ctrl[19].r.part0[26] );
tran (\sa_ctrl[19][26] , \sa_ctrl[19].f.spare[21] );
tran (\sa_ctrl[19][25] , \sa_ctrl[19].r.part0[25] );
tran (\sa_ctrl[19][25] , \sa_ctrl[19].f.spare[20] );
tran (\sa_ctrl[19][24] , \sa_ctrl[19].r.part0[24] );
tran (\sa_ctrl[19][24] , \sa_ctrl[19].f.spare[19] );
tran (\sa_ctrl[19][23] , \sa_ctrl[19].r.part0[23] );
tran (\sa_ctrl[19][23] , \sa_ctrl[19].f.spare[18] );
tran (\sa_ctrl[19][22] , \sa_ctrl[19].r.part0[22] );
tran (\sa_ctrl[19][22] , \sa_ctrl[19].f.spare[17] );
tran (\sa_ctrl[19][21] , \sa_ctrl[19].r.part0[21] );
tran (\sa_ctrl[19][21] , \sa_ctrl[19].f.spare[16] );
tran (\sa_ctrl[19][20] , \sa_ctrl[19].r.part0[20] );
tran (\sa_ctrl[19][20] , \sa_ctrl[19].f.spare[15] );
tran (\sa_ctrl[19][19] , \sa_ctrl[19].r.part0[19] );
tran (\sa_ctrl[19][19] , \sa_ctrl[19].f.spare[14] );
tran (\sa_ctrl[19][18] , \sa_ctrl[19].r.part0[18] );
tran (\sa_ctrl[19][18] , \sa_ctrl[19].f.spare[13] );
tran (\sa_ctrl[19][17] , \sa_ctrl[19].r.part0[17] );
tran (\sa_ctrl[19][17] , \sa_ctrl[19].f.spare[12] );
tran (\sa_ctrl[19][16] , \sa_ctrl[19].r.part0[16] );
tran (\sa_ctrl[19][16] , \sa_ctrl[19].f.spare[11] );
tran (\sa_ctrl[19][15] , \sa_ctrl[19].r.part0[15] );
tran (\sa_ctrl[19][15] , \sa_ctrl[19].f.spare[10] );
tran (\sa_ctrl[19][14] , \sa_ctrl[19].r.part0[14] );
tran (\sa_ctrl[19][14] , \sa_ctrl[19].f.spare[9] );
tran (\sa_ctrl[19][13] , \sa_ctrl[19].r.part0[13] );
tran (\sa_ctrl[19][13] , \sa_ctrl[19].f.spare[8] );
tran (\sa_ctrl[19][12] , \sa_ctrl[19].r.part0[12] );
tran (\sa_ctrl[19][12] , \sa_ctrl[19].f.spare[7] );
tran (\sa_ctrl[19][11] , \sa_ctrl[19].r.part0[11] );
tran (\sa_ctrl[19][11] , \sa_ctrl[19].f.spare[6] );
tran (\sa_ctrl[19][10] , \sa_ctrl[19].r.part0[10] );
tran (\sa_ctrl[19][10] , \sa_ctrl[19].f.spare[5] );
tran (\sa_ctrl[19][9] , \sa_ctrl[19].r.part0[9] );
tran (\sa_ctrl[19][9] , \sa_ctrl[19].f.spare[4] );
tran (\sa_ctrl[19][8] , \sa_ctrl[19].r.part0[8] );
tran (\sa_ctrl[19][8] , \sa_ctrl[19].f.spare[3] );
tran (\sa_ctrl[19][7] , \sa_ctrl[19].r.part0[7] );
tran (\sa_ctrl[19][7] , \sa_ctrl[19].f.spare[2] );
tran (\sa_ctrl[19][6] , \sa_ctrl[19].r.part0[6] );
tran (\sa_ctrl[19][6] , \sa_ctrl[19].f.spare[1] );
tran (\sa_ctrl[19][5] , \sa_ctrl[19].r.part0[5] );
tran (\sa_ctrl[19][5] , \sa_ctrl[19].f.spare[0] );
tran (\sa_ctrl[19][4] , \sa_ctrl[19].r.part0[4] );
tran (\sa_ctrl[19][4] , \sa_ctrl[19].f.sa_event_sel[4] );
tran (\sa_ctrl[19][3] , \sa_ctrl[19].r.part0[3] );
tran (\sa_ctrl[19][3] , \sa_ctrl[19].f.sa_event_sel[3] );
tran (\sa_ctrl[19][2] , \sa_ctrl[19].r.part0[2] );
tran (\sa_ctrl[19][2] , \sa_ctrl[19].f.sa_event_sel[2] );
tran (\sa_ctrl[19][1] , \sa_ctrl[19].r.part0[1] );
tran (\sa_ctrl[19][1] , \sa_ctrl[19].f.sa_event_sel[1] );
tran (\sa_ctrl[19][0] , \sa_ctrl[19].r.part0[0] );
tran (\sa_ctrl[19][0] , \sa_ctrl[19].f.sa_event_sel[0] );
tran (\sa_ctrl[18][31] , \sa_ctrl[18].r.part0[31] );
tran (\sa_ctrl[18][31] , \sa_ctrl[18].f.spare[26] );
tran (\sa_ctrl[18][30] , \sa_ctrl[18].r.part0[30] );
tran (\sa_ctrl[18][30] , \sa_ctrl[18].f.spare[25] );
tran (\sa_ctrl[18][29] , \sa_ctrl[18].r.part0[29] );
tran (\sa_ctrl[18][29] , \sa_ctrl[18].f.spare[24] );
tran (\sa_ctrl[18][28] , \sa_ctrl[18].r.part0[28] );
tran (\sa_ctrl[18][28] , \sa_ctrl[18].f.spare[23] );
tran (\sa_ctrl[18][27] , \sa_ctrl[18].r.part0[27] );
tran (\sa_ctrl[18][27] , \sa_ctrl[18].f.spare[22] );
tran (\sa_ctrl[18][26] , \sa_ctrl[18].r.part0[26] );
tran (\sa_ctrl[18][26] , \sa_ctrl[18].f.spare[21] );
tran (\sa_ctrl[18][25] , \sa_ctrl[18].r.part0[25] );
tran (\sa_ctrl[18][25] , \sa_ctrl[18].f.spare[20] );
tran (\sa_ctrl[18][24] , \sa_ctrl[18].r.part0[24] );
tran (\sa_ctrl[18][24] , \sa_ctrl[18].f.spare[19] );
tran (\sa_ctrl[18][23] , \sa_ctrl[18].r.part0[23] );
tran (\sa_ctrl[18][23] , \sa_ctrl[18].f.spare[18] );
tran (\sa_ctrl[18][22] , \sa_ctrl[18].r.part0[22] );
tran (\sa_ctrl[18][22] , \sa_ctrl[18].f.spare[17] );
tran (\sa_ctrl[18][21] , \sa_ctrl[18].r.part0[21] );
tran (\sa_ctrl[18][21] , \sa_ctrl[18].f.spare[16] );
tran (\sa_ctrl[18][20] , \sa_ctrl[18].r.part0[20] );
tran (\sa_ctrl[18][20] , \sa_ctrl[18].f.spare[15] );
tran (\sa_ctrl[18][19] , \sa_ctrl[18].r.part0[19] );
tran (\sa_ctrl[18][19] , \sa_ctrl[18].f.spare[14] );
tran (\sa_ctrl[18][18] , \sa_ctrl[18].r.part0[18] );
tran (\sa_ctrl[18][18] , \sa_ctrl[18].f.spare[13] );
tran (\sa_ctrl[18][17] , \sa_ctrl[18].r.part0[17] );
tran (\sa_ctrl[18][17] , \sa_ctrl[18].f.spare[12] );
tran (\sa_ctrl[18][16] , \sa_ctrl[18].r.part0[16] );
tran (\sa_ctrl[18][16] , \sa_ctrl[18].f.spare[11] );
tran (\sa_ctrl[18][15] , \sa_ctrl[18].r.part0[15] );
tran (\sa_ctrl[18][15] , \sa_ctrl[18].f.spare[10] );
tran (\sa_ctrl[18][14] , \sa_ctrl[18].r.part0[14] );
tran (\sa_ctrl[18][14] , \sa_ctrl[18].f.spare[9] );
tran (\sa_ctrl[18][13] , \sa_ctrl[18].r.part0[13] );
tran (\sa_ctrl[18][13] , \sa_ctrl[18].f.spare[8] );
tran (\sa_ctrl[18][12] , \sa_ctrl[18].r.part0[12] );
tran (\sa_ctrl[18][12] , \sa_ctrl[18].f.spare[7] );
tran (\sa_ctrl[18][11] , \sa_ctrl[18].r.part0[11] );
tran (\sa_ctrl[18][11] , \sa_ctrl[18].f.spare[6] );
tran (\sa_ctrl[18][10] , \sa_ctrl[18].r.part0[10] );
tran (\sa_ctrl[18][10] , \sa_ctrl[18].f.spare[5] );
tran (\sa_ctrl[18][9] , \sa_ctrl[18].r.part0[9] );
tran (\sa_ctrl[18][9] , \sa_ctrl[18].f.spare[4] );
tran (\sa_ctrl[18][8] , \sa_ctrl[18].r.part0[8] );
tran (\sa_ctrl[18][8] , \sa_ctrl[18].f.spare[3] );
tran (\sa_ctrl[18][7] , \sa_ctrl[18].r.part0[7] );
tran (\sa_ctrl[18][7] , \sa_ctrl[18].f.spare[2] );
tran (\sa_ctrl[18][6] , \sa_ctrl[18].r.part0[6] );
tran (\sa_ctrl[18][6] , \sa_ctrl[18].f.spare[1] );
tran (\sa_ctrl[18][5] , \sa_ctrl[18].r.part0[5] );
tran (\sa_ctrl[18][5] , \sa_ctrl[18].f.spare[0] );
tran (\sa_ctrl[18][4] , \sa_ctrl[18].r.part0[4] );
tran (\sa_ctrl[18][4] , \sa_ctrl[18].f.sa_event_sel[4] );
tran (\sa_ctrl[18][3] , \sa_ctrl[18].r.part0[3] );
tran (\sa_ctrl[18][3] , \sa_ctrl[18].f.sa_event_sel[3] );
tran (\sa_ctrl[18][2] , \sa_ctrl[18].r.part0[2] );
tran (\sa_ctrl[18][2] , \sa_ctrl[18].f.sa_event_sel[2] );
tran (\sa_ctrl[18][1] , \sa_ctrl[18].r.part0[1] );
tran (\sa_ctrl[18][1] , \sa_ctrl[18].f.sa_event_sel[1] );
tran (\sa_ctrl[18][0] , \sa_ctrl[18].r.part0[0] );
tran (\sa_ctrl[18][0] , \sa_ctrl[18].f.sa_event_sel[0] );
tran (\sa_ctrl[17][31] , \sa_ctrl[17].r.part0[31] );
tran (\sa_ctrl[17][31] , \sa_ctrl[17].f.spare[26] );
tran (\sa_ctrl[17][30] , \sa_ctrl[17].r.part0[30] );
tran (\sa_ctrl[17][30] , \sa_ctrl[17].f.spare[25] );
tran (\sa_ctrl[17][29] , \sa_ctrl[17].r.part0[29] );
tran (\sa_ctrl[17][29] , \sa_ctrl[17].f.spare[24] );
tran (\sa_ctrl[17][28] , \sa_ctrl[17].r.part0[28] );
tran (\sa_ctrl[17][28] , \sa_ctrl[17].f.spare[23] );
tran (\sa_ctrl[17][27] , \sa_ctrl[17].r.part0[27] );
tran (\sa_ctrl[17][27] , \sa_ctrl[17].f.spare[22] );
tran (\sa_ctrl[17][26] , \sa_ctrl[17].r.part0[26] );
tran (\sa_ctrl[17][26] , \sa_ctrl[17].f.spare[21] );
tran (\sa_ctrl[17][25] , \sa_ctrl[17].r.part0[25] );
tran (\sa_ctrl[17][25] , \sa_ctrl[17].f.spare[20] );
tran (\sa_ctrl[17][24] , \sa_ctrl[17].r.part0[24] );
tran (\sa_ctrl[17][24] , \sa_ctrl[17].f.spare[19] );
tran (\sa_ctrl[17][23] , \sa_ctrl[17].r.part0[23] );
tran (\sa_ctrl[17][23] , \sa_ctrl[17].f.spare[18] );
tran (\sa_ctrl[17][22] , \sa_ctrl[17].r.part0[22] );
tran (\sa_ctrl[17][22] , \sa_ctrl[17].f.spare[17] );
tran (\sa_ctrl[17][21] , \sa_ctrl[17].r.part0[21] );
tran (\sa_ctrl[17][21] , \sa_ctrl[17].f.spare[16] );
tran (\sa_ctrl[17][20] , \sa_ctrl[17].r.part0[20] );
tran (\sa_ctrl[17][20] , \sa_ctrl[17].f.spare[15] );
tran (\sa_ctrl[17][19] , \sa_ctrl[17].r.part0[19] );
tran (\sa_ctrl[17][19] , \sa_ctrl[17].f.spare[14] );
tran (\sa_ctrl[17][18] , \sa_ctrl[17].r.part0[18] );
tran (\sa_ctrl[17][18] , \sa_ctrl[17].f.spare[13] );
tran (\sa_ctrl[17][17] , \sa_ctrl[17].r.part0[17] );
tran (\sa_ctrl[17][17] , \sa_ctrl[17].f.spare[12] );
tran (\sa_ctrl[17][16] , \sa_ctrl[17].r.part0[16] );
tran (\sa_ctrl[17][16] , \sa_ctrl[17].f.spare[11] );
tran (\sa_ctrl[17][15] , \sa_ctrl[17].r.part0[15] );
tran (\sa_ctrl[17][15] , \sa_ctrl[17].f.spare[10] );
tran (\sa_ctrl[17][14] , \sa_ctrl[17].r.part0[14] );
tran (\sa_ctrl[17][14] , \sa_ctrl[17].f.spare[9] );
tran (\sa_ctrl[17][13] , \sa_ctrl[17].r.part0[13] );
tran (\sa_ctrl[17][13] , \sa_ctrl[17].f.spare[8] );
tran (\sa_ctrl[17][12] , \sa_ctrl[17].r.part0[12] );
tran (\sa_ctrl[17][12] , \sa_ctrl[17].f.spare[7] );
tran (\sa_ctrl[17][11] , \sa_ctrl[17].r.part0[11] );
tran (\sa_ctrl[17][11] , \sa_ctrl[17].f.spare[6] );
tran (\sa_ctrl[17][10] , \sa_ctrl[17].r.part0[10] );
tran (\sa_ctrl[17][10] , \sa_ctrl[17].f.spare[5] );
tran (\sa_ctrl[17][9] , \sa_ctrl[17].r.part0[9] );
tran (\sa_ctrl[17][9] , \sa_ctrl[17].f.spare[4] );
tran (\sa_ctrl[17][8] , \sa_ctrl[17].r.part0[8] );
tran (\sa_ctrl[17][8] , \sa_ctrl[17].f.spare[3] );
tran (\sa_ctrl[17][7] , \sa_ctrl[17].r.part0[7] );
tran (\sa_ctrl[17][7] , \sa_ctrl[17].f.spare[2] );
tran (\sa_ctrl[17][6] , \sa_ctrl[17].r.part0[6] );
tran (\sa_ctrl[17][6] , \sa_ctrl[17].f.spare[1] );
tran (\sa_ctrl[17][5] , \sa_ctrl[17].r.part0[5] );
tran (\sa_ctrl[17][5] , \sa_ctrl[17].f.spare[0] );
tran (\sa_ctrl[17][4] , \sa_ctrl[17].r.part0[4] );
tran (\sa_ctrl[17][4] , \sa_ctrl[17].f.sa_event_sel[4] );
tran (\sa_ctrl[17][3] , \sa_ctrl[17].r.part0[3] );
tran (\sa_ctrl[17][3] , \sa_ctrl[17].f.sa_event_sel[3] );
tran (\sa_ctrl[17][2] , \sa_ctrl[17].r.part0[2] );
tran (\sa_ctrl[17][2] , \sa_ctrl[17].f.sa_event_sel[2] );
tran (\sa_ctrl[17][1] , \sa_ctrl[17].r.part0[1] );
tran (\sa_ctrl[17][1] , \sa_ctrl[17].f.sa_event_sel[1] );
tran (\sa_ctrl[17][0] , \sa_ctrl[17].r.part0[0] );
tran (\sa_ctrl[17][0] , \sa_ctrl[17].f.sa_event_sel[0] );
tran (\sa_ctrl[16][31] , \sa_ctrl[16].r.part0[31] );
tran (\sa_ctrl[16][31] , \sa_ctrl[16].f.spare[26] );
tran (\sa_ctrl[16][30] , \sa_ctrl[16].r.part0[30] );
tran (\sa_ctrl[16][30] , \sa_ctrl[16].f.spare[25] );
tran (\sa_ctrl[16][29] , \sa_ctrl[16].r.part0[29] );
tran (\sa_ctrl[16][29] , \sa_ctrl[16].f.spare[24] );
tran (\sa_ctrl[16][28] , \sa_ctrl[16].r.part0[28] );
tran (\sa_ctrl[16][28] , \sa_ctrl[16].f.spare[23] );
tran (\sa_ctrl[16][27] , \sa_ctrl[16].r.part0[27] );
tran (\sa_ctrl[16][27] , \sa_ctrl[16].f.spare[22] );
tran (\sa_ctrl[16][26] , \sa_ctrl[16].r.part0[26] );
tran (\sa_ctrl[16][26] , \sa_ctrl[16].f.spare[21] );
tran (\sa_ctrl[16][25] , \sa_ctrl[16].r.part0[25] );
tran (\sa_ctrl[16][25] , \sa_ctrl[16].f.spare[20] );
tran (\sa_ctrl[16][24] , \sa_ctrl[16].r.part0[24] );
tran (\sa_ctrl[16][24] , \sa_ctrl[16].f.spare[19] );
tran (\sa_ctrl[16][23] , \sa_ctrl[16].r.part0[23] );
tran (\sa_ctrl[16][23] , \sa_ctrl[16].f.spare[18] );
tran (\sa_ctrl[16][22] , \sa_ctrl[16].r.part0[22] );
tran (\sa_ctrl[16][22] , \sa_ctrl[16].f.spare[17] );
tran (\sa_ctrl[16][21] , \sa_ctrl[16].r.part0[21] );
tran (\sa_ctrl[16][21] , \sa_ctrl[16].f.spare[16] );
tran (\sa_ctrl[16][20] , \sa_ctrl[16].r.part0[20] );
tran (\sa_ctrl[16][20] , \sa_ctrl[16].f.spare[15] );
tran (\sa_ctrl[16][19] , \sa_ctrl[16].r.part0[19] );
tran (\sa_ctrl[16][19] , \sa_ctrl[16].f.spare[14] );
tran (\sa_ctrl[16][18] , \sa_ctrl[16].r.part0[18] );
tran (\sa_ctrl[16][18] , \sa_ctrl[16].f.spare[13] );
tran (\sa_ctrl[16][17] , \sa_ctrl[16].r.part0[17] );
tran (\sa_ctrl[16][17] , \sa_ctrl[16].f.spare[12] );
tran (\sa_ctrl[16][16] , \sa_ctrl[16].r.part0[16] );
tran (\sa_ctrl[16][16] , \sa_ctrl[16].f.spare[11] );
tran (\sa_ctrl[16][15] , \sa_ctrl[16].r.part0[15] );
tran (\sa_ctrl[16][15] , \sa_ctrl[16].f.spare[10] );
tran (\sa_ctrl[16][14] , \sa_ctrl[16].r.part0[14] );
tran (\sa_ctrl[16][14] , \sa_ctrl[16].f.spare[9] );
tran (\sa_ctrl[16][13] , \sa_ctrl[16].r.part0[13] );
tran (\sa_ctrl[16][13] , \sa_ctrl[16].f.spare[8] );
tran (\sa_ctrl[16][12] , \sa_ctrl[16].r.part0[12] );
tran (\sa_ctrl[16][12] , \sa_ctrl[16].f.spare[7] );
tran (\sa_ctrl[16][11] , \sa_ctrl[16].r.part0[11] );
tran (\sa_ctrl[16][11] , \sa_ctrl[16].f.spare[6] );
tran (\sa_ctrl[16][10] , \sa_ctrl[16].r.part0[10] );
tran (\sa_ctrl[16][10] , \sa_ctrl[16].f.spare[5] );
tran (\sa_ctrl[16][9] , \sa_ctrl[16].r.part0[9] );
tran (\sa_ctrl[16][9] , \sa_ctrl[16].f.spare[4] );
tran (\sa_ctrl[16][8] , \sa_ctrl[16].r.part0[8] );
tran (\sa_ctrl[16][8] , \sa_ctrl[16].f.spare[3] );
tran (\sa_ctrl[16][7] , \sa_ctrl[16].r.part0[7] );
tran (\sa_ctrl[16][7] , \sa_ctrl[16].f.spare[2] );
tran (\sa_ctrl[16][6] , \sa_ctrl[16].r.part0[6] );
tran (\sa_ctrl[16][6] , \sa_ctrl[16].f.spare[1] );
tran (\sa_ctrl[16][5] , \sa_ctrl[16].r.part0[5] );
tran (\sa_ctrl[16][5] , \sa_ctrl[16].f.spare[0] );
tran (\sa_ctrl[16][4] , \sa_ctrl[16].r.part0[4] );
tran (\sa_ctrl[16][4] , \sa_ctrl[16].f.sa_event_sel[4] );
tran (\sa_ctrl[16][3] , \sa_ctrl[16].r.part0[3] );
tran (\sa_ctrl[16][3] , \sa_ctrl[16].f.sa_event_sel[3] );
tran (\sa_ctrl[16][2] , \sa_ctrl[16].r.part0[2] );
tran (\sa_ctrl[16][2] , \sa_ctrl[16].f.sa_event_sel[2] );
tran (\sa_ctrl[16][1] , \sa_ctrl[16].r.part0[1] );
tran (\sa_ctrl[16][1] , \sa_ctrl[16].f.sa_event_sel[1] );
tran (\sa_ctrl[16][0] , \sa_ctrl[16].r.part0[0] );
tran (\sa_ctrl[16][0] , \sa_ctrl[16].f.sa_event_sel[0] );
tran (\sa_ctrl[15][31] , \sa_ctrl[15].r.part0[31] );
tran (\sa_ctrl[15][31] , \sa_ctrl[15].f.spare[26] );
tran (\sa_ctrl[15][30] , \sa_ctrl[15].r.part0[30] );
tran (\sa_ctrl[15][30] , \sa_ctrl[15].f.spare[25] );
tran (\sa_ctrl[15][29] , \sa_ctrl[15].r.part0[29] );
tran (\sa_ctrl[15][29] , \sa_ctrl[15].f.spare[24] );
tran (\sa_ctrl[15][28] , \sa_ctrl[15].r.part0[28] );
tran (\sa_ctrl[15][28] , \sa_ctrl[15].f.spare[23] );
tran (\sa_ctrl[15][27] , \sa_ctrl[15].r.part0[27] );
tran (\sa_ctrl[15][27] , \sa_ctrl[15].f.spare[22] );
tran (\sa_ctrl[15][26] , \sa_ctrl[15].r.part0[26] );
tran (\sa_ctrl[15][26] , \sa_ctrl[15].f.spare[21] );
tran (\sa_ctrl[15][25] , \sa_ctrl[15].r.part0[25] );
tran (\sa_ctrl[15][25] , \sa_ctrl[15].f.spare[20] );
tran (\sa_ctrl[15][24] , \sa_ctrl[15].r.part0[24] );
tran (\sa_ctrl[15][24] , \sa_ctrl[15].f.spare[19] );
tran (\sa_ctrl[15][23] , \sa_ctrl[15].r.part0[23] );
tran (\sa_ctrl[15][23] , \sa_ctrl[15].f.spare[18] );
tran (\sa_ctrl[15][22] , \sa_ctrl[15].r.part0[22] );
tran (\sa_ctrl[15][22] , \sa_ctrl[15].f.spare[17] );
tran (\sa_ctrl[15][21] , \sa_ctrl[15].r.part0[21] );
tran (\sa_ctrl[15][21] , \sa_ctrl[15].f.spare[16] );
tran (\sa_ctrl[15][20] , \sa_ctrl[15].r.part0[20] );
tran (\sa_ctrl[15][20] , \sa_ctrl[15].f.spare[15] );
tran (\sa_ctrl[15][19] , \sa_ctrl[15].r.part0[19] );
tran (\sa_ctrl[15][19] , \sa_ctrl[15].f.spare[14] );
tran (\sa_ctrl[15][18] , \sa_ctrl[15].r.part0[18] );
tran (\sa_ctrl[15][18] , \sa_ctrl[15].f.spare[13] );
tran (\sa_ctrl[15][17] , \sa_ctrl[15].r.part0[17] );
tran (\sa_ctrl[15][17] , \sa_ctrl[15].f.spare[12] );
tran (\sa_ctrl[15][16] , \sa_ctrl[15].r.part0[16] );
tran (\sa_ctrl[15][16] , \sa_ctrl[15].f.spare[11] );
tran (\sa_ctrl[15][15] , \sa_ctrl[15].r.part0[15] );
tran (\sa_ctrl[15][15] , \sa_ctrl[15].f.spare[10] );
tran (\sa_ctrl[15][14] , \sa_ctrl[15].r.part0[14] );
tran (\sa_ctrl[15][14] , \sa_ctrl[15].f.spare[9] );
tran (\sa_ctrl[15][13] , \sa_ctrl[15].r.part0[13] );
tran (\sa_ctrl[15][13] , \sa_ctrl[15].f.spare[8] );
tran (\sa_ctrl[15][12] , \sa_ctrl[15].r.part0[12] );
tran (\sa_ctrl[15][12] , \sa_ctrl[15].f.spare[7] );
tran (\sa_ctrl[15][11] , \sa_ctrl[15].r.part0[11] );
tran (\sa_ctrl[15][11] , \sa_ctrl[15].f.spare[6] );
tran (\sa_ctrl[15][10] , \sa_ctrl[15].r.part0[10] );
tran (\sa_ctrl[15][10] , \sa_ctrl[15].f.spare[5] );
tran (\sa_ctrl[15][9] , \sa_ctrl[15].r.part0[9] );
tran (\sa_ctrl[15][9] , \sa_ctrl[15].f.spare[4] );
tran (\sa_ctrl[15][8] , \sa_ctrl[15].r.part0[8] );
tran (\sa_ctrl[15][8] , \sa_ctrl[15].f.spare[3] );
tran (\sa_ctrl[15][7] , \sa_ctrl[15].r.part0[7] );
tran (\sa_ctrl[15][7] , \sa_ctrl[15].f.spare[2] );
tran (\sa_ctrl[15][6] , \sa_ctrl[15].r.part0[6] );
tran (\sa_ctrl[15][6] , \sa_ctrl[15].f.spare[1] );
tran (\sa_ctrl[15][5] , \sa_ctrl[15].r.part0[5] );
tran (\sa_ctrl[15][5] , \sa_ctrl[15].f.spare[0] );
tran (\sa_ctrl[15][4] , \sa_ctrl[15].r.part0[4] );
tran (\sa_ctrl[15][4] , \sa_ctrl[15].f.sa_event_sel[4] );
tran (\sa_ctrl[15][3] , \sa_ctrl[15].r.part0[3] );
tran (\sa_ctrl[15][3] , \sa_ctrl[15].f.sa_event_sel[3] );
tran (\sa_ctrl[15][2] , \sa_ctrl[15].r.part0[2] );
tran (\sa_ctrl[15][2] , \sa_ctrl[15].f.sa_event_sel[2] );
tran (\sa_ctrl[15][1] , \sa_ctrl[15].r.part0[1] );
tran (\sa_ctrl[15][1] , \sa_ctrl[15].f.sa_event_sel[1] );
tran (\sa_ctrl[15][0] , \sa_ctrl[15].r.part0[0] );
tran (\sa_ctrl[15][0] , \sa_ctrl[15].f.sa_event_sel[0] );
tran (\sa_ctrl[14][31] , \sa_ctrl[14].r.part0[31] );
tran (\sa_ctrl[14][31] , \sa_ctrl[14].f.spare[26] );
tran (\sa_ctrl[14][30] , \sa_ctrl[14].r.part0[30] );
tran (\sa_ctrl[14][30] , \sa_ctrl[14].f.spare[25] );
tran (\sa_ctrl[14][29] , \sa_ctrl[14].r.part0[29] );
tran (\sa_ctrl[14][29] , \sa_ctrl[14].f.spare[24] );
tran (\sa_ctrl[14][28] , \sa_ctrl[14].r.part0[28] );
tran (\sa_ctrl[14][28] , \sa_ctrl[14].f.spare[23] );
tran (\sa_ctrl[14][27] , \sa_ctrl[14].r.part0[27] );
tran (\sa_ctrl[14][27] , \sa_ctrl[14].f.spare[22] );
tran (\sa_ctrl[14][26] , \sa_ctrl[14].r.part0[26] );
tran (\sa_ctrl[14][26] , \sa_ctrl[14].f.spare[21] );
tran (\sa_ctrl[14][25] , \sa_ctrl[14].r.part0[25] );
tran (\sa_ctrl[14][25] , \sa_ctrl[14].f.spare[20] );
tran (\sa_ctrl[14][24] , \sa_ctrl[14].r.part0[24] );
tran (\sa_ctrl[14][24] , \sa_ctrl[14].f.spare[19] );
tran (\sa_ctrl[14][23] , \sa_ctrl[14].r.part0[23] );
tran (\sa_ctrl[14][23] , \sa_ctrl[14].f.spare[18] );
tran (\sa_ctrl[14][22] , \sa_ctrl[14].r.part0[22] );
tran (\sa_ctrl[14][22] , \sa_ctrl[14].f.spare[17] );
tran (\sa_ctrl[14][21] , \sa_ctrl[14].r.part0[21] );
tran (\sa_ctrl[14][21] , \sa_ctrl[14].f.spare[16] );
tran (\sa_ctrl[14][20] , \sa_ctrl[14].r.part0[20] );
tran (\sa_ctrl[14][20] , \sa_ctrl[14].f.spare[15] );
tran (\sa_ctrl[14][19] , \sa_ctrl[14].r.part0[19] );
tran (\sa_ctrl[14][19] , \sa_ctrl[14].f.spare[14] );
tran (\sa_ctrl[14][18] , \sa_ctrl[14].r.part0[18] );
tran (\sa_ctrl[14][18] , \sa_ctrl[14].f.spare[13] );
tran (\sa_ctrl[14][17] , \sa_ctrl[14].r.part0[17] );
tran (\sa_ctrl[14][17] , \sa_ctrl[14].f.spare[12] );
tran (\sa_ctrl[14][16] , \sa_ctrl[14].r.part0[16] );
tran (\sa_ctrl[14][16] , \sa_ctrl[14].f.spare[11] );
tran (\sa_ctrl[14][15] , \sa_ctrl[14].r.part0[15] );
tran (\sa_ctrl[14][15] , \sa_ctrl[14].f.spare[10] );
tran (\sa_ctrl[14][14] , \sa_ctrl[14].r.part0[14] );
tran (\sa_ctrl[14][14] , \sa_ctrl[14].f.spare[9] );
tran (\sa_ctrl[14][13] , \sa_ctrl[14].r.part0[13] );
tran (\sa_ctrl[14][13] , \sa_ctrl[14].f.spare[8] );
tran (\sa_ctrl[14][12] , \sa_ctrl[14].r.part0[12] );
tran (\sa_ctrl[14][12] , \sa_ctrl[14].f.spare[7] );
tran (\sa_ctrl[14][11] , \sa_ctrl[14].r.part0[11] );
tran (\sa_ctrl[14][11] , \sa_ctrl[14].f.spare[6] );
tran (\sa_ctrl[14][10] , \sa_ctrl[14].r.part0[10] );
tran (\sa_ctrl[14][10] , \sa_ctrl[14].f.spare[5] );
tran (\sa_ctrl[14][9] , \sa_ctrl[14].r.part0[9] );
tran (\sa_ctrl[14][9] , \sa_ctrl[14].f.spare[4] );
tran (\sa_ctrl[14][8] , \sa_ctrl[14].r.part0[8] );
tran (\sa_ctrl[14][8] , \sa_ctrl[14].f.spare[3] );
tran (\sa_ctrl[14][7] , \sa_ctrl[14].r.part0[7] );
tran (\sa_ctrl[14][7] , \sa_ctrl[14].f.spare[2] );
tran (\sa_ctrl[14][6] , \sa_ctrl[14].r.part0[6] );
tran (\sa_ctrl[14][6] , \sa_ctrl[14].f.spare[1] );
tran (\sa_ctrl[14][5] , \sa_ctrl[14].r.part0[5] );
tran (\sa_ctrl[14][5] , \sa_ctrl[14].f.spare[0] );
tran (\sa_ctrl[14][4] , \sa_ctrl[14].r.part0[4] );
tran (\sa_ctrl[14][4] , \sa_ctrl[14].f.sa_event_sel[4] );
tran (\sa_ctrl[14][3] , \sa_ctrl[14].r.part0[3] );
tran (\sa_ctrl[14][3] , \sa_ctrl[14].f.sa_event_sel[3] );
tran (\sa_ctrl[14][2] , \sa_ctrl[14].r.part0[2] );
tran (\sa_ctrl[14][2] , \sa_ctrl[14].f.sa_event_sel[2] );
tran (\sa_ctrl[14][1] , \sa_ctrl[14].r.part0[1] );
tran (\sa_ctrl[14][1] , \sa_ctrl[14].f.sa_event_sel[1] );
tran (\sa_ctrl[14][0] , \sa_ctrl[14].r.part0[0] );
tran (\sa_ctrl[14][0] , \sa_ctrl[14].f.sa_event_sel[0] );
tran (\sa_ctrl[13][31] , \sa_ctrl[13].r.part0[31] );
tran (\sa_ctrl[13][31] , \sa_ctrl[13].f.spare[26] );
tran (\sa_ctrl[13][30] , \sa_ctrl[13].r.part0[30] );
tran (\sa_ctrl[13][30] , \sa_ctrl[13].f.spare[25] );
tran (\sa_ctrl[13][29] , \sa_ctrl[13].r.part0[29] );
tran (\sa_ctrl[13][29] , \sa_ctrl[13].f.spare[24] );
tran (\sa_ctrl[13][28] , \sa_ctrl[13].r.part0[28] );
tran (\sa_ctrl[13][28] , \sa_ctrl[13].f.spare[23] );
tran (\sa_ctrl[13][27] , \sa_ctrl[13].r.part0[27] );
tran (\sa_ctrl[13][27] , \sa_ctrl[13].f.spare[22] );
tran (\sa_ctrl[13][26] , \sa_ctrl[13].r.part0[26] );
tran (\sa_ctrl[13][26] , \sa_ctrl[13].f.spare[21] );
tran (\sa_ctrl[13][25] , \sa_ctrl[13].r.part0[25] );
tran (\sa_ctrl[13][25] , \sa_ctrl[13].f.spare[20] );
tran (\sa_ctrl[13][24] , \sa_ctrl[13].r.part0[24] );
tran (\sa_ctrl[13][24] , \sa_ctrl[13].f.spare[19] );
tran (\sa_ctrl[13][23] , \sa_ctrl[13].r.part0[23] );
tran (\sa_ctrl[13][23] , \sa_ctrl[13].f.spare[18] );
tran (\sa_ctrl[13][22] , \sa_ctrl[13].r.part0[22] );
tran (\sa_ctrl[13][22] , \sa_ctrl[13].f.spare[17] );
tran (\sa_ctrl[13][21] , \sa_ctrl[13].r.part0[21] );
tran (\sa_ctrl[13][21] , \sa_ctrl[13].f.spare[16] );
tran (\sa_ctrl[13][20] , \sa_ctrl[13].r.part0[20] );
tran (\sa_ctrl[13][20] , \sa_ctrl[13].f.spare[15] );
tran (\sa_ctrl[13][19] , \sa_ctrl[13].r.part0[19] );
tran (\sa_ctrl[13][19] , \sa_ctrl[13].f.spare[14] );
tran (\sa_ctrl[13][18] , \sa_ctrl[13].r.part0[18] );
tran (\sa_ctrl[13][18] , \sa_ctrl[13].f.spare[13] );
tran (\sa_ctrl[13][17] , \sa_ctrl[13].r.part0[17] );
tran (\sa_ctrl[13][17] , \sa_ctrl[13].f.spare[12] );
tran (\sa_ctrl[13][16] , \sa_ctrl[13].r.part0[16] );
tran (\sa_ctrl[13][16] , \sa_ctrl[13].f.spare[11] );
tran (\sa_ctrl[13][15] , \sa_ctrl[13].r.part0[15] );
tran (\sa_ctrl[13][15] , \sa_ctrl[13].f.spare[10] );
tran (\sa_ctrl[13][14] , \sa_ctrl[13].r.part0[14] );
tran (\sa_ctrl[13][14] , \sa_ctrl[13].f.spare[9] );
tran (\sa_ctrl[13][13] , \sa_ctrl[13].r.part0[13] );
tran (\sa_ctrl[13][13] , \sa_ctrl[13].f.spare[8] );
tran (\sa_ctrl[13][12] , \sa_ctrl[13].r.part0[12] );
tran (\sa_ctrl[13][12] , \sa_ctrl[13].f.spare[7] );
tran (\sa_ctrl[13][11] , \sa_ctrl[13].r.part0[11] );
tran (\sa_ctrl[13][11] , \sa_ctrl[13].f.spare[6] );
tran (\sa_ctrl[13][10] , \sa_ctrl[13].r.part0[10] );
tran (\sa_ctrl[13][10] , \sa_ctrl[13].f.spare[5] );
tran (\sa_ctrl[13][9] , \sa_ctrl[13].r.part0[9] );
tran (\sa_ctrl[13][9] , \sa_ctrl[13].f.spare[4] );
tran (\sa_ctrl[13][8] , \sa_ctrl[13].r.part0[8] );
tran (\sa_ctrl[13][8] , \sa_ctrl[13].f.spare[3] );
tran (\sa_ctrl[13][7] , \sa_ctrl[13].r.part0[7] );
tran (\sa_ctrl[13][7] , \sa_ctrl[13].f.spare[2] );
tran (\sa_ctrl[13][6] , \sa_ctrl[13].r.part0[6] );
tran (\sa_ctrl[13][6] , \sa_ctrl[13].f.spare[1] );
tran (\sa_ctrl[13][5] , \sa_ctrl[13].r.part0[5] );
tran (\sa_ctrl[13][5] , \sa_ctrl[13].f.spare[0] );
tran (\sa_ctrl[13][4] , \sa_ctrl[13].r.part0[4] );
tran (\sa_ctrl[13][4] , \sa_ctrl[13].f.sa_event_sel[4] );
tran (\sa_ctrl[13][3] , \sa_ctrl[13].r.part0[3] );
tran (\sa_ctrl[13][3] , \sa_ctrl[13].f.sa_event_sel[3] );
tran (\sa_ctrl[13][2] , \sa_ctrl[13].r.part0[2] );
tran (\sa_ctrl[13][2] , \sa_ctrl[13].f.sa_event_sel[2] );
tran (\sa_ctrl[13][1] , \sa_ctrl[13].r.part0[1] );
tran (\sa_ctrl[13][1] , \sa_ctrl[13].f.sa_event_sel[1] );
tran (\sa_ctrl[13][0] , \sa_ctrl[13].r.part0[0] );
tran (\sa_ctrl[13][0] , \sa_ctrl[13].f.sa_event_sel[0] );
tran (\sa_ctrl[12][31] , \sa_ctrl[12].r.part0[31] );
tran (\sa_ctrl[12][31] , \sa_ctrl[12].f.spare[26] );
tran (\sa_ctrl[12][30] , \sa_ctrl[12].r.part0[30] );
tran (\sa_ctrl[12][30] , \sa_ctrl[12].f.spare[25] );
tran (\sa_ctrl[12][29] , \sa_ctrl[12].r.part0[29] );
tran (\sa_ctrl[12][29] , \sa_ctrl[12].f.spare[24] );
tran (\sa_ctrl[12][28] , \sa_ctrl[12].r.part0[28] );
tran (\sa_ctrl[12][28] , \sa_ctrl[12].f.spare[23] );
tran (\sa_ctrl[12][27] , \sa_ctrl[12].r.part0[27] );
tran (\sa_ctrl[12][27] , \sa_ctrl[12].f.spare[22] );
tran (\sa_ctrl[12][26] , \sa_ctrl[12].r.part0[26] );
tran (\sa_ctrl[12][26] , \sa_ctrl[12].f.spare[21] );
tran (\sa_ctrl[12][25] , \sa_ctrl[12].r.part0[25] );
tran (\sa_ctrl[12][25] , \sa_ctrl[12].f.spare[20] );
tran (\sa_ctrl[12][24] , \sa_ctrl[12].r.part0[24] );
tran (\sa_ctrl[12][24] , \sa_ctrl[12].f.spare[19] );
tran (\sa_ctrl[12][23] , \sa_ctrl[12].r.part0[23] );
tran (\sa_ctrl[12][23] , \sa_ctrl[12].f.spare[18] );
tran (\sa_ctrl[12][22] , \sa_ctrl[12].r.part0[22] );
tran (\sa_ctrl[12][22] , \sa_ctrl[12].f.spare[17] );
tran (\sa_ctrl[12][21] , \sa_ctrl[12].r.part0[21] );
tran (\sa_ctrl[12][21] , \sa_ctrl[12].f.spare[16] );
tran (\sa_ctrl[12][20] , \sa_ctrl[12].r.part0[20] );
tran (\sa_ctrl[12][20] , \sa_ctrl[12].f.spare[15] );
tran (\sa_ctrl[12][19] , \sa_ctrl[12].r.part0[19] );
tran (\sa_ctrl[12][19] , \sa_ctrl[12].f.spare[14] );
tran (\sa_ctrl[12][18] , \sa_ctrl[12].r.part0[18] );
tran (\sa_ctrl[12][18] , \sa_ctrl[12].f.spare[13] );
tran (\sa_ctrl[12][17] , \sa_ctrl[12].r.part0[17] );
tran (\sa_ctrl[12][17] , \sa_ctrl[12].f.spare[12] );
tran (\sa_ctrl[12][16] , \sa_ctrl[12].r.part0[16] );
tran (\sa_ctrl[12][16] , \sa_ctrl[12].f.spare[11] );
tran (\sa_ctrl[12][15] , \sa_ctrl[12].r.part0[15] );
tran (\sa_ctrl[12][15] , \sa_ctrl[12].f.spare[10] );
tran (\sa_ctrl[12][14] , \sa_ctrl[12].r.part0[14] );
tran (\sa_ctrl[12][14] , \sa_ctrl[12].f.spare[9] );
tran (\sa_ctrl[12][13] , \sa_ctrl[12].r.part0[13] );
tran (\sa_ctrl[12][13] , \sa_ctrl[12].f.spare[8] );
tran (\sa_ctrl[12][12] , \sa_ctrl[12].r.part0[12] );
tran (\sa_ctrl[12][12] , \sa_ctrl[12].f.spare[7] );
tran (\sa_ctrl[12][11] , \sa_ctrl[12].r.part0[11] );
tran (\sa_ctrl[12][11] , \sa_ctrl[12].f.spare[6] );
tran (\sa_ctrl[12][10] , \sa_ctrl[12].r.part0[10] );
tran (\sa_ctrl[12][10] , \sa_ctrl[12].f.spare[5] );
tran (\sa_ctrl[12][9] , \sa_ctrl[12].r.part0[9] );
tran (\sa_ctrl[12][9] , \sa_ctrl[12].f.spare[4] );
tran (\sa_ctrl[12][8] , \sa_ctrl[12].r.part0[8] );
tran (\sa_ctrl[12][8] , \sa_ctrl[12].f.spare[3] );
tran (\sa_ctrl[12][7] , \sa_ctrl[12].r.part0[7] );
tran (\sa_ctrl[12][7] , \sa_ctrl[12].f.spare[2] );
tran (\sa_ctrl[12][6] , \sa_ctrl[12].r.part0[6] );
tran (\sa_ctrl[12][6] , \sa_ctrl[12].f.spare[1] );
tran (\sa_ctrl[12][5] , \sa_ctrl[12].r.part0[5] );
tran (\sa_ctrl[12][5] , \sa_ctrl[12].f.spare[0] );
tran (\sa_ctrl[12][4] , \sa_ctrl[12].r.part0[4] );
tran (\sa_ctrl[12][4] , \sa_ctrl[12].f.sa_event_sel[4] );
tran (\sa_ctrl[12][3] , \sa_ctrl[12].r.part0[3] );
tran (\sa_ctrl[12][3] , \sa_ctrl[12].f.sa_event_sel[3] );
tran (\sa_ctrl[12][2] , \sa_ctrl[12].r.part0[2] );
tran (\sa_ctrl[12][2] , \sa_ctrl[12].f.sa_event_sel[2] );
tran (\sa_ctrl[12][1] , \sa_ctrl[12].r.part0[1] );
tran (\sa_ctrl[12][1] , \sa_ctrl[12].f.sa_event_sel[1] );
tran (\sa_ctrl[12][0] , \sa_ctrl[12].r.part0[0] );
tran (\sa_ctrl[12][0] , \sa_ctrl[12].f.sa_event_sel[0] );
tran (\sa_ctrl[11][31] , \sa_ctrl[11].r.part0[31] );
tran (\sa_ctrl[11][31] , \sa_ctrl[11].f.spare[26] );
tran (\sa_ctrl[11][30] , \sa_ctrl[11].r.part0[30] );
tran (\sa_ctrl[11][30] , \sa_ctrl[11].f.spare[25] );
tran (\sa_ctrl[11][29] , \sa_ctrl[11].r.part0[29] );
tran (\sa_ctrl[11][29] , \sa_ctrl[11].f.spare[24] );
tran (\sa_ctrl[11][28] , \sa_ctrl[11].r.part0[28] );
tran (\sa_ctrl[11][28] , \sa_ctrl[11].f.spare[23] );
tran (\sa_ctrl[11][27] , \sa_ctrl[11].r.part0[27] );
tran (\sa_ctrl[11][27] , \sa_ctrl[11].f.spare[22] );
tran (\sa_ctrl[11][26] , \sa_ctrl[11].r.part0[26] );
tran (\sa_ctrl[11][26] , \sa_ctrl[11].f.spare[21] );
tran (\sa_ctrl[11][25] , \sa_ctrl[11].r.part0[25] );
tran (\sa_ctrl[11][25] , \sa_ctrl[11].f.spare[20] );
tran (\sa_ctrl[11][24] , \sa_ctrl[11].r.part0[24] );
tran (\sa_ctrl[11][24] , \sa_ctrl[11].f.spare[19] );
tran (\sa_ctrl[11][23] , \sa_ctrl[11].r.part0[23] );
tran (\sa_ctrl[11][23] , \sa_ctrl[11].f.spare[18] );
tran (\sa_ctrl[11][22] , \sa_ctrl[11].r.part0[22] );
tran (\sa_ctrl[11][22] , \sa_ctrl[11].f.spare[17] );
tran (\sa_ctrl[11][21] , \sa_ctrl[11].r.part0[21] );
tran (\sa_ctrl[11][21] , \sa_ctrl[11].f.spare[16] );
tran (\sa_ctrl[11][20] , \sa_ctrl[11].r.part0[20] );
tran (\sa_ctrl[11][20] , \sa_ctrl[11].f.spare[15] );
tran (\sa_ctrl[11][19] , \sa_ctrl[11].r.part0[19] );
tran (\sa_ctrl[11][19] , \sa_ctrl[11].f.spare[14] );
tran (\sa_ctrl[11][18] , \sa_ctrl[11].r.part0[18] );
tran (\sa_ctrl[11][18] , \sa_ctrl[11].f.spare[13] );
tran (\sa_ctrl[11][17] , \sa_ctrl[11].r.part0[17] );
tran (\sa_ctrl[11][17] , \sa_ctrl[11].f.spare[12] );
tran (\sa_ctrl[11][16] , \sa_ctrl[11].r.part0[16] );
tran (\sa_ctrl[11][16] , \sa_ctrl[11].f.spare[11] );
tran (\sa_ctrl[11][15] , \sa_ctrl[11].r.part0[15] );
tran (\sa_ctrl[11][15] , \sa_ctrl[11].f.spare[10] );
tran (\sa_ctrl[11][14] , \sa_ctrl[11].r.part0[14] );
tran (\sa_ctrl[11][14] , \sa_ctrl[11].f.spare[9] );
tran (\sa_ctrl[11][13] , \sa_ctrl[11].r.part0[13] );
tran (\sa_ctrl[11][13] , \sa_ctrl[11].f.spare[8] );
tran (\sa_ctrl[11][12] , \sa_ctrl[11].r.part0[12] );
tran (\sa_ctrl[11][12] , \sa_ctrl[11].f.spare[7] );
tran (\sa_ctrl[11][11] , \sa_ctrl[11].r.part0[11] );
tran (\sa_ctrl[11][11] , \sa_ctrl[11].f.spare[6] );
tran (\sa_ctrl[11][10] , \sa_ctrl[11].r.part0[10] );
tran (\sa_ctrl[11][10] , \sa_ctrl[11].f.spare[5] );
tran (\sa_ctrl[11][9] , \sa_ctrl[11].r.part0[9] );
tran (\sa_ctrl[11][9] , \sa_ctrl[11].f.spare[4] );
tran (\sa_ctrl[11][8] , \sa_ctrl[11].r.part0[8] );
tran (\sa_ctrl[11][8] , \sa_ctrl[11].f.spare[3] );
tran (\sa_ctrl[11][7] , \sa_ctrl[11].r.part0[7] );
tran (\sa_ctrl[11][7] , \sa_ctrl[11].f.spare[2] );
tran (\sa_ctrl[11][6] , \sa_ctrl[11].r.part0[6] );
tran (\sa_ctrl[11][6] , \sa_ctrl[11].f.spare[1] );
tran (\sa_ctrl[11][5] , \sa_ctrl[11].r.part0[5] );
tran (\sa_ctrl[11][5] , \sa_ctrl[11].f.spare[0] );
tran (\sa_ctrl[11][4] , \sa_ctrl[11].r.part0[4] );
tran (\sa_ctrl[11][4] , \sa_ctrl[11].f.sa_event_sel[4] );
tran (\sa_ctrl[11][3] , \sa_ctrl[11].r.part0[3] );
tran (\sa_ctrl[11][3] , \sa_ctrl[11].f.sa_event_sel[3] );
tran (\sa_ctrl[11][2] , \sa_ctrl[11].r.part0[2] );
tran (\sa_ctrl[11][2] , \sa_ctrl[11].f.sa_event_sel[2] );
tran (\sa_ctrl[11][1] , \sa_ctrl[11].r.part0[1] );
tran (\sa_ctrl[11][1] , \sa_ctrl[11].f.sa_event_sel[1] );
tran (\sa_ctrl[11][0] , \sa_ctrl[11].r.part0[0] );
tran (\sa_ctrl[11][0] , \sa_ctrl[11].f.sa_event_sel[0] );
tran (\sa_ctrl[10][31] , \sa_ctrl[10].r.part0[31] );
tran (\sa_ctrl[10][31] , \sa_ctrl[10].f.spare[26] );
tran (\sa_ctrl[10][30] , \sa_ctrl[10].r.part0[30] );
tran (\sa_ctrl[10][30] , \sa_ctrl[10].f.spare[25] );
tran (\sa_ctrl[10][29] , \sa_ctrl[10].r.part0[29] );
tran (\sa_ctrl[10][29] , \sa_ctrl[10].f.spare[24] );
tran (\sa_ctrl[10][28] , \sa_ctrl[10].r.part0[28] );
tran (\sa_ctrl[10][28] , \sa_ctrl[10].f.spare[23] );
tran (\sa_ctrl[10][27] , \sa_ctrl[10].r.part0[27] );
tran (\sa_ctrl[10][27] , \sa_ctrl[10].f.spare[22] );
tran (\sa_ctrl[10][26] , \sa_ctrl[10].r.part0[26] );
tran (\sa_ctrl[10][26] , \sa_ctrl[10].f.spare[21] );
tran (\sa_ctrl[10][25] , \sa_ctrl[10].r.part0[25] );
tran (\sa_ctrl[10][25] , \sa_ctrl[10].f.spare[20] );
tran (\sa_ctrl[10][24] , \sa_ctrl[10].r.part0[24] );
tran (\sa_ctrl[10][24] , \sa_ctrl[10].f.spare[19] );
tran (\sa_ctrl[10][23] , \sa_ctrl[10].r.part0[23] );
tran (\sa_ctrl[10][23] , \sa_ctrl[10].f.spare[18] );
tran (\sa_ctrl[10][22] , \sa_ctrl[10].r.part0[22] );
tran (\sa_ctrl[10][22] , \sa_ctrl[10].f.spare[17] );
tran (\sa_ctrl[10][21] , \sa_ctrl[10].r.part0[21] );
tran (\sa_ctrl[10][21] , \sa_ctrl[10].f.spare[16] );
tran (\sa_ctrl[10][20] , \sa_ctrl[10].r.part0[20] );
tran (\sa_ctrl[10][20] , \sa_ctrl[10].f.spare[15] );
tran (\sa_ctrl[10][19] , \sa_ctrl[10].r.part0[19] );
tran (\sa_ctrl[10][19] , \sa_ctrl[10].f.spare[14] );
tran (\sa_ctrl[10][18] , \sa_ctrl[10].r.part0[18] );
tran (\sa_ctrl[10][18] , \sa_ctrl[10].f.spare[13] );
tran (\sa_ctrl[10][17] , \sa_ctrl[10].r.part0[17] );
tran (\sa_ctrl[10][17] , \sa_ctrl[10].f.spare[12] );
tran (\sa_ctrl[10][16] , \sa_ctrl[10].r.part0[16] );
tran (\sa_ctrl[10][16] , \sa_ctrl[10].f.spare[11] );
tran (\sa_ctrl[10][15] , \sa_ctrl[10].r.part0[15] );
tran (\sa_ctrl[10][15] , \sa_ctrl[10].f.spare[10] );
tran (\sa_ctrl[10][14] , \sa_ctrl[10].r.part0[14] );
tran (\sa_ctrl[10][14] , \sa_ctrl[10].f.spare[9] );
tran (\sa_ctrl[10][13] , \sa_ctrl[10].r.part0[13] );
tran (\sa_ctrl[10][13] , \sa_ctrl[10].f.spare[8] );
tran (\sa_ctrl[10][12] , \sa_ctrl[10].r.part0[12] );
tran (\sa_ctrl[10][12] , \sa_ctrl[10].f.spare[7] );
tran (\sa_ctrl[10][11] , \sa_ctrl[10].r.part0[11] );
tran (\sa_ctrl[10][11] , \sa_ctrl[10].f.spare[6] );
tran (\sa_ctrl[10][10] , \sa_ctrl[10].r.part0[10] );
tran (\sa_ctrl[10][10] , \sa_ctrl[10].f.spare[5] );
tran (\sa_ctrl[10][9] , \sa_ctrl[10].r.part0[9] );
tran (\sa_ctrl[10][9] , \sa_ctrl[10].f.spare[4] );
tran (\sa_ctrl[10][8] , \sa_ctrl[10].r.part0[8] );
tran (\sa_ctrl[10][8] , \sa_ctrl[10].f.spare[3] );
tran (\sa_ctrl[10][7] , \sa_ctrl[10].r.part0[7] );
tran (\sa_ctrl[10][7] , \sa_ctrl[10].f.spare[2] );
tran (\sa_ctrl[10][6] , \sa_ctrl[10].r.part0[6] );
tran (\sa_ctrl[10][6] , \sa_ctrl[10].f.spare[1] );
tran (\sa_ctrl[10][5] , \sa_ctrl[10].r.part0[5] );
tran (\sa_ctrl[10][5] , \sa_ctrl[10].f.spare[0] );
tran (\sa_ctrl[10][4] , \sa_ctrl[10].r.part0[4] );
tran (\sa_ctrl[10][4] , \sa_ctrl[10].f.sa_event_sel[4] );
tran (\sa_ctrl[10][3] , \sa_ctrl[10].r.part0[3] );
tran (\sa_ctrl[10][3] , \sa_ctrl[10].f.sa_event_sel[3] );
tran (\sa_ctrl[10][2] , \sa_ctrl[10].r.part0[2] );
tran (\sa_ctrl[10][2] , \sa_ctrl[10].f.sa_event_sel[2] );
tran (\sa_ctrl[10][1] , \sa_ctrl[10].r.part0[1] );
tran (\sa_ctrl[10][1] , \sa_ctrl[10].f.sa_event_sel[1] );
tran (\sa_ctrl[10][0] , \sa_ctrl[10].r.part0[0] );
tran (\sa_ctrl[10][0] , \sa_ctrl[10].f.sa_event_sel[0] );
tran (\sa_ctrl[9][31] , \sa_ctrl[9].r.part0[31] );
tran (\sa_ctrl[9][31] , \sa_ctrl[9].f.spare[26] );
tran (\sa_ctrl[9][30] , \sa_ctrl[9].r.part0[30] );
tran (\sa_ctrl[9][30] , \sa_ctrl[9].f.spare[25] );
tran (\sa_ctrl[9][29] , \sa_ctrl[9].r.part0[29] );
tran (\sa_ctrl[9][29] , \sa_ctrl[9].f.spare[24] );
tran (\sa_ctrl[9][28] , \sa_ctrl[9].r.part0[28] );
tran (\sa_ctrl[9][28] , \sa_ctrl[9].f.spare[23] );
tran (\sa_ctrl[9][27] , \sa_ctrl[9].r.part0[27] );
tran (\sa_ctrl[9][27] , \sa_ctrl[9].f.spare[22] );
tran (\sa_ctrl[9][26] , \sa_ctrl[9].r.part0[26] );
tran (\sa_ctrl[9][26] , \sa_ctrl[9].f.spare[21] );
tran (\sa_ctrl[9][25] , \sa_ctrl[9].r.part0[25] );
tran (\sa_ctrl[9][25] , \sa_ctrl[9].f.spare[20] );
tran (\sa_ctrl[9][24] , \sa_ctrl[9].r.part0[24] );
tran (\sa_ctrl[9][24] , \sa_ctrl[9].f.spare[19] );
tran (\sa_ctrl[9][23] , \sa_ctrl[9].r.part0[23] );
tran (\sa_ctrl[9][23] , \sa_ctrl[9].f.spare[18] );
tran (\sa_ctrl[9][22] , \sa_ctrl[9].r.part0[22] );
tran (\sa_ctrl[9][22] , \sa_ctrl[9].f.spare[17] );
tran (\sa_ctrl[9][21] , \sa_ctrl[9].r.part0[21] );
tran (\sa_ctrl[9][21] , \sa_ctrl[9].f.spare[16] );
tran (\sa_ctrl[9][20] , \sa_ctrl[9].r.part0[20] );
tran (\sa_ctrl[9][20] , \sa_ctrl[9].f.spare[15] );
tran (\sa_ctrl[9][19] , \sa_ctrl[9].r.part0[19] );
tran (\sa_ctrl[9][19] , \sa_ctrl[9].f.spare[14] );
tran (\sa_ctrl[9][18] , \sa_ctrl[9].r.part0[18] );
tran (\sa_ctrl[9][18] , \sa_ctrl[9].f.spare[13] );
tran (\sa_ctrl[9][17] , \sa_ctrl[9].r.part0[17] );
tran (\sa_ctrl[9][17] , \sa_ctrl[9].f.spare[12] );
tran (\sa_ctrl[9][16] , \sa_ctrl[9].r.part0[16] );
tran (\sa_ctrl[9][16] , \sa_ctrl[9].f.spare[11] );
tran (\sa_ctrl[9][15] , \sa_ctrl[9].r.part0[15] );
tran (\sa_ctrl[9][15] , \sa_ctrl[9].f.spare[10] );
tran (\sa_ctrl[9][14] , \sa_ctrl[9].r.part0[14] );
tran (\sa_ctrl[9][14] , \sa_ctrl[9].f.spare[9] );
tran (\sa_ctrl[9][13] , \sa_ctrl[9].r.part0[13] );
tran (\sa_ctrl[9][13] , \sa_ctrl[9].f.spare[8] );
tran (\sa_ctrl[9][12] , \sa_ctrl[9].r.part0[12] );
tran (\sa_ctrl[9][12] , \sa_ctrl[9].f.spare[7] );
tran (\sa_ctrl[9][11] , \sa_ctrl[9].r.part0[11] );
tran (\sa_ctrl[9][11] , \sa_ctrl[9].f.spare[6] );
tran (\sa_ctrl[9][10] , \sa_ctrl[9].r.part0[10] );
tran (\sa_ctrl[9][10] , \sa_ctrl[9].f.spare[5] );
tran (\sa_ctrl[9][9] , \sa_ctrl[9].r.part0[9] );
tran (\sa_ctrl[9][9] , \sa_ctrl[9].f.spare[4] );
tran (\sa_ctrl[9][8] , \sa_ctrl[9].r.part0[8] );
tran (\sa_ctrl[9][8] , \sa_ctrl[9].f.spare[3] );
tran (\sa_ctrl[9][7] , \sa_ctrl[9].r.part0[7] );
tran (\sa_ctrl[9][7] , \sa_ctrl[9].f.spare[2] );
tran (\sa_ctrl[9][6] , \sa_ctrl[9].r.part0[6] );
tran (\sa_ctrl[9][6] , \sa_ctrl[9].f.spare[1] );
tran (\sa_ctrl[9][5] , \sa_ctrl[9].r.part0[5] );
tran (\sa_ctrl[9][5] , \sa_ctrl[9].f.spare[0] );
tran (\sa_ctrl[9][4] , \sa_ctrl[9].r.part0[4] );
tran (\sa_ctrl[9][4] , \sa_ctrl[9].f.sa_event_sel[4] );
tran (\sa_ctrl[9][3] , \sa_ctrl[9].r.part0[3] );
tran (\sa_ctrl[9][3] , \sa_ctrl[9].f.sa_event_sel[3] );
tran (\sa_ctrl[9][2] , \sa_ctrl[9].r.part0[2] );
tran (\sa_ctrl[9][2] , \sa_ctrl[9].f.sa_event_sel[2] );
tran (\sa_ctrl[9][1] , \sa_ctrl[9].r.part0[1] );
tran (\sa_ctrl[9][1] , \sa_ctrl[9].f.sa_event_sel[1] );
tran (\sa_ctrl[9][0] , \sa_ctrl[9].r.part0[0] );
tran (\sa_ctrl[9][0] , \sa_ctrl[9].f.sa_event_sel[0] );
tran (\sa_ctrl[8][31] , \sa_ctrl[8].r.part0[31] );
tran (\sa_ctrl[8][31] , \sa_ctrl[8].f.spare[26] );
tran (\sa_ctrl[8][30] , \sa_ctrl[8].r.part0[30] );
tran (\sa_ctrl[8][30] , \sa_ctrl[8].f.spare[25] );
tran (\sa_ctrl[8][29] , \sa_ctrl[8].r.part0[29] );
tran (\sa_ctrl[8][29] , \sa_ctrl[8].f.spare[24] );
tran (\sa_ctrl[8][28] , \sa_ctrl[8].r.part0[28] );
tran (\sa_ctrl[8][28] , \sa_ctrl[8].f.spare[23] );
tran (\sa_ctrl[8][27] , \sa_ctrl[8].r.part0[27] );
tran (\sa_ctrl[8][27] , \sa_ctrl[8].f.spare[22] );
tran (\sa_ctrl[8][26] , \sa_ctrl[8].r.part0[26] );
tran (\sa_ctrl[8][26] , \sa_ctrl[8].f.spare[21] );
tran (\sa_ctrl[8][25] , \sa_ctrl[8].r.part0[25] );
tran (\sa_ctrl[8][25] , \sa_ctrl[8].f.spare[20] );
tran (\sa_ctrl[8][24] , \sa_ctrl[8].r.part0[24] );
tran (\sa_ctrl[8][24] , \sa_ctrl[8].f.spare[19] );
tran (\sa_ctrl[8][23] , \sa_ctrl[8].r.part0[23] );
tran (\sa_ctrl[8][23] , \sa_ctrl[8].f.spare[18] );
tran (\sa_ctrl[8][22] , \sa_ctrl[8].r.part0[22] );
tran (\sa_ctrl[8][22] , \sa_ctrl[8].f.spare[17] );
tran (\sa_ctrl[8][21] , \sa_ctrl[8].r.part0[21] );
tran (\sa_ctrl[8][21] , \sa_ctrl[8].f.spare[16] );
tran (\sa_ctrl[8][20] , \sa_ctrl[8].r.part0[20] );
tran (\sa_ctrl[8][20] , \sa_ctrl[8].f.spare[15] );
tran (\sa_ctrl[8][19] , \sa_ctrl[8].r.part0[19] );
tran (\sa_ctrl[8][19] , \sa_ctrl[8].f.spare[14] );
tran (\sa_ctrl[8][18] , \sa_ctrl[8].r.part0[18] );
tran (\sa_ctrl[8][18] , \sa_ctrl[8].f.spare[13] );
tran (\sa_ctrl[8][17] , \sa_ctrl[8].r.part0[17] );
tran (\sa_ctrl[8][17] , \sa_ctrl[8].f.spare[12] );
tran (\sa_ctrl[8][16] , \sa_ctrl[8].r.part0[16] );
tran (\sa_ctrl[8][16] , \sa_ctrl[8].f.spare[11] );
tran (\sa_ctrl[8][15] , \sa_ctrl[8].r.part0[15] );
tran (\sa_ctrl[8][15] , \sa_ctrl[8].f.spare[10] );
tran (\sa_ctrl[8][14] , \sa_ctrl[8].r.part0[14] );
tran (\sa_ctrl[8][14] , \sa_ctrl[8].f.spare[9] );
tran (\sa_ctrl[8][13] , \sa_ctrl[8].r.part0[13] );
tran (\sa_ctrl[8][13] , \sa_ctrl[8].f.spare[8] );
tran (\sa_ctrl[8][12] , \sa_ctrl[8].r.part0[12] );
tran (\sa_ctrl[8][12] , \sa_ctrl[8].f.spare[7] );
tran (\sa_ctrl[8][11] , \sa_ctrl[8].r.part0[11] );
tran (\sa_ctrl[8][11] , \sa_ctrl[8].f.spare[6] );
tran (\sa_ctrl[8][10] , \sa_ctrl[8].r.part0[10] );
tran (\sa_ctrl[8][10] , \sa_ctrl[8].f.spare[5] );
tran (\sa_ctrl[8][9] , \sa_ctrl[8].r.part0[9] );
tran (\sa_ctrl[8][9] , \sa_ctrl[8].f.spare[4] );
tran (\sa_ctrl[8][8] , \sa_ctrl[8].r.part0[8] );
tran (\sa_ctrl[8][8] , \sa_ctrl[8].f.spare[3] );
tran (\sa_ctrl[8][7] , \sa_ctrl[8].r.part0[7] );
tran (\sa_ctrl[8][7] , \sa_ctrl[8].f.spare[2] );
tran (\sa_ctrl[8][6] , \sa_ctrl[8].r.part0[6] );
tran (\sa_ctrl[8][6] , \sa_ctrl[8].f.spare[1] );
tran (\sa_ctrl[8][5] , \sa_ctrl[8].r.part0[5] );
tran (\sa_ctrl[8][5] , \sa_ctrl[8].f.spare[0] );
tran (\sa_ctrl[8][4] , \sa_ctrl[8].r.part0[4] );
tran (\sa_ctrl[8][4] , \sa_ctrl[8].f.sa_event_sel[4] );
tran (\sa_ctrl[8][3] , \sa_ctrl[8].r.part0[3] );
tran (\sa_ctrl[8][3] , \sa_ctrl[8].f.sa_event_sel[3] );
tran (\sa_ctrl[8][2] , \sa_ctrl[8].r.part0[2] );
tran (\sa_ctrl[8][2] , \sa_ctrl[8].f.sa_event_sel[2] );
tran (\sa_ctrl[8][1] , \sa_ctrl[8].r.part0[1] );
tran (\sa_ctrl[8][1] , \sa_ctrl[8].f.sa_event_sel[1] );
tran (\sa_ctrl[8][0] , \sa_ctrl[8].r.part0[0] );
tran (\sa_ctrl[8][0] , \sa_ctrl[8].f.sa_event_sel[0] );
tran (\sa_ctrl[7][31] , \sa_ctrl[7].r.part0[31] );
tran (\sa_ctrl[7][31] , \sa_ctrl[7].f.spare[26] );
tran (\sa_ctrl[7][30] , \sa_ctrl[7].r.part0[30] );
tran (\sa_ctrl[7][30] , \sa_ctrl[7].f.spare[25] );
tran (\sa_ctrl[7][29] , \sa_ctrl[7].r.part0[29] );
tran (\sa_ctrl[7][29] , \sa_ctrl[7].f.spare[24] );
tran (\sa_ctrl[7][28] , \sa_ctrl[7].r.part0[28] );
tran (\sa_ctrl[7][28] , \sa_ctrl[7].f.spare[23] );
tran (\sa_ctrl[7][27] , \sa_ctrl[7].r.part0[27] );
tran (\sa_ctrl[7][27] , \sa_ctrl[7].f.spare[22] );
tran (\sa_ctrl[7][26] , \sa_ctrl[7].r.part0[26] );
tran (\sa_ctrl[7][26] , \sa_ctrl[7].f.spare[21] );
tran (\sa_ctrl[7][25] , \sa_ctrl[7].r.part0[25] );
tran (\sa_ctrl[7][25] , \sa_ctrl[7].f.spare[20] );
tran (\sa_ctrl[7][24] , \sa_ctrl[7].r.part0[24] );
tran (\sa_ctrl[7][24] , \sa_ctrl[7].f.spare[19] );
tran (\sa_ctrl[7][23] , \sa_ctrl[7].r.part0[23] );
tran (\sa_ctrl[7][23] , \sa_ctrl[7].f.spare[18] );
tran (\sa_ctrl[7][22] , \sa_ctrl[7].r.part0[22] );
tran (\sa_ctrl[7][22] , \sa_ctrl[7].f.spare[17] );
tran (\sa_ctrl[7][21] , \sa_ctrl[7].r.part0[21] );
tran (\sa_ctrl[7][21] , \sa_ctrl[7].f.spare[16] );
tran (\sa_ctrl[7][20] , \sa_ctrl[7].r.part0[20] );
tran (\sa_ctrl[7][20] , \sa_ctrl[7].f.spare[15] );
tran (\sa_ctrl[7][19] , \sa_ctrl[7].r.part0[19] );
tran (\sa_ctrl[7][19] , \sa_ctrl[7].f.spare[14] );
tran (\sa_ctrl[7][18] , \sa_ctrl[7].r.part0[18] );
tran (\sa_ctrl[7][18] , \sa_ctrl[7].f.spare[13] );
tran (\sa_ctrl[7][17] , \sa_ctrl[7].r.part0[17] );
tran (\sa_ctrl[7][17] , \sa_ctrl[7].f.spare[12] );
tran (\sa_ctrl[7][16] , \sa_ctrl[7].r.part0[16] );
tran (\sa_ctrl[7][16] , \sa_ctrl[7].f.spare[11] );
tran (\sa_ctrl[7][15] , \sa_ctrl[7].r.part0[15] );
tran (\sa_ctrl[7][15] , \sa_ctrl[7].f.spare[10] );
tran (\sa_ctrl[7][14] , \sa_ctrl[7].r.part0[14] );
tran (\sa_ctrl[7][14] , \sa_ctrl[7].f.spare[9] );
tran (\sa_ctrl[7][13] , \sa_ctrl[7].r.part0[13] );
tran (\sa_ctrl[7][13] , \sa_ctrl[7].f.spare[8] );
tran (\sa_ctrl[7][12] , \sa_ctrl[7].r.part0[12] );
tran (\sa_ctrl[7][12] , \sa_ctrl[7].f.spare[7] );
tran (\sa_ctrl[7][11] , \sa_ctrl[7].r.part0[11] );
tran (\sa_ctrl[7][11] , \sa_ctrl[7].f.spare[6] );
tran (\sa_ctrl[7][10] , \sa_ctrl[7].r.part0[10] );
tran (\sa_ctrl[7][10] , \sa_ctrl[7].f.spare[5] );
tran (\sa_ctrl[7][9] , \sa_ctrl[7].r.part0[9] );
tran (\sa_ctrl[7][9] , \sa_ctrl[7].f.spare[4] );
tran (\sa_ctrl[7][8] , \sa_ctrl[7].r.part0[8] );
tran (\sa_ctrl[7][8] , \sa_ctrl[7].f.spare[3] );
tran (\sa_ctrl[7][7] , \sa_ctrl[7].r.part0[7] );
tran (\sa_ctrl[7][7] , \sa_ctrl[7].f.spare[2] );
tran (\sa_ctrl[7][6] , \sa_ctrl[7].r.part0[6] );
tran (\sa_ctrl[7][6] , \sa_ctrl[7].f.spare[1] );
tran (\sa_ctrl[7][5] , \sa_ctrl[7].r.part0[5] );
tran (\sa_ctrl[7][5] , \sa_ctrl[7].f.spare[0] );
tran (\sa_ctrl[7][4] , \sa_ctrl[7].r.part0[4] );
tran (\sa_ctrl[7][4] , \sa_ctrl[7].f.sa_event_sel[4] );
tran (\sa_ctrl[7][3] , \sa_ctrl[7].r.part0[3] );
tran (\sa_ctrl[7][3] , \sa_ctrl[7].f.sa_event_sel[3] );
tran (\sa_ctrl[7][2] , \sa_ctrl[7].r.part0[2] );
tran (\sa_ctrl[7][2] , \sa_ctrl[7].f.sa_event_sel[2] );
tran (\sa_ctrl[7][1] , \sa_ctrl[7].r.part0[1] );
tran (\sa_ctrl[7][1] , \sa_ctrl[7].f.sa_event_sel[1] );
tran (\sa_ctrl[7][0] , \sa_ctrl[7].r.part0[0] );
tran (\sa_ctrl[7][0] , \sa_ctrl[7].f.sa_event_sel[0] );
tran (\sa_ctrl[6][31] , \sa_ctrl[6].r.part0[31] );
tran (\sa_ctrl[6][31] , \sa_ctrl[6].f.spare[26] );
tran (\sa_ctrl[6][30] , \sa_ctrl[6].r.part0[30] );
tran (\sa_ctrl[6][30] , \sa_ctrl[6].f.spare[25] );
tran (\sa_ctrl[6][29] , \sa_ctrl[6].r.part0[29] );
tran (\sa_ctrl[6][29] , \sa_ctrl[6].f.spare[24] );
tran (\sa_ctrl[6][28] , \sa_ctrl[6].r.part0[28] );
tran (\sa_ctrl[6][28] , \sa_ctrl[6].f.spare[23] );
tran (\sa_ctrl[6][27] , \sa_ctrl[6].r.part0[27] );
tran (\sa_ctrl[6][27] , \sa_ctrl[6].f.spare[22] );
tran (\sa_ctrl[6][26] , \sa_ctrl[6].r.part0[26] );
tran (\sa_ctrl[6][26] , \sa_ctrl[6].f.spare[21] );
tran (\sa_ctrl[6][25] , \sa_ctrl[6].r.part0[25] );
tran (\sa_ctrl[6][25] , \sa_ctrl[6].f.spare[20] );
tran (\sa_ctrl[6][24] , \sa_ctrl[6].r.part0[24] );
tran (\sa_ctrl[6][24] , \sa_ctrl[6].f.spare[19] );
tran (\sa_ctrl[6][23] , \sa_ctrl[6].r.part0[23] );
tran (\sa_ctrl[6][23] , \sa_ctrl[6].f.spare[18] );
tran (\sa_ctrl[6][22] , \sa_ctrl[6].r.part0[22] );
tran (\sa_ctrl[6][22] , \sa_ctrl[6].f.spare[17] );
tran (\sa_ctrl[6][21] , \sa_ctrl[6].r.part0[21] );
tran (\sa_ctrl[6][21] , \sa_ctrl[6].f.spare[16] );
tran (\sa_ctrl[6][20] , \sa_ctrl[6].r.part0[20] );
tran (\sa_ctrl[6][20] , \sa_ctrl[6].f.spare[15] );
tran (\sa_ctrl[6][19] , \sa_ctrl[6].r.part0[19] );
tran (\sa_ctrl[6][19] , \sa_ctrl[6].f.spare[14] );
tran (\sa_ctrl[6][18] , \sa_ctrl[6].r.part0[18] );
tran (\sa_ctrl[6][18] , \sa_ctrl[6].f.spare[13] );
tran (\sa_ctrl[6][17] , \sa_ctrl[6].r.part0[17] );
tran (\sa_ctrl[6][17] , \sa_ctrl[6].f.spare[12] );
tran (\sa_ctrl[6][16] , \sa_ctrl[6].r.part0[16] );
tran (\sa_ctrl[6][16] , \sa_ctrl[6].f.spare[11] );
tran (\sa_ctrl[6][15] , \sa_ctrl[6].r.part0[15] );
tran (\sa_ctrl[6][15] , \sa_ctrl[6].f.spare[10] );
tran (\sa_ctrl[6][14] , \sa_ctrl[6].r.part0[14] );
tran (\sa_ctrl[6][14] , \sa_ctrl[6].f.spare[9] );
tran (\sa_ctrl[6][13] , \sa_ctrl[6].r.part0[13] );
tran (\sa_ctrl[6][13] , \sa_ctrl[6].f.spare[8] );
tran (\sa_ctrl[6][12] , \sa_ctrl[6].r.part0[12] );
tran (\sa_ctrl[6][12] , \sa_ctrl[6].f.spare[7] );
tran (\sa_ctrl[6][11] , \sa_ctrl[6].r.part0[11] );
tran (\sa_ctrl[6][11] , \sa_ctrl[6].f.spare[6] );
tran (\sa_ctrl[6][10] , \sa_ctrl[6].r.part0[10] );
tran (\sa_ctrl[6][10] , \sa_ctrl[6].f.spare[5] );
tran (\sa_ctrl[6][9] , \sa_ctrl[6].r.part0[9] );
tran (\sa_ctrl[6][9] , \sa_ctrl[6].f.spare[4] );
tran (\sa_ctrl[6][8] , \sa_ctrl[6].r.part0[8] );
tran (\sa_ctrl[6][8] , \sa_ctrl[6].f.spare[3] );
tran (\sa_ctrl[6][7] , \sa_ctrl[6].r.part0[7] );
tran (\sa_ctrl[6][7] , \sa_ctrl[6].f.spare[2] );
tran (\sa_ctrl[6][6] , \sa_ctrl[6].r.part0[6] );
tran (\sa_ctrl[6][6] , \sa_ctrl[6].f.spare[1] );
tran (\sa_ctrl[6][5] , \sa_ctrl[6].r.part0[5] );
tran (\sa_ctrl[6][5] , \sa_ctrl[6].f.spare[0] );
tran (\sa_ctrl[6][4] , \sa_ctrl[6].r.part0[4] );
tran (\sa_ctrl[6][4] , \sa_ctrl[6].f.sa_event_sel[4] );
tran (\sa_ctrl[6][3] , \sa_ctrl[6].r.part0[3] );
tran (\sa_ctrl[6][3] , \sa_ctrl[6].f.sa_event_sel[3] );
tran (\sa_ctrl[6][2] , \sa_ctrl[6].r.part0[2] );
tran (\sa_ctrl[6][2] , \sa_ctrl[6].f.sa_event_sel[2] );
tran (\sa_ctrl[6][1] , \sa_ctrl[6].r.part0[1] );
tran (\sa_ctrl[6][1] , \sa_ctrl[6].f.sa_event_sel[1] );
tran (\sa_ctrl[6][0] , \sa_ctrl[6].r.part0[0] );
tran (\sa_ctrl[6][0] , \sa_ctrl[6].f.sa_event_sel[0] );
tran (\sa_ctrl[5][31] , \sa_ctrl[5].r.part0[31] );
tran (\sa_ctrl[5][31] , \sa_ctrl[5].f.spare[26] );
tran (\sa_ctrl[5][30] , \sa_ctrl[5].r.part0[30] );
tran (\sa_ctrl[5][30] , \sa_ctrl[5].f.spare[25] );
tran (\sa_ctrl[5][29] , \sa_ctrl[5].r.part0[29] );
tran (\sa_ctrl[5][29] , \sa_ctrl[5].f.spare[24] );
tran (\sa_ctrl[5][28] , \sa_ctrl[5].r.part0[28] );
tran (\sa_ctrl[5][28] , \sa_ctrl[5].f.spare[23] );
tran (\sa_ctrl[5][27] , \sa_ctrl[5].r.part0[27] );
tran (\sa_ctrl[5][27] , \sa_ctrl[5].f.spare[22] );
tran (\sa_ctrl[5][26] , \sa_ctrl[5].r.part0[26] );
tran (\sa_ctrl[5][26] , \sa_ctrl[5].f.spare[21] );
tran (\sa_ctrl[5][25] , \sa_ctrl[5].r.part0[25] );
tran (\sa_ctrl[5][25] , \sa_ctrl[5].f.spare[20] );
tran (\sa_ctrl[5][24] , \sa_ctrl[5].r.part0[24] );
tran (\sa_ctrl[5][24] , \sa_ctrl[5].f.spare[19] );
tran (\sa_ctrl[5][23] , \sa_ctrl[5].r.part0[23] );
tran (\sa_ctrl[5][23] , \sa_ctrl[5].f.spare[18] );
tran (\sa_ctrl[5][22] , \sa_ctrl[5].r.part0[22] );
tran (\sa_ctrl[5][22] , \sa_ctrl[5].f.spare[17] );
tran (\sa_ctrl[5][21] , \sa_ctrl[5].r.part0[21] );
tran (\sa_ctrl[5][21] , \sa_ctrl[5].f.spare[16] );
tran (\sa_ctrl[5][20] , \sa_ctrl[5].r.part0[20] );
tran (\sa_ctrl[5][20] , \sa_ctrl[5].f.spare[15] );
tran (\sa_ctrl[5][19] , \sa_ctrl[5].r.part0[19] );
tran (\sa_ctrl[5][19] , \sa_ctrl[5].f.spare[14] );
tran (\sa_ctrl[5][18] , \sa_ctrl[5].r.part0[18] );
tran (\sa_ctrl[5][18] , \sa_ctrl[5].f.spare[13] );
tran (\sa_ctrl[5][17] , \sa_ctrl[5].r.part0[17] );
tran (\sa_ctrl[5][17] , \sa_ctrl[5].f.spare[12] );
tran (\sa_ctrl[5][16] , \sa_ctrl[5].r.part0[16] );
tran (\sa_ctrl[5][16] , \sa_ctrl[5].f.spare[11] );
tran (\sa_ctrl[5][15] , \sa_ctrl[5].r.part0[15] );
tran (\sa_ctrl[5][15] , \sa_ctrl[5].f.spare[10] );
tran (\sa_ctrl[5][14] , \sa_ctrl[5].r.part0[14] );
tran (\sa_ctrl[5][14] , \sa_ctrl[5].f.spare[9] );
tran (\sa_ctrl[5][13] , \sa_ctrl[5].r.part0[13] );
tran (\sa_ctrl[5][13] , \sa_ctrl[5].f.spare[8] );
tran (\sa_ctrl[5][12] , \sa_ctrl[5].r.part0[12] );
tran (\sa_ctrl[5][12] , \sa_ctrl[5].f.spare[7] );
tran (\sa_ctrl[5][11] , \sa_ctrl[5].r.part0[11] );
tran (\sa_ctrl[5][11] , \sa_ctrl[5].f.spare[6] );
tran (\sa_ctrl[5][10] , \sa_ctrl[5].r.part0[10] );
tran (\sa_ctrl[5][10] , \sa_ctrl[5].f.spare[5] );
tran (\sa_ctrl[5][9] , \sa_ctrl[5].r.part0[9] );
tran (\sa_ctrl[5][9] , \sa_ctrl[5].f.spare[4] );
tran (\sa_ctrl[5][8] , \sa_ctrl[5].r.part0[8] );
tran (\sa_ctrl[5][8] , \sa_ctrl[5].f.spare[3] );
tran (\sa_ctrl[5][7] , \sa_ctrl[5].r.part0[7] );
tran (\sa_ctrl[5][7] , \sa_ctrl[5].f.spare[2] );
tran (\sa_ctrl[5][6] , \sa_ctrl[5].r.part0[6] );
tran (\sa_ctrl[5][6] , \sa_ctrl[5].f.spare[1] );
tran (\sa_ctrl[5][5] , \sa_ctrl[5].r.part0[5] );
tran (\sa_ctrl[5][5] , \sa_ctrl[5].f.spare[0] );
tran (\sa_ctrl[5][4] , \sa_ctrl[5].r.part0[4] );
tran (\sa_ctrl[5][4] , \sa_ctrl[5].f.sa_event_sel[4] );
tran (\sa_ctrl[5][3] , \sa_ctrl[5].r.part0[3] );
tran (\sa_ctrl[5][3] , \sa_ctrl[5].f.sa_event_sel[3] );
tran (\sa_ctrl[5][2] , \sa_ctrl[5].r.part0[2] );
tran (\sa_ctrl[5][2] , \sa_ctrl[5].f.sa_event_sel[2] );
tran (\sa_ctrl[5][1] , \sa_ctrl[5].r.part0[1] );
tran (\sa_ctrl[5][1] , \sa_ctrl[5].f.sa_event_sel[1] );
tran (\sa_ctrl[5][0] , \sa_ctrl[5].r.part0[0] );
tran (\sa_ctrl[5][0] , \sa_ctrl[5].f.sa_event_sel[0] );
tran (\sa_ctrl[4][31] , \sa_ctrl[4].r.part0[31] );
tran (\sa_ctrl[4][31] , \sa_ctrl[4].f.spare[26] );
tran (\sa_ctrl[4][30] , \sa_ctrl[4].r.part0[30] );
tran (\sa_ctrl[4][30] , \sa_ctrl[4].f.spare[25] );
tran (\sa_ctrl[4][29] , \sa_ctrl[4].r.part0[29] );
tran (\sa_ctrl[4][29] , \sa_ctrl[4].f.spare[24] );
tran (\sa_ctrl[4][28] , \sa_ctrl[4].r.part0[28] );
tran (\sa_ctrl[4][28] , \sa_ctrl[4].f.spare[23] );
tran (\sa_ctrl[4][27] , \sa_ctrl[4].r.part0[27] );
tran (\sa_ctrl[4][27] , \sa_ctrl[4].f.spare[22] );
tran (\sa_ctrl[4][26] , \sa_ctrl[4].r.part0[26] );
tran (\sa_ctrl[4][26] , \sa_ctrl[4].f.spare[21] );
tran (\sa_ctrl[4][25] , \sa_ctrl[4].r.part0[25] );
tran (\sa_ctrl[4][25] , \sa_ctrl[4].f.spare[20] );
tran (\sa_ctrl[4][24] , \sa_ctrl[4].r.part0[24] );
tran (\sa_ctrl[4][24] , \sa_ctrl[4].f.spare[19] );
tran (\sa_ctrl[4][23] , \sa_ctrl[4].r.part0[23] );
tran (\sa_ctrl[4][23] , \sa_ctrl[4].f.spare[18] );
tran (\sa_ctrl[4][22] , \sa_ctrl[4].r.part0[22] );
tran (\sa_ctrl[4][22] , \sa_ctrl[4].f.spare[17] );
tran (\sa_ctrl[4][21] , \sa_ctrl[4].r.part0[21] );
tran (\sa_ctrl[4][21] , \sa_ctrl[4].f.spare[16] );
tran (\sa_ctrl[4][20] , \sa_ctrl[4].r.part0[20] );
tran (\sa_ctrl[4][20] , \sa_ctrl[4].f.spare[15] );
tran (\sa_ctrl[4][19] , \sa_ctrl[4].r.part0[19] );
tran (\sa_ctrl[4][19] , \sa_ctrl[4].f.spare[14] );
tran (\sa_ctrl[4][18] , \sa_ctrl[4].r.part0[18] );
tran (\sa_ctrl[4][18] , \sa_ctrl[4].f.spare[13] );
tran (\sa_ctrl[4][17] , \sa_ctrl[4].r.part0[17] );
tran (\sa_ctrl[4][17] , \sa_ctrl[4].f.spare[12] );
tran (\sa_ctrl[4][16] , \sa_ctrl[4].r.part0[16] );
tran (\sa_ctrl[4][16] , \sa_ctrl[4].f.spare[11] );
tran (\sa_ctrl[4][15] , \sa_ctrl[4].r.part0[15] );
tran (\sa_ctrl[4][15] , \sa_ctrl[4].f.spare[10] );
tran (\sa_ctrl[4][14] , \sa_ctrl[4].r.part0[14] );
tran (\sa_ctrl[4][14] , \sa_ctrl[4].f.spare[9] );
tran (\sa_ctrl[4][13] , \sa_ctrl[4].r.part0[13] );
tran (\sa_ctrl[4][13] , \sa_ctrl[4].f.spare[8] );
tran (\sa_ctrl[4][12] , \sa_ctrl[4].r.part0[12] );
tran (\sa_ctrl[4][12] , \sa_ctrl[4].f.spare[7] );
tran (\sa_ctrl[4][11] , \sa_ctrl[4].r.part0[11] );
tran (\sa_ctrl[4][11] , \sa_ctrl[4].f.spare[6] );
tran (\sa_ctrl[4][10] , \sa_ctrl[4].r.part0[10] );
tran (\sa_ctrl[4][10] , \sa_ctrl[4].f.spare[5] );
tran (\sa_ctrl[4][9] , \sa_ctrl[4].r.part0[9] );
tran (\sa_ctrl[4][9] , \sa_ctrl[4].f.spare[4] );
tran (\sa_ctrl[4][8] , \sa_ctrl[4].r.part0[8] );
tran (\sa_ctrl[4][8] , \sa_ctrl[4].f.spare[3] );
tran (\sa_ctrl[4][7] , \sa_ctrl[4].r.part0[7] );
tran (\sa_ctrl[4][7] , \sa_ctrl[4].f.spare[2] );
tran (\sa_ctrl[4][6] , \sa_ctrl[4].r.part0[6] );
tran (\sa_ctrl[4][6] , \sa_ctrl[4].f.spare[1] );
tran (\sa_ctrl[4][5] , \sa_ctrl[4].r.part0[5] );
tran (\sa_ctrl[4][5] , \sa_ctrl[4].f.spare[0] );
tran (\sa_ctrl[4][4] , \sa_ctrl[4].r.part0[4] );
tran (\sa_ctrl[4][4] , \sa_ctrl[4].f.sa_event_sel[4] );
tran (\sa_ctrl[4][3] , \sa_ctrl[4].r.part0[3] );
tran (\sa_ctrl[4][3] , \sa_ctrl[4].f.sa_event_sel[3] );
tran (\sa_ctrl[4][2] , \sa_ctrl[4].r.part0[2] );
tran (\sa_ctrl[4][2] , \sa_ctrl[4].f.sa_event_sel[2] );
tran (\sa_ctrl[4][1] , \sa_ctrl[4].r.part0[1] );
tran (\sa_ctrl[4][1] , \sa_ctrl[4].f.sa_event_sel[1] );
tran (\sa_ctrl[4][0] , \sa_ctrl[4].r.part0[0] );
tran (\sa_ctrl[4][0] , \sa_ctrl[4].f.sa_event_sel[0] );
tran (\sa_ctrl[3][31] , \sa_ctrl[3].r.part0[31] );
tran (\sa_ctrl[3][31] , \sa_ctrl[3].f.spare[26] );
tran (\sa_ctrl[3][30] , \sa_ctrl[3].r.part0[30] );
tran (\sa_ctrl[3][30] , \sa_ctrl[3].f.spare[25] );
tran (\sa_ctrl[3][29] , \sa_ctrl[3].r.part0[29] );
tran (\sa_ctrl[3][29] , \sa_ctrl[3].f.spare[24] );
tran (\sa_ctrl[3][28] , \sa_ctrl[3].r.part0[28] );
tran (\sa_ctrl[3][28] , \sa_ctrl[3].f.spare[23] );
tran (\sa_ctrl[3][27] , \sa_ctrl[3].r.part0[27] );
tran (\sa_ctrl[3][27] , \sa_ctrl[3].f.spare[22] );
tran (\sa_ctrl[3][26] , \sa_ctrl[3].r.part0[26] );
tran (\sa_ctrl[3][26] , \sa_ctrl[3].f.spare[21] );
tran (\sa_ctrl[3][25] , \sa_ctrl[3].r.part0[25] );
tran (\sa_ctrl[3][25] , \sa_ctrl[3].f.spare[20] );
tran (\sa_ctrl[3][24] , \sa_ctrl[3].r.part0[24] );
tran (\sa_ctrl[3][24] , \sa_ctrl[3].f.spare[19] );
tran (\sa_ctrl[3][23] , \sa_ctrl[3].r.part0[23] );
tran (\sa_ctrl[3][23] , \sa_ctrl[3].f.spare[18] );
tran (\sa_ctrl[3][22] , \sa_ctrl[3].r.part0[22] );
tran (\sa_ctrl[3][22] , \sa_ctrl[3].f.spare[17] );
tran (\sa_ctrl[3][21] , \sa_ctrl[3].r.part0[21] );
tran (\sa_ctrl[3][21] , \sa_ctrl[3].f.spare[16] );
tran (\sa_ctrl[3][20] , \sa_ctrl[3].r.part0[20] );
tran (\sa_ctrl[3][20] , \sa_ctrl[3].f.spare[15] );
tran (\sa_ctrl[3][19] , \sa_ctrl[3].r.part0[19] );
tran (\sa_ctrl[3][19] , \sa_ctrl[3].f.spare[14] );
tran (\sa_ctrl[3][18] , \sa_ctrl[3].r.part0[18] );
tran (\sa_ctrl[3][18] , \sa_ctrl[3].f.spare[13] );
tran (\sa_ctrl[3][17] , \sa_ctrl[3].r.part0[17] );
tran (\sa_ctrl[3][17] , \sa_ctrl[3].f.spare[12] );
tran (\sa_ctrl[3][16] , \sa_ctrl[3].r.part0[16] );
tran (\sa_ctrl[3][16] , \sa_ctrl[3].f.spare[11] );
tran (\sa_ctrl[3][15] , \sa_ctrl[3].r.part0[15] );
tran (\sa_ctrl[3][15] , \sa_ctrl[3].f.spare[10] );
tran (\sa_ctrl[3][14] , \sa_ctrl[3].r.part0[14] );
tran (\sa_ctrl[3][14] , \sa_ctrl[3].f.spare[9] );
tran (\sa_ctrl[3][13] , \sa_ctrl[3].r.part0[13] );
tran (\sa_ctrl[3][13] , \sa_ctrl[3].f.spare[8] );
tran (\sa_ctrl[3][12] , \sa_ctrl[3].r.part0[12] );
tran (\sa_ctrl[3][12] , \sa_ctrl[3].f.spare[7] );
tran (\sa_ctrl[3][11] , \sa_ctrl[3].r.part0[11] );
tran (\sa_ctrl[3][11] , \sa_ctrl[3].f.spare[6] );
tran (\sa_ctrl[3][10] , \sa_ctrl[3].r.part0[10] );
tran (\sa_ctrl[3][10] , \sa_ctrl[3].f.spare[5] );
tran (\sa_ctrl[3][9] , \sa_ctrl[3].r.part0[9] );
tran (\sa_ctrl[3][9] , \sa_ctrl[3].f.spare[4] );
tran (\sa_ctrl[3][8] , \sa_ctrl[3].r.part0[8] );
tran (\sa_ctrl[3][8] , \sa_ctrl[3].f.spare[3] );
tran (\sa_ctrl[3][7] , \sa_ctrl[3].r.part0[7] );
tran (\sa_ctrl[3][7] , \sa_ctrl[3].f.spare[2] );
tran (\sa_ctrl[3][6] , \sa_ctrl[3].r.part0[6] );
tran (\sa_ctrl[3][6] , \sa_ctrl[3].f.spare[1] );
tran (\sa_ctrl[3][5] , \sa_ctrl[3].r.part0[5] );
tran (\sa_ctrl[3][5] , \sa_ctrl[3].f.spare[0] );
tran (\sa_ctrl[3][4] , \sa_ctrl[3].r.part0[4] );
tran (\sa_ctrl[3][4] , \sa_ctrl[3].f.sa_event_sel[4] );
tran (\sa_ctrl[3][3] , \sa_ctrl[3].r.part0[3] );
tran (\sa_ctrl[3][3] , \sa_ctrl[3].f.sa_event_sel[3] );
tran (\sa_ctrl[3][2] , \sa_ctrl[3].r.part0[2] );
tran (\sa_ctrl[3][2] , \sa_ctrl[3].f.sa_event_sel[2] );
tran (\sa_ctrl[3][1] , \sa_ctrl[3].r.part0[1] );
tran (\sa_ctrl[3][1] , \sa_ctrl[3].f.sa_event_sel[1] );
tran (\sa_ctrl[3][0] , \sa_ctrl[3].r.part0[0] );
tran (\sa_ctrl[3][0] , \sa_ctrl[3].f.sa_event_sel[0] );
tran (\sa_ctrl[2][31] , \sa_ctrl[2].r.part0[31] );
tran (\sa_ctrl[2][31] , \sa_ctrl[2].f.spare[26] );
tran (\sa_ctrl[2][30] , \sa_ctrl[2].r.part0[30] );
tran (\sa_ctrl[2][30] , \sa_ctrl[2].f.spare[25] );
tran (\sa_ctrl[2][29] , \sa_ctrl[2].r.part0[29] );
tran (\sa_ctrl[2][29] , \sa_ctrl[2].f.spare[24] );
tran (\sa_ctrl[2][28] , \sa_ctrl[2].r.part0[28] );
tran (\sa_ctrl[2][28] , \sa_ctrl[2].f.spare[23] );
tran (\sa_ctrl[2][27] , \sa_ctrl[2].r.part0[27] );
tran (\sa_ctrl[2][27] , \sa_ctrl[2].f.spare[22] );
tran (\sa_ctrl[2][26] , \sa_ctrl[2].r.part0[26] );
tran (\sa_ctrl[2][26] , \sa_ctrl[2].f.spare[21] );
tran (\sa_ctrl[2][25] , \sa_ctrl[2].r.part0[25] );
tran (\sa_ctrl[2][25] , \sa_ctrl[2].f.spare[20] );
tran (\sa_ctrl[2][24] , \sa_ctrl[2].r.part0[24] );
tran (\sa_ctrl[2][24] , \sa_ctrl[2].f.spare[19] );
tran (\sa_ctrl[2][23] , \sa_ctrl[2].r.part0[23] );
tran (\sa_ctrl[2][23] , \sa_ctrl[2].f.spare[18] );
tran (\sa_ctrl[2][22] , \sa_ctrl[2].r.part0[22] );
tran (\sa_ctrl[2][22] , \sa_ctrl[2].f.spare[17] );
tran (\sa_ctrl[2][21] , \sa_ctrl[2].r.part0[21] );
tran (\sa_ctrl[2][21] , \sa_ctrl[2].f.spare[16] );
tran (\sa_ctrl[2][20] , \sa_ctrl[2].r.part0[20] );
tran (\sa_ctrl[2][20] , \sa_ctrl[2].f.spare[15] );
tran (\sa_ctrl[2][19] , \sa_ctrl[2].r.part0[19] );
tran (\sa_ctrl[2][19] , \sa_ctrl[2].f.spare[14] );
tran (\sa_ctrl[2][18] , \sa_ctrl[2].r.part0[18] );
tran (\sa_ctrl[2][18] , \sa_ctrl[2].f.spare[13] );
tran (\sa_ctrl[2][17] , \sa_ctrl[2].r.part0[17] );
tran (\sa_ctrl[2][17] , \sa_ctrl[2].f.spare[12] );
tran (\sa_ctrl[2][16] , \sa_ctrl[2].r.part0[16] );
tran (\sa_ctrl[2][16] , \sa_ctrl[2].f.spare[11] );
tran (\sa_ctrl[2][15] , \sa_ctrl[2].r.part0[15] );
tran (\sa_ctrl[2][15] , \sa_ctrl[2].f.spare[10] );
tran (\sa_ctrl[2][14] , \sa_ctrl[2].r.part0[14] );
tran (\sa_ctrl[2][14] , \sa_ctrl[2].f.spare[9] );
tran (\sa_ctrl[2][13] , \sa_ctrl[2].r.part0[13] );
tran (\sa_ctrl[2][13] , \sa_ctrl[2].f.spare[8] );
tran (\sa_ctrl[2][12] , \sa_ctrl[2].r.part0[12] );
tran (\sa_ctrl[2][12] , \sa_ctrl[2].f.spare[7] );
tran (\sa_ctrl[2][11] , \sa_ctrl[2].r.part0[11] );
tran (\sa_ctrl[2][11] , \sa_ctrl[2].f.spare[6] );
tran (\sa_ctrl[2][10] , \sa_ctrl[2].r.part0[10] );
tran (\sa_ctrl[2][10] , \sa_ctrl[2].f.spare[5] );
tran (\sa_ctrl[2][9] , \sa_ctrl[2].r.part0[9] );
tran (\sa_ctrl[2][9] , \sa_ctrl[2].f.spare[4] );
tran (\sa_ctrl[2][8] , \sa_ctrl[2].r.part0[8] );
tran (\sa_ctrl[2][8] , \sa_ctrl[2].f.spare[3] );
tran (\sa_ctrl[2][7] , \sa_ctrl[2].r.part0[7] );
tran (\sa_ctrl[2][7] , \sa_ctrl[2].f.spare[2] );
tran (\sa_ctrl[2][6] , \sa_ctrl[2].r.part0[6] );
tran (\sa_ctrl[2][6] , \sa_ctrl[2].f.spare[1] );
tran (\sa_ctrl[2][5] , \sa_ctrl[2].r.part0[5] );
tran (\sa_ctrl[2][5] , \sa_ctrl[2].f.spare[0] );
tran (\sa_ctrl[2][4] , \sa_ctrl[2].r.part0[4] );
tran (\sa_ctrl[2][4] , \sa_ctrl[2].f.sa_event_sel[4] );
tran (\sa_ctrl[2][3] , \sa_ctrl[2].r.part0[3] );
tran (\sa_ctrl[2][3] , \sa_ctrl[2].f.sa_event_sel[3] );
tran (\sa_ctrl[2][2] , \sa_ctrl[2].r.part0[2] );
tran (\sa_ctrl[2][2] , \sa_ctrl[2].f.sa_event_sel[2] );
tran (\sa_ctrl[2][1] , \sa_ctrl[2].r.part0[1] );
tran (\sa_ctrl[2][1] , \sa_ctrl[2].f.sa_event_sel[1] );
tran (\sa_ctrl[2][0] , \sa_ctrl[2].r.part0[0] );
tran (\sa_ctrl[2][0] , \sa_ctrl[2].f.sa_event_sel[0] );
tran (\sa_ctrl[1][31] , \sa_ctrl[1].r.part0[31] );
tran (\sa_ctrl[1][31] , \sa_ctrl[1].f.spare[26] );
tran (\sa_ctrl[1][30] , \sa_ctrl[1].r.part0[30] );
tran (\sa_ctrl[1][30] , \sa_ctrl[1].f.spare[25] );
tran (\sa_ctrl[1][29] , \sa_ctrl[1].r.part0[29] );
tran (\sa_ctrl[1][29] , \sa_ctrl[1].f.spare[24] );
tran (\sa_ctrl[1][28] , \sa_ctrl[1].r.part0[28] );
tran (\sa_ctrl[1][28] , \sa_ctrl[1].f.spare[23] );
tran (\sa_ctrl[1][27] , \sa_ctrl[1].r.part0[27] );
tran (\sa_ctrl[1][27] , \sa_ctrl[1].f.spare[22] );
tran (\sa_ctrl[1][26] , \sa_ctrl[1].r.part0[26] );
tran (\sa_ctrl[1][26] , \sa_ctrl[1].f.spare[21] );
tran (\sa_ctrl[1][25] , \sa_ctrl[1].r.part0[25] );
tran (\sa_ctrl[1][25] , \sa_ctrl[1].f.spare[20] );
tran (\sa_ctrl[1][24] , \sa_ctrl[1].r.part0[24] );
tran (\sa_ctrl[1][24] , \sa_ctrl[1].f.spare[19] );
tran (\sa_ctrl[1][23] , \sa_ctrl[1].r.part0[23] );
tran (\sa_ctrl[1][23] , \sa_ctrl[1].f.spare[18] );
tran (\sa_ctrl[1][22] , \sa_ctrl[1].r.part0[22] );
tran (\sa_ctrl[1][22] , \sa_ctrl[1].f.spare[17] );
tran (\sa_ctrl[1][21] , \sa_ctrl[1].r.part0[21] );
tran (\sa_ctrl[1][21] , \sa_ctrl[1].f.spare[16] );
tran (\sa_ctrl[1][20] , \sa_ctrl[1].r.part0[20] );
tran (\sa_ctrl[1][20] , \sa_ctrl[1].f.spare[15] );
tran (\sa_ctrl[1][19] , \sa_ctrl[1].r.part0[19] );
tran (\sa_ctrl[1][19] , \sa_ctrl[1].f.spare[14] );
tran (\sa_ctrl[1][18] , \sa_ctrl[1].r.part0[18] );
tran (\sa_ctrl[1][18] , \sa_ctrl[1].f.spare[13] );
tran (\sa_ctrl[1][17] , \sa_ctrl[1].r.part0[17] );
tran (\sa_ctrl[1][17] , \sa_ctrl[1].f.spare[12] );
tran (\sa_ctrl[1][16] , \sa_ctrl[1].r.part0[16] );
tran (\sa_ctrl[1][16] , \sa_ctrl[1].f.spare[11] );
tran (\sa_ctrl[1][15] , \sa_ctrl[1].r.part0[15] );
tran (\sa_ctrl[1][15] , \sa_ctrl[1].f.spare[10] );
tran (\sa_ctrl[1][14] , \sa_ctrl[1].r.part0[14] );
tran (\sa_ctrl[1][14] , \sa_ctrl[1].f.spare[9] );
tran (\sa_ctrl[1][13] , \sa_ctrl[1].r.part0[13] );
tran (\sa_ctrl[1][13] , \sa_ctrl[1].f.spare[8] );
tran (\sa_ctrl[1][12] , \sa_ctrl[1].r.part0[12] );
tran (\sa_ctrl[1][12] , \sa_ctrl[1].f.spare[7] );
tran (\sa_ctrl[1][11] , \sa_ctrl[1].r.part0[11] );
tran (\sa_ctrl[1][11] , \sa_ctrl[1].f.spare[6] );
tran (\sa_ctrl[1][10] , \sa_ctrl[1].r.part0[10] );
tran (\sa_ctrl[1][10] , \sa_ctrl[1].f.spare[5] );
tran (\sa_ctrl[1][9] , \sa_ctrl[1].r.part0[9] );
tran (\sa_ctrl[1][9] , \sa_ctrl[1].f.spare[4] );
tran (\sa_ctrl[1][8] , \sa_ctrl[1].r.part0[8] );
tran (\sa_ctrl[1][8] , \sa_ctrl[1].f.spare[3] );
tran (\sa_ctrl[1][7] , \sa_ctrl[1].r.part0[7] );
tran (\sa_ctrl[1][7] , \sa_ctrl[1].f.spare[2] );
tran (\sa_ctrl[1][6] , \sa_ctrl[1].r.part0[6] );
tran (\sa_ctrl[1][6] , \sa_ctrl[1].f.spare[1] );
tran (\sa_ctrl[1][5] , \sa_ctrl[1].r.part0[5] );
tran (\sa_ctrl[1][5] , \sa_ctrl[1].f.spare[0] );
tran (\sa_ctrl[1][4] , \sa_ctrl[1].r.part0[4] );
tran (\sa_ctrl[1][4] , \sa_ctrl[1].f.sa_event_sel[4] );
tran (\sa_ctrl[1][3] , \sa_ctrl[1].r.part0[3] );
tran (\sa_ctrl[1][3] , \sa_ctrl[1].f.sa_event_sel[3] );
tran (\sa_ctrl[1][2] , \sa_ctrl[1].r.part0[2] );
tran (\sa_ctrl[1][2] , \sa_ctrl[1].f.sa_event_sel[2] );
tran (\sa_ctrl[1][1] , \sa_ctrl[1].r.part0[1] );
tran (\sa_ctrl[1][1] , \sa_ctrl[1].f.sa_event_sel[1] );
tran (\sa_ctrl[1][0] , \sa_ctrl[1].r.part0[0] );
tran (\sa_ctrl[1][0] , \sa_ctrl[1].f.sa_event_sel[0] );
tran (\sa_ctrl[0][31] , \sa_ctrl[0].r.part0[31] );
tran (\sa_ctrl[0][31] , \sa_ctrl[0].f.spare[26] );
tran (\sa_ctrl[0][30] , \sa_ctrl[0].r.part0[30] );
tran (\sa_ctrl[0][30] , \sa_ctrl[0].f.spare[25] );
tran (\sa_ctrl[0][29] , \sa_ctrl[0].r.part0[29] );
tran (\sa_ctrl[0][29] , \sa_ctrl[0].f.spare[24] );
tran (\sa_ctrl[0][28] , \sa_ctrl[0].r.part0[28] );
tran (\sa_ctrl[0][28] , \sa_ctrl[0].f.spare[23] );
tran (\sa_ctrl[0][27] , \sa_ctrl[0].r.part0[27] );
tran (\sa_ctrl[0][27] , \sa_ctrl[0].f.spare[22] );
tran (\sa_ctrl[0][26] , \sa_ctrl[0].r.part0[26] );
tran (\sa_ctrl[0][26] , \sa_ctrl[0].f.spare[21] );
tran (\sa_ctrl[0][25] , \sa_ctrl[0].r.part0[25] );
tran (\sa_ctrl[0][25] , \sa_ctrl[0].f.spare[20] );
tran (\sa_ctrl[0][24] , \sa_ctrl[0].r.part0[24] );
tran (\sa_ctrl[0][24] , \sa_ctrl[0].f.spare[19] );
tran (\sa_ctrl[0][23] , \sa_ctrl[0].r.part0[23] );
tran (\sa_ctrl[0][23] , \sa_ctrl[0].f.spare[18] );
tran (\sa_ctrl[0][22] , \sa_ctrl[0].r.part0[22] );
tran (\sa_ctrl[0][22] , \sa_ctrl[0].f.spare[17] );
tran (\sa_ctrl[0][21] , \sa_ctrl[0].r.part0[21] );
tran (\sa_ctrl[0][21] , \sa_ctrl[0].f.spare[16] );
tran (\sa_ctrl[0][20] , \sa_ctrl[0].r.part0[20] );
tran (\sa_ctrl[0][20] , \sa_ctrl[0].f.spare[15] );
tran (\sa_ctrl[0][19] , \sa_ctrl[0].r.part0[19] );
tran (\sa_ctrl[0][19] , \sa_ctrl[0].f.spare[14] );
tran (\sa_ctrl[0][18] , \sa_ctrl[0].r.part0[18] );
tran (\sa_ctrl[0][18] , \sa_ctrl[0].f.spare[13] );
tran (\sa_ctrl[0][17] , \sa_ctrl[0].r.part0[17] );
tran (\sa_ctrl[0][17] , \sa_ctrl[0].f.spare[12] );
tran (\sa_ctrl[0][16] , \sa_ctrl[0].r.part0[16] );
tran (\sa_ctrl[0][16] , \sa_ctrl[0].f.spare[11] );
tran (\sa_ctrl[0][15] , \sa_ctrl[0].r.part0[15] );
tran (\sa_ctrl[0][15] , \sa_ctrl[0].f.spare[10] );
tran (\sa_ctrl[0][14] , \sa_ctrl[0].r.part0[14] );
tran (\sa_ctrl[0][14] , \sa_ctrl[0].f.spare[9] );
tran (\sa_ctrl[0][13] , \sa_ctrl[0].r.part0[13] );
tran (\sa_ctrl[0][13] , \sa_ctrl[0].f.spare[8] );
tran (\sa_ctrl[0][12] , \sa_ctrl[0].r.part0[12] );
tran (\sa_ctrl[0][12] , \sa_ctrl[0].f.spare[7] );
tran (\sa_ctrl[0][11] , \sa_ctrl[0].r.part0[11] );
tran (\sa_ctrl[0][11] , \sa_ctrl[0].f.spare[6] );
tran (\sa_ctrl[0][10] , \sa_ctrl[0].r.part0[10] );
tran (\sa_ctrl[0][10] , \sa_ctrl[0].f.spare[5] );
tran (\sa_ctrl[0][9] , \sa_ctrl[0].r.part0[9] );
tran (\sa_ctrl[0][9] , \sa_ctrl[0].f.spare[4] );
tran (\sa_ctrl[0][8] , \sa_ctrl[0].r.part0[8] );
tran (\sa_ctrl[0][8] , \sa_ctrl[0].f.spare[3] );
tran (\sa_ctrl[0][7] , \sa_ctrl[0].r.part0[7] );
tran (\sa_ctrl[0][7] , \sa_ctrl[0].f.spare[2] );
tran (\sa_ctrl[0][6] , \sa_ctrl[0].r.part0[6] );
tran (\sa_ctrl[0][6] , \sa_ctrl[0].f.spare[1] );
tran (\sa_ctrl[0][5] , \sa_ctrl[0].r.part0[5] );
tran (\sa_ctrl[0][5] , \sa_ctrl[0].f.spare[0] );
tran (\sa_ctrl[0][4] , \sa_ctrl[0].r.part0[4] );
tran (\sa_ctrl[0][4] , \sa_ctrl[0].f.sa_event_sel[4] );
tran (\sa_ctrl[0][3] , \sa_ctrl[0].r.part0[3] );
tran (\sa_ctrl[0][3] , \sa_ctrl[0].f.sa_event_sel[3] );
tran (\sa_ctrl[0][2] , \sa_ctrl[0].r.part0[2] );
tran (\sa_ctrl[0][2] , \sa_ctrl[0].f.sa_event_sel[2] );
tran (\sa_ctrl[0][1] , \sa_ctrl[0].r.part0[1] );
tran (\sa_ctrl[0][1] , \sa_ctrl[0].f.sa_event_sel[1] );
tran (\sa_ctrl[0][0] , \sa_ctrl[0].r.part0[0] );
tran (\sa_ctrl[0][0] , \sa_ctrl[0].f.sa_event_sel[0] );
Q_BUF U0 ( .A(n1), .Z(rbus_ring_i[2]));
Q_BUF U1 ( .A(n1), .Z(rbus_ring_i[3]));
Q_BUF U2 ( .A(n1), .Z(rbus_ring_i[4]));
Q_BUF U3 ( .A(n1), .Z(rbus_ring_i[5]));
Q_BUF U4 ( .A(n1), .Z(rbus_ring_i[6]));
Q_BUF U5 ( .A(n1), .Z(rbus_ring_i[7]));
Q_BUF U6 ( .A(n1), .Z(rbus_ring_i[8]));
Q_BUF U7 ( .A(n1), .Z(rbus_ring_i[9]));
Q_BUF U8 ( .A(n1), .Z(rbus_ring_i[10]));
Q_BUF U9 ( .A(n1), .Z(rbus_ring_i[11]));
Q_BUF U10 ( .A(n1), .Z(rbus_ring_i[12]));
Q_BUF U11 ( .A(n1), .Z(rbus_ring_i[13]));
Q_BUF U12 ( .A(n1), .Z(rbus_ring_i[14]));
Q_BUF U13 ( .A(n1), .Z(rbus_ring_i[15]));
Q_BUF U14 ( .A(n1), .Z(rbus_ring_i[16]));
Q_BUF U15 ( .A(n1), .Z(rbus_ring_i[17]));
Q_BUF U16 ( .A(n1), .Z(rbus_ring_i[18]));
Q_BUF U17 ( .A(n1), .Z(rbus_ring_i[19]));
Q_BUF U18 ( .A(n1), .Z(rbus_ring_i[20]));
Q_BUF U19 ( .A(n1), .Z(rbus_ring_i[21]));
Q_BUF U20 ( .A(n1), .Z(rbus_ring_i[22]));
Q_BUF U21 ( .A(n1), .Z(rbus_ring_i[23]));
Q_BUF U22 ( .A(n1), .Z(rbus_ring_i[24]));
Q_BUF U23 ( .A(n1), .Z(rbus_ring_i[25]));
Q_BUF U24 ( .A(n1), .Z(rbus_ring_i[26]));
Q_BUF U25 ( .A(n1), .Z(rbus_ring_i[27]));
Q_BUF U26 ( .A(n1), .Z(rbus_ring_i[28]));
Q_BUF U27 ( .A(n1), .Z(rbus_ring_i[29]));
Q_BUF U28 ( .A(n1), .Z(rbus_ring_i[30]));
Q_BUF U29 ( .A(n1), .Z(rbus_ring_i[31]));
Q_BUF U30 ( .A(n1), .Z(rbus_ring_i[32]));
Q_BUF U31 ( .A(n1), .Z(rbus_ring_i[33]));
Q_BUF U32 ( .A(n1), .Z(rbus_ring_i[0]));
Q_BUF U33 ( .A(n1), .Z(rbus_ring_i[1]));
Q_BUF U34 ( .A(n1), .Z(_zy_simnet_cio_61[15]));
Q_BUF U35 ( .A(n1), .Z(_zy_simnet_cio_61[14]));
Q_BUF U36 ( .A(n2), .Z(_zy_simnet_cio_61[13]));
Q_BUF U37 ( .A(n2), .Z(_zy_simnet_cio_61[12]));
Q_BUF U38 ( .A(n2), .Z(_zy_simnet_cio_61[11]));
Q_BUF U39 ( .A(n1), .Z(_zy_simnet_cio_61[10]));
Q_BUF U40 ( .A(n2), .Z(_zy_simnet_cio_61[9]));
Q_BUF U41 ( .A(n1), .Z(_zy_simnet_cio_61[8]));
Q_BUF U42 ( .A(n1), .Z(_zy_simnet_cio_61[7]));
Q_BUF U43 ( .A(n1), .Z(_zy_simnet_cio_61[6]));
Q_BUF U44 ( .A(n2), .Z(_zy_simnet_cio_61[5]));
Q_BUF U45 ( .A(n1), .Z(_zy_simnet_cio_61[4]));
Q_BUF U46 ( .A(n1), .Z(_zy_simnet_cio_61[3]));
Q_BUF U47 ( .A(n1), .Z(_zy_simnet_cio_61[2]));
Q_BUF U48 ( .A(n1), .Z(_zy_simnet_cio_61[1]));
Q_BUF U49 ( .A(n1), .Z(_zy_simnet_cio_61[0]));
Q_BUF U50 ( .A(n1), .Z(_zy_simnet_cio_60[15]));
Q_BUF U51 ( .A(n1), .Z(_zy_simnet_cio_60[14]));
Q_BUF U52 ( .A(n1), .Z(_zy_simnet_cio_60[13]));
Q_BUF U53 ( .A(n1), .Z(_zy_simnet_cio_60[12]));
Q_BUF U54 ( .A(n1), .Z(_zy_simnet_cio_60[11]));
Q_BUF U55 ( .A(n1), .Z(_zy_simnet_cio_60[10]));
Q_BUF U56 ( .A(n1), .Z(_zy_simnet_cio_60[9]));
Q_BUF U57 ( .A(n1), .Z(_zy_simnet_cio_60[8]));
Q_BUF U58 ( .A(n1), .Z(_zy_simnet_cio_60[7]));
Q_BUF U59 ( .A(n1), .Z(_zy_simnet_cio_60[6]));
Q_BUF U60 ( .A(n1), .Z(_zy_simnet_cio_60[5]));
Q_BUF U61 ( .A(n1), .Z(_zy_simnet_cio_60[4]));
Q_BUF U62 ( .A(n1), .Z(_zy_simnet_cio_60[3]));
Q_BUF U63 ( .A(n1), .Z(_zy_simnet_cio_60[2]));
Q_BUF U64 ( .A(n1), .Z(_zy_simnet_cio_60[1]));
Q_BUF U65 ( .A(n1), .Z(_zy_simnet_cio_60[0]));
Q_BUF U66 ( .A(n2), .Z(kme_cddip3_ob_tready));
Q_BUF U67 ( .A(n2), .Z(kme_cddip2_ob_tready));
Q_BUF U68 ( .A(n2), .Z(kme_cddip1_ob_tready));
Q_BUF U69 ( .A(n2), .Z(kme_cddip0_ob_tready));
Q_BUF U70 ( .A(n2), .Z(kme_cceip3_ob_tready));
Q_BUF U71 ( .A(n2), .Z(kme_cceip2_ob_tready));
Q_BUF U72 ( .A(n2), .Z(kme_cceip1_ob_tready));
ixc_assign_2176 _zz_strnp_62 ( { \labels[7][271] , \labels[7][270] , 
	\labels[7][269] , \labels[7][268] , \labels[7][267] , 
	\labels[7][266] , \labels[7][265] , \labels[7][264] , 
	\labels[7][263] , \labels[7][262] , \labels[7][261] , 
	\labels[7][260] , \labels[7][259] , \labels[7][258] , 
	\labels[7][257] , \labels[7][256] , \labels[7][255] , 
	\labels[7][254] , \labels[7][253] , \labels[7][252] , 
	\labels[7][251] , \labels[7][250] , \labels[7][249] , 
	\labels[7][248] , \labels[7][247] , \labels[7][246] , 
	\labels[7][245] , \labels[7][244] , \labels[7][243] , 
	\labels[7][242] , \labels[7][241] , \labels[7][240] , 
	\labels[7][239] , \labels[7][238] , \labels[7][237] , 
	\labels[7][236] , \labels[7][235] , \labels[7][234] , 
	\labels[7][233] , \labels[7][232] , \labels[7][231] , 
	\labels[7][230] , \labels[7][229] , \labels[7][228] , 
	\labels[7][227] , \labels[7][226] , \labels[7][225] , 
	\labels[7][224] , \labels[7][223] , \labels[7][222] , 
	\labels[7][221] , \labels[7][220] , \labels[7][219] , 
	\labels[7][218] , \labels[7][217] , \labels[7][216] , 
	\labels[7][215] , \labels[7][214] , \labels[7][213] , 
	\labels[7][212] , \labels[7][211] , \labels[7][210] , 
	\labels[7][209] , \labels[7][208] , \labels[7][207] , 
	\labels[7][206] , \labels[7][205] , \labels[7][204] , 
	\labels[7][203] , \labels[7][202] , \labels[7][201] , 
	\labels[7][200] , \labels[7][199] , \labels[7][198] , 
	\labels[7][197] , \labels[7][196] , \labels[7][195] , 
	\labels[7][194] , \labels[7][193] , \labels[7][192] , 
	\labels[7][191] , \labels[7][190] , \labels[7][189] , 
	\labels[7][188] , \labels[7][187] , \labels[7][186] , 
	\labels[7][185] , \labels[7][184] , \labels[7][183] , 
	\labels[7][182] , \labels[7][181] , \labels[7][180] , 
	\labels[7][179] , \labels[7][178] , \labels[7][177] , 
	\labels[7][176] , \labels[7][175] , \labels[7][174] , 
	\labels[7][173] , \labels[7][172] , \labels[7][171] , 
	\labels[7][170] , \labels[7][169] , \labels[7][168] , 
	\labels[7][167] , \labels[7][166] , \labels[7][165] , 
	\labels[7][164] , \labels[7][163] , \labels[7][162] , 
	\labels[7][161] , \labels[7][160] , \labels[7][159] , 
	\labels[7][158] , \labels[7][157] , \labels[7][156] , 
	\labels[7][155] , \labels[7][154] , \labels[7][153] , 
	\labels[7][152] , \labels[7][151] , \labels[7][150] , 
	\labels[7][149] , \labels[7][148] , \labels[7][147] , 
	\labels[7][146] , \labels[7][145] , \labels[7][144] , 
	\labels[7][143] , \labels[7][142] , \labels[7][141] , 
	\labels[7][140] , \labels[7][139] , \labels[7][138] , 
	\labels[7][137] , \labels[7][136] , \labels[7][135] , 
	\labels[7][134] , \labels[7][133] , \labels[7][132] , 
	\labels[7][131] , \labels[7][130] , \labels[7][129] , 
	\labels[7][128] , \labels[7][127] , \labels[7][126] , 
	\labels[7][125] , \labels[7][124] , \labels[7][123] , 
	\labels[7][122] , \labels[7][121] , \labels[7][120] , 
	\labels[7][119] , \labels[7][118] , \labels[7][117] , 
	\labels[7][116] , \labels[7][115] , \labels[7][114] , 
	\labels[7][113] , \labels[7][112] , \labels[7][111] , 
	\labels[7][110] , \labels[7][109] , \labels[7][108] , 
	\labels[7][107] , \labels[7][106] , \labels[7][105] , 
	\labels[7][104] , \labels[7][103] , \labels[7][102] , 
	\labels[7][101] , \labels[7][100] , \labels[7][99] , \labels[7][98] , 
	\labels[7][97] , \labels[7][96] , \labels[7][95] , \labels[7][94] , 
	\labels[7][93] , \labels[7][92] , \labels[7][91] , \labels[7][90] , 
	\labels[7][89] , \labels[7][88] , \labels[7][87] , \labels[7][86] , 
	\labels[7][85] , \labels[7][84] , \labels[7][83] , \labels[7][82] , 
	\labels[7][81] , \labels[7][80] , \labels[7][79] , \labels[7][78] , 
	\labels[7][77] , \labels[7][76] , \labels[7][75] , \labels[7][74] , 
	\labels[7][73] , \labels[7][72] , \labels[7][71] , \labels[7][70] , 
	\labels[7][69] , \labels[7][68] , \labels[7][67] , \labels[7][66] , 
	\labels[7][65] , \labels[7][64] , \labels[7][63] , \labels[7][62] , 
	\labels[7][61] , \labels[7][60] , \labels[7][59] , \labels[7][58] , 
	\labels[7][57] , \labels[7][56] , \labels[7][55] , \labels[7][54] , 
	\labels[7][53] , \labels[7][52] , \labels[7][51] , \labels[7][50] , 
	\labels[7][49] , \labels[7][48] , \labels[7][47] , \labels[7][46] , 
	\labels[7][45] , \labels[7][44] , \labels[7][43] , \labels[7][42] , 
	\labels[7][41] , \labels[7][40] , \labels[7][39] , \labels[7][38] , 
	\labels[7][37] , \labels[7][36] , \labels[7][35] , \labels[7][34] , 
	\labels[7][33] , \labels[7][32] , \labels[7][31] , \labels[7][30] , 
	\labels[7][29] , \labels[7][28] , \labels[7][27] , \labels[7][26] , 
	\labels[7][25] , \labels[7][24] , \labels[7][23] , \labels[7][22] , 
	\labels[7][21] , \labels[7][20] , \labels[7][19] , \labels[7][18] , 
	\labels[7][17] , \labels[7][16] , \labels[7][15] , \labels[7][14] , 
	\labels[7][13] , \labels[7][12] , \labels[7][11] , \labels[7][10] , 
	\labels[7][9] , \labels[7][8] , \labels[7][7] , \labels[7][6] , 
	\labels[7][5] , \labels[7][4] , \labels[7][3] , \labels[7][2] , 
	\labels[7][1] , \labels[7][0] , \labels[6][271] , \labels[6][270] , 
	\labels[6][269] , \labels[6][268] , \labels[6][267] , 
	\labels[6][266] , \labels[6][265] , \labels[6][264] , 
	\labels[6][263] , \labels[6][262] , \labels[6][261] , 
	\labels[6][260] , \labels[6][259] , \labels[6][258] , 
	\labels[6][257] , \labels[6][256] , \labels[6][255] , 
	\labels[6][254] , \labels[6][253] , \labels[6][252] , 
	\labels[6][251] , \labels[6][250] , \labels[6][249] , 
	\labels[6][248] , \labels[6][247] , \labels[6][246] , 
	\labels[6][245] , \labels[6][244] , \labels[6][243] , 
	\labels[6][242] , \labels[6][241] , \labels[6][240] , 
	\labels[6][239] , \labels[6][238] , \labels[6][237] , 
	\labels[6][236] , \labels[6][235] , \labels[6][234] , 
	\labels[6][233] , \labels[6][232] , \labels[6][231] , 
	\labels[6][230] , \labels[6][229] , \labels[6][228] , 
	\labels[6][227] , \labels[6][226] , \labels[6][225] , 
	\labels[6][224] , \labels[6][223] , \labels[6][222] , 
	\labels[6][221] , \labels[6][220] , \labels[6][219] , 
	\labels[6][218] , \labels[6][217] , \labels[6][216] , 
	\labels[6][215] , \labels[6][214] , \labels[6][213] , 
	\labels[6][212] , \labels[6][211] , \labels[6][210] , 
	\labels[6][209] , \labels[6][208] , \labels[6][207] , 
	\labels[6][206] , \labels[6][205] , \labels[6][204] , 
	\labels[6][203] , \labels[6][202] , \labels[6][201] , 
	\labels[6][200] , \labels[6][199] , \labels[6][198] , 
	\labels[6][197] , \labels[6][196] , \labels[6][195] , 
	\labels[6][194] , \labels[6][193] , \labels[6][192] , 
	\labels[6][191] , \labels[6][190] , \labels[6][189] , 
	\labels[6][188] , \labels[6][187] , \labels[6][186] , 
	\labels[6][185] , \labels[6][184] , \labels[6][183] , 
	\labels[6][182] , \labels[6][181] , \labels[6][180] , 
	\labels[6][179] , \labels[6][178] , \labels[6][177] , 
	\labels[6][176] , \labels[6][175] , \labels[6][174] , 
	\labels[6][173] , \labels[6][172] , \labels[6][171] , 
	\labels[6][170] , \labels[6][169] , \labels[6][168] , 
	\labels[6][167] , \labels[6][166] , \labels[6][165] , 
	\labels[6][164] , \labels[6][163] , \labels[6][162] , 
	\labels[6][161] , \labels[6][160] , \labels[6][159] , 
	\labels[6][158] , \labels[6][157] , \labels[6][156] , 
	\labels[6][155] , \labels[6][154] , \labels[6][153] , 
	\labels[6][152] , \labels[6][151] , \labels[6][150] , 
	\labels[6][149] , \labels[6][148] , \labels[6][147] , 
	\labels[6][146] , \labels[6][145] , \labels[6][144] , 
	\labels[6][143] , \labels[6][142] , \labels[6][141] , 
	\labels[6][140] , \labels[6][139] , \labels[6][138] , 
	\labels[6][137] , \labels[6][136] , \labels[6][135] , 
	\labels[6][134] , \labels[6][133] , \labels[6][132] , 
	\labels[6][131] , \labels[6][130] , \labels[6][129] , 
	\labels[6][128] , \labels[6][127] , \labels[6][126] , 
	\labels[6][125] , \labels[6][124] , \labels[6][123] , 
	\labels[6][122] , \labels[6][121] , \labels[6][120] , 
	\labels[6][119] , \labels[6][118] , \labels[6][117] , 
	\labels[6][116] , \labels[6][115] , \labels[6][114] , 
	\labels[6][113] , \labels[6][112] , \labels[6][111] , 
	\labels[6][110] , \labels[6][109] , \labels[6][108] , 
	\labels[6][107] , \labels[6][106] , \labels[6][105] , 
	\labels[6][104] , \labels[6][103] , \labels[6][102] , 
	\labels[6][101] , \labels[6][100] , \labels[6][99] , \labels[6][98] , 
	\labels[6][97] , \labels[6][96] , \labels[6][95] , \labels[6][94] , 
	\labels[6][93] , \labels[6][92] , \labels[6][91] , \labels[6][90] , 
	\labels[6][89] , \labels[6][88] , \labels[6][87] , \labels[6][86] , 
	\labels[6][85] , \labels[6][84] , \labels[6][83] , \labels[6][82] , 
	\labels[6][81] , \labels[6][80] , \labels[6][79] , \labels[6][78] , 
	\labels[6][77] , \labels[6][76] , \labels[6][75] , \labels[6][74] , 
	\labels[6][73] , \labels[6][72] , \labels[6][71] , \labels[6][70] , 
	\labels[6][69] , \labels[6][68] , \labels[6][67] , \labels[6][66] , 
	\labels[6][65] , \labels[6][64] , \labels[6][63] , \labels[6][62] , 
	\labels[6][61] , \labels[6][60] , \labels[6][59] , \labels[6][58] , 
	\labels[6][57] , \labels[6][56] , \labels[6][55] , \labels[6][54] , 
	\labels[6][53] , \labels[6][52] , \labels[6][51] , \labels[6][50] , 
	\labels[6][49] , \labels[6][48] , \labels[6][47] , \labels[6][46] , 
	\labels[6][45] , \labels[6][44] , \labels[6][43] , \labels[6][42] , 
	\labels[6][41] , \labels[6][40] , \labels[6][39] , \labels[6][38] , 
	\labels[6][37] , \labels[6][36] , \labels[6][35] , \labels[6][34] , 
	\labels[6][33] , \labels[6][32] , \labels[6][31] , \labels[6][30] , 
	\labels[6][29] , \labels[6][28] , \labels[6][27] , \labels[6][26] , 
	\labels[6][25] , \labels[6][24] , \labels[6][23] , \labels[6][22] , 
	\labels[6][21] , \labels[6][20] , \labels[6][19] , \labels[6][18] , 
	\labels[6][17] , \labels[6][16] , \labels[6][15] , \labels[6][14] , 
	\labels[6][13] , \labels[6][12] , \labels[6][11] , \labels[6][10] , 
	\labels[6][9] , \labels[6][8] , \labels[6][7] , \labels[6][6] , 
	\labels[6][5] , \labels[6][4] , \labels[6][3] , \labels[6][2] , 
	\labels[6][1] , \labels[6][0] , \labels[5][271] , \labels[5][270] , 
	\labels[5][269] , \labels[5][268] , \labels[5][267] , 
	\labels[5][266] , \labels[5][265] , \labels[5][264] , 
	\labels[5][263] , \labels[5][262] , \labels[5][261] , 
	\labels[5][260] , \labels[5][259] , \labels[5][258] , 
	\labels[5][257] , \labels[5][256] , \labels[5][255] , 
	\labels[5][254] , \labels[5][253] , \labels[5][252] , 
	\labels[5][251] , \labels[5][250] , \labels[5][249] , 
	\labels[5][248] , \labels[5][247] , \labels[5][246] , 
	\labels[5][245] , \labels[5][244] , \labels[5][243] , 
	\labels[5][242] , \labels[5][241] , \labels[5][240] , 
	\labels[5][239] , \labels[5][238] , \labels[5][237] , 
	\labels[5][236] , \labels[5][235] , \labels[5][234] , 
	\labels[5][233] , \labels[5][232] , \labels[5][231] , 
	\labels[5][230] , \labels[5][229] , \labels[5][228] , 
	\labels[5][227] , \labels[5][226] , \labels[5][225] , 
	\labels[5][224] , \labels[5][223] , \labels[5][222] , 
	\labels[5][221] , \labels[5][220] , \labels[5][219] , 
	\labels[5][218] , \labels[5][217] , \labels[5][216] , 
	\labels[5][215] , \labels[5][214] , \labels[5][213] , 
	\labels[5][212] , \labels[5][211] , \labels[5][210] , 
	\labels[5][209] , \labels[5][208] , \labels[5][207] , 
	\labels[5][206] , \labels[5][205] , \labels[5][204] , 
	\labels[5][203] , \labels[5][202] , \labels[5][201] , 
	\labels[5][200] , \labels[5][199] , \labels[5][198] , 
	\labels[5][197] , \labels[5][196] , \labels[5][195] , 
	\labels[5][194] , \labels[5][193] , \labels[5][192] , 
	\labels[5][191] , \labels[5][190] , \labels[5][189] , 
	\labels[5][188] , \labels[5][187] , \labels[5][186] , 
	\labels[5][185] , \labels[5][184] , \labels[5][183] , 
	\labels[5][182] , \labels[5][181] , \labels[5][180] , 
	\labels[5][179] , \labels[5][178] , \labels[5][177] , 
	\labels[5][176] , \labels[5][175] , \labels[5][174] , 
	\labels[5][173] , \labels[5][172] , \labels[5][171] , 
	\labels[5][170] , \labels[5][169] , \labels[5][168] , 
	\labels[5][167] , \labels[5][166] , \labels[5][165] , 
	\labels[5][164] , \labels[5][163] , \labels[5][162] , 
	\labels[5][161] , \labels[5][160] , \labels[5][159] , 
	\labels[5][158] , \labels[5][157] , \labels[5][156] , 
	\labels[5][155] , \labels[5][154] , \labels[5][153] , 
	\labels[5][152] , \labels[5][151] , \labels[5][150] , 
	\labels[5][149] , \labels[5][148] , \labels[5][147] , 
	\labels[5][146] , \labels[5][145] , \labels[5][144] , 
	\labels[5][143] , \labels[5][142] , \labels[5][141] , 
	\labels[5][140] , \labels[5][139] , \labels[5][138] , 
	\labels[5][137] , \labels[5][136] , \labels[5][135] , 
	\labels[5][134] , \labels[5][133] , \labels[5][132] , 
	\labels[5][131] , \labels[5][130] , \labels[5][129] , 
	\labels[5][128] , \labels[5][127] , \labels[5][126] , 
	\labels[5][125] , \labels[5][124] , \labels[5][123] , 
	\labels[5][122] , \labels[5][121] , \labels[5][120] , 
	\labels[5][119] , \labels[5][118] , \labels[5][117] , 
	\labels[5][116] , \labels[5][115] , \labels[5][114] , 
	\labels[5][113] , \labels[5][112] , \labels[5][111] , 
	\labels[5][110] , \labels[5][109] , \labels[5][108] , 
	\labels[5][107] , \labels[5][106] , \labels[5][105] , 
	\labels[5][104] , \labels[5][103] , \labels[5][102] , 
	\labels[5][101] , \labels[5][100] , \labels[5][99] , \labels[5][98] , 
	\labels[5][97] , \labels[5][96] , \labels[5][95] , \labels[5][94] , 
	\labels[5][93] , \labels[5][92] , \labels[5][91] , \labels[5][90] , 
	\labels[5][89] , \labels[5][88] , \labels[5][87] , \labels[5][86] , 
	\labels[5][85] , \labels[5][84] , \labels[5][83] , \labels[5][82] , 
	\labels[5][81] , \labels[5][80] , \labels[5][79] , \labels[5][78] , 
	\labels[5][77] , \labels[5][76] , \labels[5][75] , \labels[5][74] , 
	\labels[5][73] , \labels[5][72] , \labels[5][71] , \labels[5][70] , 
	\labels[5][69] , \labels[5][68] , \labels[5][67] , \labels[5][66] , 
	\labels[5][65] , \labels[5][64] , \labels[5][63] , \labels[5][62] , 
	\labels[5][61] , \labels[5][60] , \labels[5][59] , \labels[5][58] , 
	\labels[5][57] , \labels[5][56] , \labels[5][55] , \labels[5][54] , 
	\labels[5][53] , \labels[5][52] , \labels[5][51] , \labels[5][50] , 
	\labels[5][49] , \labels[5][48] , \labels[5][47] , \labels[5][46] , 
	\labels[5][45] , \labels[5][44] , \labels[5][43] , \labels[5][42] , 
	\labels[5][41] , \labels[5][40] , \labels[5][39] , \labels[5][38] , 
	\labels[5][37] , \labels[5][36] , \labels[5][35] , \labels[5][34] , 
	\labels[5][33] , \labels[5][32] , \labels[5][31] , \labels[5][30] , 
	\labels[5][29] , \labels[5][28] , \labels[5][27] , \labels[5][26] , 
	\labels[5][25] , \labels[5][24] , \labels[5][23] , \labels[5][22] , 
	\labels[5][21] , \labels[5][20] , \labels[5][19] , \labels[5][18] , 
	\labels[5][17] , \labels[5][16] , \labels[5][15] , \labels[5][14] , 
	\labels[5][13] , \labels[5][12] , \labels[5][11] , \labels[5][10] , 
	\labels[5][9] , \labels[5][8] , \labels[5][7] , \labels[5][6] , 
	\labels[5][5] , \labels[5][4] , \labels[5][3] , \labels[5][2] , 
	\labels[5][1] , \labels[5][0] , \labels[4][271] , \labels[4][270] , 
	\labels[4][269] , \labels[4][268] , \labels[4][267] , 
	\labels[4][266] , \labels[4][265] , \labels[4][264] , 
	\labels[4][263] , \labels[4][262] , \labels[4][261] , 
	\labels[4][260] , \labels[4][259] , \labels[4][258] , 
	\labels[4][257] , \labels[4][256] , \labels[4][255] , 
	\labels[4][254] , \labels[4][253] , \labels[4][252] , 
	\labels[4][251] , \labels[4][250] , \labels[4][249] , 
	\labels[4][248] , \labels[4][247] , \labels[4][246] , 
	\labels[4][245] , \labels[4][244] , \labels[4][243] , 
	\labels[4][242] , \labels[4][241] , \labels[4][240] , 
	\labels[4][239] , \labels[4][238] , \labels[4][237] , 
	\labels[4][236] , \labels[4][235] , \labels[4][234] , 
	\labels[4][233] , \labels[4][232] , \labels[4][231] , 
	\labels[4][230] , \labels[4][229] , \labels[4][228] , 
	\labels[4][227] , \labels[4][226] , \labels[4][225] , 
	\labels[4][224] , \labels[4][223] , \labels[4][222] , 
	\labels[4][221] , \labels[4][220] , \labels[4][219] , 
	\labels[4][218] , \labels[4][217] , \labels[4][216] , 
	\labels[4][215] , \labels[4][214] , \labels[4][213] , 
	\labels[4][212] , \labels[4][211] , \labels[4][210] , 
	\labels[4][209] , \labels[4][208] , \labels[4][207] , 
	\labels[4][206] , \labels[4][205] , \labels[4][204] , 
	\labels[4][203] , \labels[4][202] , \labels[4][201] , 
	\labels[4][200] , \labels[4][199] , \labels[4][198] , 
	\labels[4][197] , \labels[4][196] , \labels[4][195] , 
	\labels[4][194] , \labels[4][193] , \labels[4][192] , 
	\labels[4][191] , \labels[4][190] , \labels[4][189] , 
	\labels[4][188] , \labels[4][187] , \labels[4][186] , 
	\labels[4][185] , \labels[4][184] , \labels[4][183] , 
	\labels[4][182] , \labels[4][181] , \labels[4][180] , 
	\labels[4][179] , \labels[4][178] , \labels[4][177] , 
	\labels[4][176] , \labels[4][175] , \labels[4][174] , 
	\labels[4][173] , \labels[4][172] , \labels[4][171] , 
	\labels[4][170] , \labels[4][169] , \labels[4][168] , 
	\labels[4][167] , \labels[4][166] , \labels[4][165] , 
	\labels[4][164] , \labels[4][163] , \labels[4][162] , 
	\labels[4][161] , \labels[4][160] , \labels[4][159] , 
	\labels[4][158] , \labels[4][157] , \labels[4][156] , 
	\labels[4][155] , \labels[4][154] , \labels[4][153] , 
	\labels[4][152] , \labels[4][151] , \labels[4][150] , 
	\labels[4][149] , \labels[4][148] , \labels[4][147] , 
	\labels[4][146] , \labels[4][145] , \labels[4][144] , 
	\labels[4][143] , \labels[4][142] , \labels[4][141] , 
	\labels[4][140] , \labels[4][139] , \labels[4][138] , 
	\labels[4][137] , \labels[4][136] , \labels[4][135] , 
	\labels[4][134] , \labels[4][133] , \labels[4][132] , 
	\labels[4][131] , \labels[4][130] , \labels[4][129] , 
	\labels[4][128] , \labels[4][127] , \labels[4][126] , 
	\labels[4][125] , \labels[4][124] , \labels[4][123] , 
	\labels[4][122] , \labels[4][121] , \labels[4][120] , 
	\labels[4][119] , \labels[4][118] , \labels[4][117] , 
	\labels[4][116] , \labels[4][115] , \labels[4][114] , 
	\labels[4][113] , \labels[4][112] , \labels[4][111] , 
	\labels[4][110] , \labels[4][109] , \labels[4][108] , 
	\labels[4][107] , \labels[4][106] , \labels[4][105] , 
	\labels[4][104] , \labels[4][103] , \labels[4][102] , 
	\labels[4][101] , \labels[4][100] , \labels[4][99] , \labels[4][98] , 
	\labels[4][97] , \labels[4][96] , \labels[4][95] , \labels[4][94] , 
	\labels[4][93] , \labels[4][92] , \labels[4][91] , \labels[4][90] , 
	\labels[4][89] , \labels[4][88] , \labels[4][87] , \labels[4][86] , 
	\labels[4][85] , \labels[4][84] , \labels[4][83] , \labels[4][82] , 
	\labels[4][81] , \labels[4][80] , \labels[4][79] , \labels[4][78] , 
	\labels[4][77] , \labels[4][76] , \labels[4][75] , \labels[4][74] , 
	\labels[4][73] , \labels[4][72] , \labels[4][71] , \labels[4][70] , 
	\labels[4][69] , \labels[4][68] , \labels[4][67] , \labels[4][66] , 
	\labels[4][65] , \labels[4][64] , \labels[4][63] , \labels[4][62] , 
	\labels[4][61] , \labels[4][60] , \labels[4][59] , \labels[4][58] , 
	\labels[4][57] , \labels[4][56] , \labels[4][55] , \labels[4][54] , 
	\labels[4][53] , \labels[4][52] , \labels[4][51] , \labels[4][50] , 
	\labels[4][49] , \labels[4][48] , \labels[4][47] , \labels[4][46] , 
	\labels[4][45] , \labels[4][44] , \labels[4][43] , \labels[4][42] , 
	\labels[4][41] , \labels[4][40] , \labels[4][39] , \labels[4][38] , 
	\labels[4][37] , \labels[4][36] , \labels[4][35] , \labels[4][34] , 
	\labels[4][33] , \labels[4][32] , \labels[4][31] , \labels[4][30] , 
	\labels[4][29] , \labels[4][28] , \labels[4][27] , \labels[4][26] , 
	\labels[4][25] , \labels[4][24] , \labels[4][23] , \labels[4][22] , 
	\labels[4][21] , \labels[4][20] , \labels[4][19] , \labels[4][18] , 
	\labels[4][17] , \labels[4][16] , \labels[4][15] , \labels[4][14] , 
	\labels[4][13] , \labels[4][12] , \labels[4][11] , \labels[4][10] , 
	\labels[4][9] , \labels[4][8] , \labels[4][7] , \labels[4][6] , 
	\labels[4][5] , \labels[4][4] , \labels[4][3] , \labels[4][2] , 
	\labels[4][1] , \labels[4][0] , \labels[3][271] , \labels[3][270] , 
	\labels[3][269] , \labels[3][268] , \labels[3][267] , 
	\labels[3][266] , \labels[3][265] , \labels[3][264] , 
	\labels[3][263] , \labels[3][262] , \labels[3][261] , 
	\labels[3][260] , \labels[3][259] , \labels[3][258] , 
	\labels[3][257] , \labels[3][256] , \labels[3][255] , 
	\labels[3][254] , \labels[3][253] , \labels[3][252] , 
	\labels[3][251] , \labels[3][250] , \labels[3][249] , 
	\labels[3][248] , \labels[3][247] , \labels[3][246] , 
	\labels[3][245] , \labels[3][244] , \labels[3][243] , 
	\labels[3][242] , \labels[3][241] , \labels[3][240] , 
	\labels[3][239] , \labels[3][238] , \labels[3][237] , 
	\labels[3][236] , \labels[3][235] , \labels[3][234] , 
	\labels[3][233] , \labels[3][232] , \labels[3][231] , 
	\labels[3][230] , \labels[3][229] , \labels[3][228] , 
	\labels[3][227] , \labels[3][226] , \labels[3][225] , 
	\labels[3][224] , \labels[3][223] , \labels[3][222] , 
	\labels[3][221] , \labels[3][220] , \labels[3][219] , 
	\labels[3][218] , \labels[3][217] , \labels[3][216] , 
	\labels[3][215] , \labels[3][214] , \labels[3][213] , 
	\labels[3][212] , \labels[3][211] , \labels[3][210] , 
	\labels[3][209] , \labels[3][208] , \labels[3][207] , 
	\labels[3][206] , \labels[3][205] , \labels[3][204] , 
	\labels[3][203] , \labels[3][202] , \labels[3][201] , 
	\labels[3][200] , \labels[3][199] , \labels[3][198] , 
	\labels[3][197] , \labels[3][196] , \labels[3][195] , 
	\labels[3][194] , \labels[3][193] , \labels[3][192] , 
	\labels[3][191] , \labels[3][190] , \labels[3][189] , 
	\labels[3][188] , \labels[3][187] , \labels[3][186] , 
	\labels[3][185] , \labels[3][184] , \labels[3][183] , 
	\labels[3][182] , \labels[3][181] , \labels[3][180] , 
	\labels[3][179] , \labels[3][178] , \labels[3][177] , 
	\labels[3][176] , \labels[3][175] , \labels[3][174] , 
	\labels[3][173] , \labels[3][172] , \labels[3][171] , 
	\labels[3][170] , \labels[3][169] , \labels[3][168] , 
	\labels[3][167] , \labels[3][166] , \labels[3][165] , 
	\labels[3][164] , \labels[3][163] , \labels[3][162] , 
	\labels[3][161] , \labels[3][160] , \labels[3][159] , 
	\labels[3][158] , \labels[3][157] , \labels[3][156] , 
	\labels[3][155] , \labels[3][154] , \labels[3][153] , 
	\labels[3][152] , \labels[3][151] , \labels[3][150] , 
	\labels[3][149] , \labels[3][148] , \labels[3][147] , 
	\labels[3][146] , \labels[3][145] , \labels[3][144] , 
	\labels[3][143] , \labels[3][142] , \labels[3][141] , 
	\labels[3][140] , \labels[3][139] , \labels[3][138] , 
	\labels[3][137] , \labels[3][136] , \labels[3][135] , 
	\labels[3][134] , \labels[3][133] , \labels[3][132] , 
	\labels[3][131] , \labels[3][130] , \labels[3][129] , 
	\labels[3][128] , \labels[3][127] , \labels[3][126] , 
	\labels[3][125] , \labels[3][124] , \labels[3][123] , 
	\labels[3][122] , \labels[3][121] , \labels[3][120] , 
	\labels[3][119] , \labels[3][118] , \labels[3][117] , 
	\labels[3][116] , \labels[3][115] , \labels[3][114] , 
	\labels[3][113] , \labels[3][112] , \labels[3][111] , 
	\labels[3][110] , \labels[3][109] , \labels[3][108] , 
	\labels[3][107] , \labels[3][106] , \labels[3][105] , 
	\labels[3][104] , \labels[3][103] , \labels[3][102] , 
	\labels[3][101] , \labels[3][100] , \labels[3][99] , \labels[3][98] , 
	\labels[3][97] , \labels[3][96] , \labels[3][95] , \labels[3][94] , 
	\labels[3][93] , \labels[3][92] , \labels[3][91] , \labels[3][90] , 
	\labels[3][89] , \labels[3][88] , \labels[3][87] , \labels[3][86] , 
	\labels[3][85] , \labels[3][84] , \labels[3][83] , \labels[3][82] , 
	\labels[3][81] , \labels[3][80] , \labels[3][79] , \labels[3][78] , 
	\labels[3][77] , \labels[3][76] , \labels[3][75] , \labels[3][74] , 
	\labels[3][73] , \labels[3][72] , \labels[3][71] , \labels[3][70] , 
	\labels[3][69] , \labels[3][68] , \labels[3][67] , \labels[3][66] , 
	\labels[3][65] , \labels[3][64] , \labels[3][63] , \labels[3][62] , 
	\labels[3][61] , \labels[3][60] , \labels[3][59] , \labels[3][58] , 
	\labels[3][57] , \labels[3][56] , \labels[3][55] , \labels[3][54] , 
	\labels[3][53] , \labels[3][52] , \labels[3][51] , \labels[3][50] , 
	\labels[3][49] , \labels[3][48] , \labels[3][47] , \labels[3][46] , 
	\labels[3][45] , \labels[3][44] , \labels[3][43] , \labels[3][42] , 
	\labels[3][41] , \labels[3][40] , \labels[3][39] , \labels[3][38] , 
	\labels[3][37] , \labels[3][36] , \labels[3][35] , \labels[3][34] , 
	\labels[3][33] , \labels[3][32] , \labels[3][31] , \labels[3][30] , 
	\labels[3][29] , \labels[3][28] , \labels[3][27] , \labels[3][26] , 
	\labels[3][25] , \labels[3][24] , \labels[3][23] , \labels[3][22] , 
	\labels[3][21] , \labels[3][20] , \labels[3][19] , \labels[3][18] , 
	\labels[3][17] , \labels[3][16] , \labels[3][15] , \labels[3][14] , 
	\labels[3][13] , \labels[3][12] , \labels[3][11] , \labels[3][10] , 
	\labels[3][9] , \labels[3][8] , \labels[3][7] , \labels[3][6] , 
	\labels[3][5] , \labels[3][4] , \labels[3][3] , \labels[3][2] , 
	\labels[3][1] , \labels[3][0] , \labels[2][271] , \labels[2][270] , 
	\labels[2][269] , \labels[2][268] , \labels[2][267] , 
	\labels[2][266] , \labels[2][265] , \labels[2][264] , 
	\labels[2][263] , \labels[2][262] , \labels[2][261] , 
	\labels[2][260] , \labels[2][259] , \labels[2][258] , 
	\labels[2][257] , \labels[2][256] , \labels[2][255] , 
	\labels[2][254] , \labels[2][253] , \labels[2][252] , 
	\labels[2][251] , \labels[2][250] , \labels[2][249] , 
	\labels[2][248] , \labels[2][247] , \labels[2][246] , 
	\labels[2][245] , \labels[2][244] , \labels[2][243] , 
	\labels[2][242] , \labels[2][241] , \labels[2][240] , 
	\labels[2][239] , \labels[2][238] , \labels[2][237] , 
	\labels[2][236] , \labels[2][235] , \labels[2][234] , 
	\labels[2][233] , \labels[2][232] , \labels[2][231] , 
	\labels[2][230] , \labels[2][229] , \labels[2][228] , 
	\labels[2][227] , \labels[2][226] , \labels[2][225] , 
	\labels[2][224] , \labels[2][223] , \labels[2][222] , 
	\labels[2][221] , \labels[2][220] , \labels[2][219] , 
	\labels[2][218] , \labels[2][217] , \labels[2][216] , 
	\labels[2][215] , \labels[2][214] , \labels[2][213] , 
	\labels[2][212] , \labels[2][211] , \labels[2][210] , 
	\labels[2][209] , \labels[2][208] , \labels[2][207] , 
	\labels[2][206] , \labels[2][205] , \labels[2][204] , 
	\labels[2][203] , \labels[2][202] , \labels[2][201] , 
	\labels[2][200] , \labels[2][199] , \labels[2][198] , 
	\labels[2][197] , \labels[2][196] , \labels[2][195] , 
	\labels[2][194] , \labels[2][193] , \labels[2][192] , 
	\labels[2][191] , \labels[2][190] , \labels[2][189] , 
	\labels[2][188] , \labels[2][187] , \labels[2][186] , 
	\labels[2][185] , \labels[2][184] , \labels[2][183] , 
	\labels[2][182] , \labels[2][181] , \labels[2][180] , 
	\labels[2][179] , \labels[2][178] , \labels[2][177] , 
	\labels[2][176] , \labels[2][175] , \labels[2][174] , 
	\labels[2][173] , \labels[2][172] , \labels[2][171] , 
	\labels[2][170] , \labels[2][169] , \labels[2][168] , 
	\labels[2][167] , \labels[2][166] , \labels[2][165] , 
	\labels[2][164] , \labels[2][163] , \labels[2][162] , 
	\labels[2][161] , \labels[2][160] , \labels[2][159] , 
	\labels[2][158] , \labels[2][157] , \labels[2][156] , 
	\labels[2][155] , \labels[2][154] , \labels[2][153] , 
	\labels[2][152] , \labels[2][151] , \labels[2][150] , 
	\labels[2][149] , \labels[2][148] , \labels[2][147] , 
	\labels[2][146] , \labels[2][145] , \labels[2][144] , 
	\labels[2][143] , \labels[2][142] , \labels[2][141] , 
	\labels[2][140] , \labels[2][139] , \labels[2][138] , 
	\labels[2][137] , \labels[2][136] , \labels[2][135] , 
	\labels[2][134] , \labels[2][133] , \labels[2][132] , 
	\labels[2][131] , \labels[2][130] , \labels[2][129] , 
	\labels[2][128] , \labels[2][127] , \labels[2][126] , 
	\labels[2][125] , \labels[2][124] , \labels[2][123] , 
	\labels[2][122] , \labels[2][121] , \labels[2][120] , 
	\labels[2][119] , \labels[2][118] , \labels[2][117] , 
	\labels[2][116] , \labels[2][115] , \labels[2][114] , 
	\labels[2][113] , \labels[2][112] , \labels[2][111] , 
	\labels[2][110] , \labels[2][109] , \labels[2][108] , 
	\labels[2][107] , \labels[2][106] , \labels[2][105] , 
	\labels[2][104] , \labels[2][103] , \labels[2][102] , 
	\labels[2][101] , \labels[2][100] , \labels[2][99] , \labels[2][98] , 
	\labels[2][97] , \labels[2][96] , \labels[2][95] , \labels[2][94] , 
	\labels[2][93] , \labels[2][92] , \labels[2][91] , \labels[2][90] , 
	\labels[2][89] , \labels[2][88] , \labels[2][87] , \labels[2][86] , 
	\labels[2][85] , \labels[2][84] , \labels[2][83] , \labels[2][82] , 
	\labels[2][81] , \labels[2][80] , \labels[2][79] , \labels[2][78] , 
	\labels[2][77] , \labels[2][76] , \labels[2][75] , \labels[2][74] , 
	\labels[2][73] , \labels[2][72] , \labels[2][71] , \labels[2][70] , 
	\labels[2][69] , \labels[2][68] , \labels[2][67] , \labels[2][66] , 
	\labels[2][65] , \labels[2][64] , \labels[2][63] , \labels[2][62] , 
	\labels[2][61] , \labels[2][60] , \labels[2][59] , \labels[2][58] , 
	\labels[2][57] , \labels[2][56] , \labels[2][55] , \labels[2][54] , 
	\labels[2][53] , \labels[2][52] , \labels[2][51] , \labels[2][50] , 
	\labels[2][49] , \labels[2][48] , \labels[2][47] , \labels[2][46] , 
	\labels[2][45] , \labels[2][44] , \labels[2][43] , \labels[2][42] , 
	\labels[2][41] , \labels[2][40] , \labels[2][39] , \labels[2][38] , 
	\labels[2][37] , \labels[2][36] , \labels[2][35] , \labels[2][34] , 
	\labels[2][33] , \labels[2][32] , \labels[2][31] , \labels[2][30] , 
	\labels[2][29] , \labels[2][28] , \labels[2][27] , \labels[2][26] , 
	\labels[2][25] , \labels[2][24] , \labels[2][23] , \labels[2][22] , 
	\labels[2][21] , \labels[2][20] , \labels[2][19] , \labels[2][18] , 
	\labels[2][17] , \labels[2][16] , \labels[2][15] , \labels[2][14] , 
	\labels[2][13] , \labels[2][12] , \labels[2][11] , \labels[2][10] , 
	\labels[2][9] , \labels[2][8] , \labels[2][7] , \labels[2][6] , 
	\labels[2][5] , \labels[2][4] , \labels[2][3] , \labels[2][2] , 
	\labels[2][1] , \labels[2][0] , \labels[1][271] , \labels[1][270] , 
	\labels[1][269] , \labels[1][268] , \labels[1][267] , 
	\labels[1][266] , \labels[1][265] , \labels[1][264] , 
	\labels[1][263] , \labels[1][262] , \labels[1][261] , 
	\labels[1][260] , \labels[1][259] , \labels[1][258] , 
	\labels[1][257] , \labels[1][256] , \labels[1][255] , 
	\labels[1][254] , \labels[1][253] , \labels[1][252] , 
	\labels[1][251] , \labels[1][250] , \labels[1][249] , 
	\labels[1][248] , \labels[1][247] , \labels[1][246] , 
	\labels[1][245] , \labels[1][244] , \labels[1][243] , 
	\labels[1][242] , \labels[1][241] , \labels[1][240] , 
	\labels[1][239] , \labels[1][238] , \labels[1][237] , 
	\labels[1][236] , \labels[1][235] , \labels[1][234] , 
	\labels[1][233] , \labels[1][232] , \labels[1][231] , 
	\labels[1][230] , \labels[1][229] , \labels[1][228] , 
	\labels[1][227] , \labels[1][226] , \labels[1][225] , 
	\labels[1][224] , \labels[1][223] , \labels[1][222] , 
	\labels[1][221] , \labels[1][220] , \labels[1][219] , 
	\labels[1][218] , \labels[1][217] , \labels[1][216] , 
	\labels[1][215] , \labels[1][214] , \labels[1][213] , 
	\labels[1][212] , \labels[1][211] , \labels[1][210] , 
	\labels[1][209] , \labels[1][208] , \labels[1][207] , 
	\labels[1][206] , \labels[1][205] , \labels[1][204] , 
	\labels[1][203] , \labels[1][202] , \labels[1][201] , 
	\labels[1][200] , \labels[1][199] , \labels[1][198] , 
	\labels[1][197] , \labels[1][196] , \labels[1][195] , 
	\labels[1][194] , \labels[1][193] , \labels[1][192] , 
	\labels[1][191] , \labels[1][190] , \labels[1][189] , 
	\labels[1][188] , \labels[1][187] , \labels[1][186] , 
	\labels[1][185] , \labels[1][184] , \labels[1][183] , 
	\labels[1][182] , \labels[1][181] , \labels[1][180] , 
	\labels[1][179] , \labels[1][178] , \labels[1][177] , 
	\labels[1][176] , \labels[1][175] , \labels[1][174] , 
	\labels[1][173] , \labels[1][172] , \labels[1][171] , 
	\labels[1][170] , \labels[1][169] , \labels[1][168] , 
	\labels[1][167] , \labels[1][166] , \labels[1][165] , 
	\labels[1][164] , \labels[1][163] , \labels[1][162] , 
	\labels[1][161] , \labels[1][160] , \labels[1][159] , 
	\labels[1][158] , \labels[1][157] , \labels[1][156] , 
	\labels[1][155] , \labels[1][154] , \labels[1][153] , 
	\labels[1][152] , \labels[1][151] , \labels[1][150] , 
	\labels[1][149] , \labels[1][148] , \labels[1][147] , 
	\labels[1][146] , \labels[1][145] , \labels[1][144] , 
	\labels[1][143] , \labels[1][142] , \labels[1][141] , 
	\labels[1][140] , \labels[1][139] , \labels[1][138] , 
	\labels[1][137] , \labels[1][136] , \labels[1][135] , 
	\labels[1][134] , \labels[1][133] , \labels[1][132] , 
	\labels[1][131] , \labels[1][130] , \labels[1][129] , 
	\labels[1][128] , \labels[1][127] , \labels[1][126] , 
	\labels[1][125] , \labels[1][124] , \labels[1][123] , 
	\labels[1][122] , \labels[1][121] , \labels[1][120] , 
	\labels[1][119] , \labels[1][118] , \labels[1][117] , 
	\labels[1][116] , \labels[1][115] , \labels[1][114] , 
	\labels[1][113] , \labels[1][112] , \labels[1][111] , 
	\labels[1][110] , \labels[1][109] , \labels[1][108] , 
	\labels[1][107] , \labels[1][106] , \labels[1][105] , 
	\labels[1][104] , \labels[1][103] , \labels[1][102] , 
	\labels[1][101] , \labels[1][100] , \labels[1][99] , \labels[1][98] , 
	\labels[1][97] , \labels[1][96] , \labels[1][95] , \labels[1][94] , 
	\labels[1][93] , \labels[1][92] , \labels[1][91] , \labels[1][90] , 
	\labels[1][89] , \labels[1][88] , \labels[1][87] , \labels[1][86] , 
	\labels[1][85] , \labels[1][84] , \labels[1][83] , \labels[1][82] , 
	\labels[1][81] , \labels[1][80] , \labels[1][79] , \labels[1][78] , 
	\labels[1][77] , \labels[1][76] , \labels[1][75] , \labels[1][74] , 
	\labels[1][73] , \labels[1][72] , \labels[1][71] , \labels[1][70] , 
	\labels[1][69] , \labels[1][68] , \labels[1][67] , \labels[1][66] , 
	\labels[1][65] , \labels[1][64] , \labels[1][63] , \labels[1][62] , 
	\labels[1][61] , \labels[1][60] , \labels[1][59] , \labels[1][58] , 
	\labels[1][57] , \labels[1][56] , \labels[1][55] , \labels[1][54] , 
	\labels[1][53] , \labels[1][52] , \labels[1][51] , \labels[1][50] , 
	\labels[1][49] , \labels[1][48] , \labels[1][47] , \labels[1][46] , 
	\labels[1][45] , \labels[1][44] , \labels[1][43] , \labels[1][42] , 
	\labels[1][41] , \labels[1][40] , \labels[1][39] , \labels[1][38] , 
	\labels[1][37] , \labels[1][36] , \labels[1][35] , \labels[1][34] , 
	\labels[1][33] , \labels[1][32] , \labels[1][31] , \labels[1][30] , 
	\labels[1][29] , \labels[1][28] , \labels[1][27] , \labels[1][26] , 
	\labels[1][25] , \labels[1][24] , \labels[1][23] , \labels[1][22] , 
	\labels[1][21] , \labels[1][20] , \labels[1][19] , \labels[1][18] , 
	\labels[1][17] , \labels[1][16] , \labels[1][15] , \labels[1][14] , 
	\labels[1][13] , \labels[1][12] , \labels[1][11] , \labels[1][10] , 
	\labels[1][9] , \labels[1][8] , \labels[1][7] , \labels[1][6] , 
	\labels[1][5] , \labels[1][4] , \labels[1][3] , \labels[1][2] , 
	\labels[1][1] , \labels[1][0] , \labels[0][271] , \labels[0][270] , 
	\labels[0][269] , \labels[0][268] , \labels[0][267] , 
	\labels[0][266] , \labels[0][265] , \labels[0][264] , 
	\labels[0][263] , \labels[0][262] , \labels[0][261] , 
	\labels[0][260] , \labels[0][259] , \labels[0][258] , 
	\labels[0][257] , \labels[0][256] , \labels[0][255] , 
	\labels[0][254] , \labels[0][253] , \labels[0][252] , 
	\labels[0][251] , \labels[0][250] , \labels[0][249] , 
	\labels[0][248] , \labels[0][247] , \labels[0][246] , 
	\labels[0][245] , \labels[0][244] , \labels[0][243] , 
	\labels[0][242] , \labels[0][241] , \labels[0][240] , 
	\labels[0][239] , \labels[0][238] , \labels[0][237] , 
	\labels[0][236] , \labels[0][235] , \labels[0][234] , 
	\labels[0][233] , \labels[0][232] , \labels[0][231] , 
	\labels[0][230] , \labels[0][229] , \labels[0][228] , 
	\labels[0][227] , \labels[0][226] , \labels[0][225] , 
	\labels[0][224] , \labels[0][223] , \labels[0][222] , 
	\labels[0][221] , \labels[0][220] , \labels[0][219] , 
	\labels[0][218] , \labels[0][217] , \labels[0][216] , 
	\labels[0][215] , \labels[0][214] , \labels[0][213] , 
	\labels[0][212] , \labels[0][211] , \labels[0][210] , 
	\labels[0][209] , \labels[0][208] , \labels[0][207] , 
	\labels[0][206] , \labels[0][205] , \labels[0][204] , 
	\labels[0][203] , \labels[0][202] , \labels[0][201] , 
	\labels[0][200] , \labels[0][199] , \labels[0][198] , 
	\labels[0][197] , \labels[0][196] , \labels[0][195] , 
	\labels[0][194] , \labels[0][193] , \labels[0][192] , 
	\labels[0][191] , \labels[0][190] , \labels[0][189] , 
	\labels[0][188] , \labels[0][187] , \labels[0][186] , 
	\labels[0][185] , \labels[0][184] , \labels[0][183] , 
	\labels[0][182] , \labels[0][181] , \labels[0][180] , 
	\labels[0][179] , \labels[0][178] , \labels[0][177] , 
	\labels[0][176] , \labels[0][175] , \labels[0][174] , 
	\labels[0][173] , \labels[0][172] , \labels[0][171] , 
	\labels[0][170] , \labels[0][169] , \labels[0][168] , 
	\labels[0][167] , \labels[0][166] , \labels[0][165] , 
	\labels[0][164] , \labels[0][163] , \labels[0][162] , 
	\labels[0][161] , \labels[0][160] , \labels[0][159] , 
	\labels[0][158] , \labels[0][157] , \labels[0][156] , 
	\labels[0][155] , \labels[0][154] , \labels[0][153] , 
	\labels[0][152] , \labels[0][151] , \labels[0][150] , 
	\labels[0][149] , \labels[0][148] , \labels[0][147] , 
	\labels[0][146] , \labels[0][145] , \labels[0][144] , 
	\labels[0][143] , \labels[0][142] , \labels[0][141] , 
	\labels[0][140] , \labels[0][139] , \labels[0][138] , 
	\labels[0][137] , \labels[0][136] , \labels[0][135] , 
	\labels[0][134] , \labels[0][133] , \labels[0][132] , 
	\labels[0][131] , \labels[0][130] , \labels[0][129] , 
	\labels[0][128] , \labels[0][127] , \labels[0][126] , 
	\labels[0][125] , \labels[0][124] , \labels[0][123] , 
	\labels[0][122] , \labels[0][121] , \labels[0][120] , 
	\labels[0][119] , \labels[0][118] , \labels[0][117] , 
	\labels[0][116] , \labels[0][115] , \labels[0][114] , 
	\labels[0][113] , \labels[0][112] , \labels[0][111] , 
	\labels[0][110] , \labels[0][109] , \labels[0][108] , 
	\labels[0][107] , \labels[0][106] , \labels[0][105] , 
	\labels[0][104] , \labels[0][103] , \labels[0][102] , 
	\labels[0][101] , \labels[0][100] , \labels[0][99] , \labels[0][98] , 
	\labels[0][97] , \labels[0][96] , \labels[0][95] , \labels[0][94] , 
	\labels[0][93] , \labels[0][92] , \labels[0][91] , \labels[0][90] , 
	\labels[0][89] , \labels[0][88] , \labels[0][87] , \labels[0][86] , 
	\labels[0][85] , \labels[0][84] , \labels[0][83] , \labels[0][82] , 
	\labels[0][81] , \labels[0][80] , \labels[0][79] , \labels[0][78] , 
	\labels[0][77] , \labels[0][76] , \labels[0][75] , \labels[0][74] , 
	\labels[0][73] , \labels[0][72] , \labels[0][71] , \labels[0][70] , 
	\labels[0][69] , \labels[0][68] , \labels[0][67] , \labels[0][66] , 
	\labels[0][65] , \labels[0][64] , \labels[0][63] , \labels[0][62] , 
	\labels[0][61] , \labels[0][60] , \labels[0][59] , \labels[0][58] , 
	\labels[0][57] , \labels[0][56] , \labels[0][55] , \labels[0][54] , 
	\labels[0][53] , \labels[0][52] , \labels[0][51] , \labels[0][50] , 
	\labels[0][49] , \labels[0][48] , \labels[0][47] , \labels[0][46] , 
	\labels[0][45] , \labels[0][44] , \labels[0][43] , \labels[0][42] , 
	\labels[0][41] , \labels[0][40] , \labels[0][39] , \labels[0][38] , 
	\labels[0][37] , \labels[0][36] , \labels[0][35] , \labels[0][34] , 
	\labels[0][33] , \labels[0][32] , \labels[0][31] , \labels[0][30] , 
	\labels[0][29] , \labels[0][28] , \labels[0][27] , \labels[0][26] , 
	\labels[0][25] , \labels[0][24] , \labels[0][23] , \labels[0][22] , 
	\labels[0][21] , \labels[0][20] , \labels[0][19] , \labels[0][18] , 
	\labels[0][17] , \labels[0][16] , \labels[0][15] , \labels[0][14] , 
	\labels[0][13] , \labels[0][12] , \labels[0][11] , \labels[0][10] , 
	\labels[0][9] , \labels[0][8] , \labels[0][7] , \labels[0][6] , 
	\labels[0][5] , \labels[0][4] , \labels[0][3] , \labels[0][2] , 
	\labels[0][1] , \labels[0][0] }, { \_zy_simnet_tvar_53[7][271] , 
	\_zy_simnet_tvar_53[7][270] , \_zy_simnet_tvar_53[7][269] , 
	\_zy_simnet_tvar_53[7][268] , \_zy_simnet_tvar_53[7][267] , 
	\_zy_simnet_tvar_53[7][266] , \_zy_simnet_tvar_53[7][265] , 
	\_zy_simnet_tvar_53[7][264] , \_zy_simnet_tvar_53[7][263] , 
	\_zy_simnet_tvar_53[7][262] , \_zy_simnet_tvar_53[7][261] , 
	\_zy_simnet_tvar_53[7][260] , \_zy_simnet_tvar_53[7][259] , 
	\_zy_simnet_tvar_53[7][258] , \_zy_simnet_tvar_53[7][257] , 
	\_zy_simnet_tvar_53[7][256] , \_zy_simnet_tvar_53[7][255] , 
	\_zy_simnet_tvar_53[7][254] , \_zy_simnet_tvar_53[7][253] , 
	\_zy_simnet_tvar_53[7][252] , \_zy_simnet_tvar_53[7][251] , 
	\_zy_simnet_tvar_53[7][250] , \_zy_simnet_tvar_53[7][249] , 
	\_zy_simnet_tvar_53[7][248] , \_zy_simnet_tvar_53[7][247] , 
	\_zy_simnet_tvar_53[7][246] , \_zy_simnet_tvar_53[7][245] , 
	\_zy_simnet_tvar_53[7][244] , \_zy_simnet_tvar_53[7][243] , 
	\_zy_simnet_tvar_53[7][242] , \_zy_simnet_tvar_53[7][241] , 
	\_zy_simnet_tvar_53[7][240] , \_zy_simnet_tvar_53[7][239] , 
	\_zy_simnet_tvar_53[7][238] , \_zy_simnet_tvar_53[7][237] , 
	\_zy_simnet_tvar_53[7][236] , \_zy_simnet_tvar_53[7][235] , 
	\_zy_simnet_tvar_53[7][234] , \_zy_simnet_tvar_53[7][233] , 
	\_zy_simnet_tvar_53[7][232] , \_zy_simnet_tvar_53[7][231] , 
	\_zy_simnet_tvar_53[7][230] , \_zy_simnet_tvar_53[7][229] , 
	\_zy_simnet_tvar_53[7][228] , \_zy_simnet_tvar_53[7][227] , 
	\_zy_simnet_tvar_53[7][226] , \_zy_simnet_tvar_53[7][225] , 
	\_zy_simnet_tvar_53[7][224] , \_zy_simnet_tvar_53[7][223] , 
	\_zy_simnet_tvar_53[7][222] , \_zy_simnet_tvar_53[7][221] , 
	\_zy_simnet_tvar_53[7][220] , \_zy_simnet_tvar_53[7][219] , 
	\_zy_simnet_tvar_53[7][218] , \_zy_simnet_tvar_53[7][217] , 
	\_zy_simnet_tvar_53[7][216] , \_zy_simnet_tvar_53[7][215] , 
	\_zy_simnet_tvar_53[7][214] , \_zy_simnet_tvar_53[7][213] , 
	\_zy_simnet_tvar_53[7][212] , \_zy_simnet_tvar_53[7][211] , 
	\_zy_simnet_tvar_53[7][210] , \_zy_simnet_tvar_53[7][209] , 
	\_zy_simnet_tvar_53[7][208] , \_zy_simnet_tvar_53[7][207] , 
	\_zy_simnet_tvar_53[7][206] , \_zy_simnet_tvar_53[7][205] , 
	\_zy_simnet_tvar_53[7][204] , \_zy_simnet_tvar_53[7][203] , 
	\_zy_simnet_tvar_53[7][202] , \_zy_simnet_tvar_53[7][201] , 
	\_zy_simnet_tvar_53[7][200] , \_zy_simnet_tvar_53[7][199] , 
	\_zy_simnet_tvar_53[7][198] , \_zy_simnet_tvar_53[7][197] , 
	\_zy_simnet_tvar_53[7][196] , \_zy_simnet_tvar_53[7][195] , 
	\_zy_simnet_tvar_53[7][194] , \_zy_simnet_tvar_53[7][193] , 
	\_zy_simnet_tvar_53[7][192] , \_zy_simnet_tvar_53[7][191] , 
	\_zy_simnet_tvar_53[7][190] , \_zy_simnet_tvar_53[7][189] , 
	\_zy_simnet_tvar_53[7][188] , \_zy_simnet_tvar_53[7][187] , 
	\_zy_simnet_tvar_53[7][186] , \_zy_simnet_tvar_53[7][185] , 
	\_zy_simnet_tvar_53[7][184] , \_zy_simnet_tvar_53[7][183] , 
	\_zy_simnet_tvar_53[7][182] , \_zy_simnet_tvar_53[7][181] , 
	\_zy_simnet_tvar_53[7][180] , \_zy_simnet_tvar_53[7][179] , 
	\_zy_simnet_tvar_53[7][178] , \_zy_simnet_tvar_53[7][177] , 
	\_zy_simnet_tvar_53[7][176] , \_zy_simnet_tvar_53[7][175] , 
	\_zy_simnet_tvar_53[7][174] , \_zy_simnet_tvar_53[7][173] , 
	\_zy_simnet_tvar_53[7][172] , \_zy_simnet_tvar_53[7][171] , 
	\_zy_simnet_tvar_53[7][170] , \_zy_simnet_tvar_53[7][169] , 
	\_zy_simnet_tvar_53[7][168] , \_zy_simnet_tvar_53[7][167] , 
	\_zy_simnet_tvar_53[7][166] , \_zy_simnet_tvar_53[7][165] , 
	\_zy_simnet_tvar_53[7][164] , \_zy_simnet_tvar_53[7][163] , 
	\_zy_simnet_tvar_53[7][162] , \_zy_simnet_tvar_53[7][161] , 
	\_zy_simnet_tvar_53[7][160] , \_zy_simnet_tvar_53[7][159] , 
	\_zy_simnet_tvar_53[7][158] , \_zy_simnet_tvar_53[7][157] , 
	\_zy_simnet_tvar_53[7][156] , \_zy_simnet_tvar_53[7][155] , 
	\_zy_simnet_tvar_53[7][154] , \_zy_simnet_tvar_53[7][153] , 
	\_zy_simnet_tvar_53[7][152] , \_zy_simnet_tvar_53[7][151] , 
	\_zy_simnet_tvar_53[7][150] , \_zy_simnet_tvar_53[7][149] , 
	\_zy_simnet_tvar_53[7][148] , \_zy_simnet_tvar_53[7][147] , 
	\_zy_simnet_tvar_53[7][146] , \_zy_simnet_tvar_53[7][145] , 
	\_zy_simnet_tvar_53[7][144] , \_zy_simnet_tvar_53[7][143] , 
	\_zy_simnet_tvar_53[7][142] , \_zy_simnet_tvar_53[7][141] , 
	\_zy_simnet_tvar_53[7][140] , \_zy_simnet_tvar_53[7][139] , 
	\_zy_simnet_tvar_53[7][138] , \_zy_simnet_tvar_53[7][137] , 
	\_zy_simnet_tvar_53[7][136] , \_zy_simnet_tvar_53[7][135] , 
	\_zy_simnet_tvar_53[7][134] , \_zy_simnet_tvar_53[7][133] , 
	\_zy_simnet_tvar_53[7][132] , \_zy_simnet_tvar_53[7][131] , 
	\_zy_simnet_tvar_53[7][130] , \_zy_simnet_tvar_53[7][129] , 
	\_zy_simnet_tvar_53[7][128] , \_zy_simnet_tvar_53[7][127] , 
	\_zy_simnet_tvar_53[7][126] , \_zy_simnet_tvar_53[7][125] , 
	\_zy_simnet_tvar_53[7][124] , \_zy_simnet_tvar_53[7][123] , 
	\_zy_simnet_tvar_53[7][122] , \_zy_simnet_tvar_53[7][121] , 
	\_zy_simnet_tvar_53[7][120] , \_zy_simnet_tvar_53[7][119] , 
	\_zy_simnet_tvar_53[7][118] , \_zy_simnet_tvar_53[7][117] , 
	\_zy_simnet_tvar_53[7][116] , \_zy_simnet_tvar_53[7][115] , 
	\_zy_simnet_tvar_53[7][114] , \_zy_simnet_tvar_53[7][113] , 
	\_zy_simnet_tvar_53[7][112] , \_zy_simnet_tvar_53[7][111] , 
	\_zy_simnet_tvar_53[7][110] , \_zy_simnet_tvar_53[7][109] , 
	\_zy_simnet_tvar_53[7][108] , \_zy_simnet_tvar_53[7][107] , 
	\_zy_simnet_tvar_53[7][106] , \_zy_simnet_tvar_53[7][105] , 
	\_zy_simnet_tvar_53[7][104] , \_zy_simnet_tvar_53[7][103] , 
	\_zy_simnet_tvar_53[7][102] , \_zy_simnet_tvar_53[7][101] , 
	\_zy_simnet_tvar_53[7][100] , \_zy_simnet_tvar_53[7][99] , 
	\_zy_simnet_tvar_53[7][98] , \_zy_simnet_tvar_53[7][97] , 
	\_zy_simnet_tvar_53[7][96] , \_zy_simnet_tvar_53[7][95] , 
	\_zy_simnet_tvar_53[7][94] , \_zy_simnet_tvar_53[7][93] , 
	\_zy_simnet_tvar_53[7][92] , \_zy_simnet_tvar_53[7][91] , 
	\_zy_simnet_tvar_53[7][90] , \_zy_simnet_tvar_53[7][89] , 
	\_zy_simnet_tvar_53[7][88] , \_zy_simnet_tvar_53[7][87] , 
	\_zy_simnet_tvar_53[7][86] , \_zy_simnet_tvar_53[7][85] , 
	\_zy_simnet_tvar_53[7][84] , \_zy_simnet_tvar_53[7][83] , 
	\_zy_simnet_tvar_53[7][82] , \_zy_simnet_tvar_53[7][81] , 
	\_zy_simnet_tvar_53[7][80] , \_zy_simnet_tvar_53[7][79] , 
	\_zy_simnet_tvar_53[7][78] , \_zy_simnet_tvar_53[7][77] , 
	\_zy_simnet_tvar_53[7][76] , \_zy_simnet_tvar_53[7][75] , 
	\_zy_simnet_tvar_53[7][74] , \_zy_simnet_tvar_53[7][73] , 
	\_zy_simnet_tvar_53[7][72] , \_zy_simnet_tvar_53[7][71] , 
	\_zy_simnet_tvar_53[7][70] , \_zy_simnet_tvar_53[7][69] , 
	\_zy_simnet_tvar_53[7][68] , \_zy_simnet_tvar_53[7][67] , 
	\_zy_simnet_tvar_53[7][66] , \_zy_simnet_tvar_53[7][65] , 
	\_zy_simnet_tvar_53[7][64] , \_zy_simnet_tvar_53[7][63] , 
	\_zy_simnet_tvar_53[7][62] , \_zy_simnet_tvar_53[7][61] , 
	\_zy_simnet_tvar_53[7][60] , \_zy_simnet_tvar_53[7][59] , 
	\_zy_simnet_tvar_53[7][58] , \_zy_simnet_tvar_53[7][57] , 
	\_zy_simnet_tvar_53[7][56] , \_zy_simnet_tvar_53[7][55] , 
	\_zy_simnet_tvar_53[7][54] , \_zy_simnet_tvar_53[7][53] , 
	\_zy_simnet_tvar_53[7][52] , \_zy_simnet_tvar_53[7][51] , 
	\_zy_simnet_tvar_53[7][50] , \_zy_simnet_tvar_53[7][49] , 
	\_zy_simnet_tvar_53[7][48] , \_zy_simnet_tvar_53[7][47] , 
	\_zy_simnet_tvar_53[7][46] , \_zy_simnet_tvar_53[7][45] , 
	\_zy_simnet_tvar_53[7][44] , \_zy_simnet_tvar_53[7][43] , 
	\_zy_simnet_tvar_53[7][42] , \_zy_simnet_tvar_53[7][41] , 
	\_zy_simnet_tvar_53[7][40] , \_zy_simnet_tvar_53[7][39] , 
	\_zy_simnet_tvar_53[7][38] , \_zy_simnet_tvar_53[7][37] , 
	\_zy_simnet_tvar_53[7][36] , \_zy_simnet_tvar_53[7][35] , 
	\_zy_simnet_tvar_53[7][34] , \_zy_simnet_tvar_53[7][33] , 
	\_zy_simnet_tvar_53[7][32] , \_zy_simnet_tvar_53[7][31] , 
	\_zy_simnet_tvar_53[7][30] , \_zy_simnet_tvar_53[7][29] , 
	\_zy_simnet_tvar_53[7][28] , \_zy_simnet_tvar_53[7][27] , 
	\_zy_simnet_tvar_53[7][26] , \_zy_simnet_tvar_53[7][25] , 
	\_zy_simnet_tvar_53[7][24] , \_zy_simnet_tvar_53[7][23] , 
	\_zy_simnet_tvar_53[7][22] , \_zy_simnet_tvar_53[7][21] , 
	\_zy_simnet_tvar_53[7][20] , \_zy_simnet_tvar_53[7][19] , 
	\_zy_simnet_tvar_53[7][18] , \_zy_simnet_tvar_53[7][17] , 
	\_zy_simnet_tvar_53[7][16] , \_zy_simnet_tvar_53[7][15] , 
	\_zy_simnet_tvar_53[7][14] , \_zy_simnet_tvar_53[7][13] , 
	\_zy_simnet_tvar_53[7][12] , \_zy_simnet_tvar_53[7][11] , 
	\_zy_simnet_tvar_53[7][10] , \_zy_simnet_tvar_53[7][9] , 
	\_zy_simnet_tvar_53[7][8] , \_zy_simnet_tvar_53[7][7] , 
	\_zy_simnet_tvar_53[7][6] , \_zy_simnet_tvar_53[7][5] , 
	\_zy_simnet_tvar_53[7][4] , \_zy_simnet_tvar_53[7][3] , 
	\_zy_simnet_tvar_53[7][2] , \_zy_simnet_tvar_53[7][1] , 
	\_zy_simnet_tvar_53[7][0] , \_zy_simnet_tvar_53[6][271] , 
	\_zy_simnet_tvar_53[6][270] , \_zy_simnet_tvar_53[6][269] , 
	\_zy_simnet_tvar_53[6][268] , \_zy_simnet_tvar_53[6][267] , 
	\_zy_simnet_tvar_53[6][266] , \_zy_simnet_tvar_53[6][265] , 
	\_zy_simnet_tvar_53[6][264] , \_zy_simnet_tvar_53[6][263] , 
	\_zy_simnet_tvar_53[6][262] , \_zy_simnet_tvar_53[6][261] , 
	\_zy_simnet_tvar_53[6][260] , \_zy_simnet_tvar_53[6][259] , 
	\_zy_simnet_tvar_53[6][258] , \_zy_simnet_tvar_53[6][257] , 
	\_zy_simnet_tvar_53[6][256] , \_zy_simnet_tvar_53[6][255] , 
	\_zy_simnet_tvar_53[6][254] , \_zy_simnet_tvar_53[6][253] , 
	\_zy_simnet_tvar_53[6][252] , \_zy_simnet_tvar_53[6][251] , 
	\_zy_simnet_tvar_53[6][250] , \_zy_simnet_tvar_53[6][249] , 
	\_zy_simnet_tvar_53[6][248] , \_zy_simnet_tvar_53[6][247] , 
	\_zy_simnet_tvar_53[6][246] , \_zy_simnet_tvar_53[6][245] , 
	\_zy_simnet_tvar_53[6][244] , \_zy_simnet_tvar_53[6][243] , 
	\_zy_simnet_tvar_53[6][242] , \_zy_simnet_tvar_53[6][241] , 
	\_zy_simnet_tvar_53[6][240] , \_zy_simnet_tvar_53[6][239] , 
	\_zy_simnet_tvar_53[6][238] , \_zy_simnet_tvar_53[6][237] , 
	\_zy_simnet_tvar_53[6][236] , \_zy_simnet_tvar_53[6][235] , 
	\_zy_simnet_tvar_53[6][234] , \_zy_simnet_tvar_53[6][233] , 
	\_zy_simnet_tvar_53[6][232] , \_zy_simnet_tvar_53[6][231] , 
	\_zy_simnet_tvar_53[6][230] , \_zy_simnet_tvar_53[6][229] , 
	\_zy_simnet_tvar_53[6][228] , \_zy_simnet_tvar_53[6][227] , 
	\_zy_simnet_tvar_53[6][226] , \_zy_simnet_tvar_53[6][225] , 
	\_zy_simnet_tvar_53[6][224] , \_zy_simnet_tvar_53[6][223] , 
	\_zy_simnet_tvar_53[6][222] , \_zy_simnet_tvar_53[6][221] , 
	\_zy_simnet_tvar_53[6][220] , \_zy_simnet_tvar_53[6][219] , 
	\_zy_simnet_tvar_53[6][218] , \_zy_simnet_tvar_53[6][217] , 
	\_zy_simnet_tvar_53[6][216] , \_zy_simnet_tvar_53[6][215] , 
	\_zy_simnet_tvar_53[6][214] , \_zy_simnet_tvar_53[6][213] , 
	\_zy_simnet_tvar_53[6][212] , \_zy_simnet_tvar_53[6][211] , 
	\_zy_simnet_tvar_53[6][210] , \_zy_simnet_tvar_53[6][209] , 
	\_zy_simnet_tvar_53[6][208] , \_zy_simnet_tvar_53[6][207] , 
	\_zy_simnet_tvar_53[6][206] , \_zy_simnet_tvar_53[6][205] , 
	\_zy_simnet_tvar_53[6][204] , \_zy_simnet_tvar_53[6][203] , 
	\_zy_simnet_tvar_53[6][202] , \_zy_simnet_tvar_53[6][201] , 
	\_zy_simnet_tvar_53[6][200] , \_zy_simnet_tvar_53[6][199] , 
	\_zy_simnet_tvar_53[6][198] , \_zy_simnet_tvar_53[6][197] , 
	\_zy_simnet_tvar_53[6][196] , \_zy_simnet_tvar_53[6][195] , 
	\_zy_simnet_tvar_53[6][194] , \_zy_simnet_tvar_53[6][193] , 
	\_zy_simnet_tvar_53[6][192] , \_zy_simnet_tvar_53[6][191] , 
	\_zy_simnet_tvar_53[6][190] , \_zy_simnet_tvar_53[6][189] , 
	\_zy_simnet_tvar_53[6][188] , \_zy_simnet_tvar_53[6][187] , 
	\_zy_simnet_tvar_53[6][186] , \_zy_simnet_tvar_53[6][185] , 
	\_zy_simnet_tvar_53[6][184] , \_zy_simnet_tvar_53[6][183] , 
	\_zy_simnet_tvar_53[6][182] , \_zy_simnet_tvar_53[6][181] , 
	\_zy_simnet_tvar_53[6][180] , \_zy_simnet_tvar_53[6][179] , 
	\_zy_simnet_tvar_53[6][178] , \_zy_simnet_tvar_53[6][177] , 
	\_zy_simnet_tvar_53[6][176] , \_zy_simnet_tvar_53[6][175] , 
	\_zy_simnet_tvar_53[6][174] , \_zy_simnet_tvar_53[6][173] , 
	\_zy_simnet_tvar_53[6][172] , \_zy_simnet_tvar_53[6][171] , 
	\_zy_simnet_tvar_53[6][170] , \_zy_simnet_tvar_53[6][169] , 
	\_zy_simnet_tvar_53[6][168] , \_zy_simnet_tvar_53[6][167] , 
	\_zy_simnet_tvar_53[6][166] , \_zy_simnet_tvar_53[6][165] , 
	\_zy_simnet_tvar_53[6][164] , \_zy_simnet_tvar_53[6][163] , 
	\_zy_simnet_tvar_53[6][162] , \_zy_simnet_tvar_53[6][161] , 
	\_zy_simnet_tvar_53[6][160] , \_zy_simnet_tvar_53[6][159] , 
	\_zy_simnet_tvar_53[6][158] , \_zy_simnet_tvar_53[6][157] , 
	\_zy_simnet_tvar_53[6][156] , \_zy_simnet_tvar_53[6][155] , 
	\_zy_simnet_tvar_53[6][154] , \_zy_simnet_tvar_53[6][153] , 
	\_zy_simnet_tvar_53[6][152] , \_zy_simnet_tvar_53[6][151] , 
	\_zy_simnet_tvar_53[6][150] , \_zy_simnet_tvar_53[6][149] , 
	\_zy_simnet_tvar_53[6][148] , \_zy_simnet_tvar_53[6][147] , 
	\_zy_simnet_tvar_53[6][146] , \_zy_simnet_tvar_53[6][145] , 
	\_zy_simnet_tvar_53[6][144] , \_zy_simnet_tvar_53[6][143] , 
	\_zy_simnet_tvar_53[6][142] , \_zy_simnet_tvar_53[6][141] , 
	\_zy_simnet_tvar_53[6][140] , \_zy_simnet_tvar_53[6][139] , 
	\_zy_simnet_tvar_53[6][138] , \_zy_simnet_tvar_53[6][137] , 
	\_zy_simnet_tvar_53[6][136] , \_zy_simnet_tvar_53[6][135] , 
	\_zy_simnet_tvar_53[6][134] , \_zy_simnet_tvar_53[6][133] , 
	\_zy_simnet_tvar_53[6][132] , \_zy_simnet_tvar_53[6][131] , 
	\_zy_simnet_tvar_53[6][130] , \_zy_simnet_tvar_53[6][129] , 
	\_zy_simnet_tvar_53[6][128] , \_zy_simnet_tvar_53[6][127] , 
	\_zy_simnet_tvar_53[6][126] , \_zy_simnet_tvar_53[6][125] , 
	\_zy_simnet_tvar_53[6][124] , \_zy_simnet_tvar_53[6][123] , 
	\_zy_simnet_tvar_53[6][122] , \_zy_simnet_tvar_53[6][121] , 
	\_zy_simnet_tvar_53[6][120] , \_zy_simnet_tvar_53[6][119] , 
	\_zy_simnet_tvar_53[6][118] , \_zy_simnet_tvar_53[6][117] , 
	\_zy_simnet_tvar_53[6][116] , \_zy_simnet_tvar_53[6][115] , 
	\_zy_simnet_tvar_53[6][114] , \_zy_simnet_tvar_53[6][113] , 
	\_zy_simnet_tvar_53[6][112] , \_zy_simnet_tvar_53[6][111] , 
	\_zy_simnet_tvar_53[6][110] , \_zy_simnet_tvar_53[6][109] , 
	\_zy_simnet_tvar_53[6][108] , \_zy_simnet_tvar_53[6][107] , 
	\_zy_simnet_tvar_53[6][106] , \_zy_simnet_tvar_53[6][105] , 
	\_zy_simnet_tvar_53[6][104] , \_zy_simnet_tvar_53[6][103] , 
	\_zy_simnet_tvar_53[6][102] , \_zy_simnet_tvar_53[6][101] , 
	\_zy_simnet_tvar_53[6][100] , \_zy_simnet_tvar_53[6][99] , 
	\_zy_simnet_tvar_53[6][98] , \_zy_simnet_tvar_53[6][97] , 
	\_zy_simnet_tvar_53[6][96] , \_zy_simnet_tvar_53[6][95] , 
	\_zy_simnet_tvar_53[6][94] , \_zy_simnet_tvar_53[6][93] , 
	\_zy_simnet_tvar_53[6][92] , \_zy_simnet_tvar_53[6][91] , 
	\_zy_simnet_tvar_53[6][90] , \_zy_simnet_tvar_53[6][89] , 
	\_zy_simnet_tvar_53[6][88] , \_zy_simnet_tvar_53[6][87] , 
	\_zy_simnet_tvar_53[6][86] , \_zy_simnet_tvar_53[6][85] , 
	\_zy_simnet_tvar_53[6][84] , \_zy_simnet_tvar_53[6][83] , 
	\_zy_simnet_tvar_53[6][82] , \_zy_simnet_tvar_53[6][81] , 
	\_zy_simnet_tvar_53[6][80] , \_zy_simnet_tvar_53[6][79] , 
	\_zy_simnet_tvar_53[6][78] , \_zy_simnet_tvar_53[6][77] , 
	\_zy_simnet_tvar_53[6][76] , \_zy_simnet_tvar_53[6][75] , 
	\_zy_simnet_tvar_53[6][74] , \_zy_simnet_tvar_53[6][73] , 
	\_zy_simnet_tvar_53[6][72] , \_zy_simnet_tvar_53[6][71] , 
	\_zy_simnet_tvar_53[6][70] , \_zy_simnet_tvar_53[6][69] , 
	\_zy_simnet_tvar_53[6][68] , \_zy_simnet_tvar_53[6][67] , 
	\_zy_simnet_tvar_53[6][66] , \_zy_simnet_tvar_53[6][65] , 
	\_zy_simnet_tvar_53[6][64] , \_zy_simnet_tvar_53[6][63] , 
	\_zy_simnet_tvar_53[6][62] , \_zy_simnet_tvar_53[6][61] , 
	\_zy_simnet_tvar_53[6][60] , \_zy_simnet_tvar_53[6][59] , 
	\_zy_simnet_tvar_53[6][58] , \_zy_simnet_tvar_53[6][57] , 
	\_zy_simnet_tvar_53[6][56] , \_zy_simnet_tvar_53[6][55] , 
	\_zy_simnet_tvar_53[6][54] , \_zy_simnet_tvar_53[6][53] , 
	\_zy_simnet_tvar_53[6][52] , \_zy_simnet_tvar_53[6][51] , 
	\_zy_simnet_tvar_53[6][50] , \_zy_simnet_tvar_53[6][49] , 
	\_zy_simnet_tvar_53[6][48] , \_zy_simnet_tvar_53[6][47] , 
	\_zy_simnet_tvar_53[6][46] , \_zy_simnet_tvar_53[6][45] , 
	\_zy_simnet_tvar_53[6][44] , \_zy_simnet_tvar_53[6][43] , 
	\_zy_simnet_tvar_53[6][42] , \_zy_simnet_tvar_53[6][41] , 
	\_zy_simnet_tvar_53[6][40] , \_zy_simnet_tvar_53[6][39] , 
	\_zy_simnet_tvar_53[6][38] , \_zy_simnet_tvar_53[6][37] , 
	\_zy_simnet_tvar_53[6][36] , \_zy_simnet_tvar_53[6][35] , 
	\_zy_simnet_tvar_53[6][34] , \_zy_simnet_tvar_53[6][33] , 
	\_zy_simnet_tvar_53[6][32] , \_zy_simnet_tvar_53[6][31] , 
	\_zy_simnet_tvar_53[6][30] , \_zy_simnet_tvar_53[6][29] , 
	\_zy_simnet_tvar_53[6][28] , \_zy_simnet_tvar_53[6][27] , 
	\_zy_simnet_tvar_53[6][26] , \_zy_simnet_tvar_53[6][25] , 
	\_zy_simnet_tvar_53[6][24] , \_zy_simnet_tvar_53[6][23] , 
	\_zy_simnet_tvar_53[6][22] , \_zy_simnet_tvar_53[6][21] , 
	\_zy_simnet_tvar_53[6][20] , \_zy_simnet_tvar_53[6][19] , 
	\_zy_simnet_tvar_53[6][18] , \_zy_simnet_tvar_53[6][17] , 
	\_zy_simnet_tvar_53[6][16] , \_zy_simnet_tvar_53[6][15] , 
	\_zy_simnet_tvar_53[6][14] , \_zy_simnet_tvar_53[6][13] , 
	\_zy_simnet_tvar_53[6][12] , \_zy_simnet_tvar_53[6][11] , 
	\_zy_simnet_tvar_53[6][10] , \_zy_simnet_tvar_53[6][9] , 
	\_zy_simnet_tvar_53[6][8] , \_zy_simnet_tvar_53[6][7] , 
	\_zy_simnet_tvar_53[6][6] , \_zy_simnet_tvar_53[6][5] , 
	\_zy_simnet_tvar_53[6][4] , \_zy_simnet_tvar_53[6][3] , 
	\_zy_simnet_tvar_53[6][2] , \_zy_simnet_tvar_53[6][1] , 
	\_zy_simnet_tvar_53[6][0] , \_zy_simnet_tvar_53[5][271] , 
	\_zy_simnet_tvar_53[5][270] , \_zy_simnet_tvar_53[5][269] , 
	\_zy_simnet_tvar_53[5][268] , \_zy_simnet_tvar_53[5][267] , 
	\_zy_simnet_tvar_53[5][266] , \_zy_simnet_tvar_53[5][265] , 
	\_zy_simnet_tvar_53[5][264] , \_zy_simnet_tvar_53[5][263] , 
	\_zy_simnet_tvar_53[5][262] , \_zy_simnet_tvar_53[5][261] , 
	\_zy_simnet_tvar_53[5][260] , \_zy_simnet_tvar_53[5][259] , 
	\_zy_simnet_tvar_53[5][258] , \_zy_simnet_tvar_53[5][257] , 
	\_zy_simnet_tvar_53[5][256] , \_zy_simnet_tvar_53[5][255] , 
	\_zy_simnet_tvar_53[5][254] , \_zy_simnet_tvar_53[5][253] , 
	\_zy_simnet_tvar_53[5][252] , \_zy_simnet_tvar_53[5][251] , 
	\_zy_simnet_tvar_53[5][250] , \_zy_simnet_tvar_53[5][249] , 
	\_zy_simnet_tvar_53[5][248] , \_zy_simnet_tvar_53[5][247] , 
	\_zy_simnet_tvar_53[5][246] , \_zy_simnet_tvar_53[5][245] , 
	\_zy_simnet_tvar_53[5][244] , \_zy_simnet_tvar_53[5][243] , 
	\_zy_simnet_tvar_53[5][242] , \_zy_simnet_tvar_53[5][241] , 
	\_zy_simnet_tvar_53[5][240] , \_zy_simnet_tvar_53[5][239] , 
	\_zy_simnet_tvar_53[5][238] , \_zy_simnet_tvar_53[5][237] , 
	\_zy_simnet_tvar_53[5][236] , \_zy_simnet_tvar_53[5][235] , 
	\_zy_simnet_tvar_53[5][234] , \_zy_simnet_tvar_53[5][233] , 
	\_zy_simnet_tvar_53[5][232] , \_zy_simnet_tvar_53[5][231] , 
	\_zy_simnet_tvar_53[5][230] , \_zy_simnet_tvar_53[5][229] , 
	\_zy_simnet_tvar_53[5][228] , \_zy_simnet_tvar_53[5][227] , 
	\_zy_simnet_tvar_53[5][226] , \_zy_simnet_tvar_53[5][225] , 
	\_zy_simnet_tvar_53[5][224] , \_zy_simnet_tvar_53[5][223] , 
	\_zy_simnet_tvar_53[5][222] , \_zy_simnet_tvar_53[5][221] , 
	\_zy_simnet_tvar_53[5][220] , \_zy_simnet_tvar_53[5][219] , 
	\_zy_simnet_tvar_53[5][218] , \_zy_simnet_tvar_53[5][217] , 
	\_zy_simnet_tvar_53[5][216] , \_zy_simnet_tvar_53[5][215] , 
	\_zy_simnet_tvar_53[5][214] , \_zy_simnet_tvar_53[5][213] , 
	\_zy_simnet_tvar_53[5][212] , \_zy_simnet_tvar_53[5][211] , 
	\_zy_simnet_tvar_53[5][210] , \_zy_simnet_tvar_53[5][209] , 
	\_zy_simnet_tvar_53[5][208] , \_zy_simnet_tvar_53[5][207] , 
	\_zy_simnet_tvar_53[5][206] , \_zy_simnet_tvar_53[5][205] , 
	\_zy_simnet_tvar_53[5][204] , \_zy_simnet_tvar_53[5][203] , 
	\_zy_simnet_tvar_53[5][202] , \_zy_simnet_tvar_53[5][201] , 
	\_zy_simnet_tvar_53[5][200] , \_zy_simnet_tvar_53[5][199] , 
	\_zy_simnet_tvar_53[5][198] , \_zy_simnet_tvar_53[5][197] , 
	\_zy_simnet_tvar_53[5][196] , \_zy_simnet_tvar_53[5][195] , 
	\_zy_simnet_tvar_53[5][194] , \_zy_simnet_tvar_53[5][193] , 
	\_zy_simnet_tvar_53[5][192] , \_zy_simnet_tvar_53[5][191] , 
	\_zy_simnet_tvar_53[5][190] , \_zy_simnet_tvar_53[5][189] , 
	\_zy_simnet_tvar_53[5][188] , \_zy_simnet_tvar_53[5][187] , 
	\_zy_simnet_tvar_53[5][186] , \_zy_simnet_tvar_53[5][185] , 
	\_zy_simnet_tvar_53[5][184] , \_zy_simnet_tvar_53[5][183] , 
	\_zy_simnet_tvar_53[5][182] , \_zy_simnet_tvar_53[5][181] , 
	\_zy_simnet_tvar_53[5][180] , \_zy_simnet_tvar_53[5][179] , 
	\_zy_simnet_tvar_53[5][178] , \_zy_simnet_tvar_53[5][177] , 
	\_zy_simnet_tvar_53[5][176] , \_zy_simnet_tvar_53[5][175] , 
	\_zy_simnet_tvar_53[5][174] , \_zy_simnet_tvar_53[5][173] , 
	\_zy_simnet_tvar_53[5][172] , \_zy_simnet_tvar_53[5][171] , 
	\_zy_simnet_tvar_53[5][170] , \_zy_simnet_tvar_53[5][169] , 
	\_zy_simnet_tvar_53[5][168] , \_zy_simnet_tvar_53[5][167] , 
	\_zy_simnet_tvar_53[5][166] , \_zy_simnet_tvar_53[5][165] , 
	\_zy_simnet_tvar_53[5][164] , \_zy_simnet_tvar_53[5][163] , 
	\_zy_simnet_tvar_53[5][162] , \_zy_simnet_tvar_53[5][161] , 
	\_zy_simnet_tvar_53[5][160] , \_zy_simnet_tvar_53[5][159] , 
	\_zy_simnet_tvar_53[5][158] , \_zy_simnet_tvar_53[5][157] , 
	\_zy_simnet_tvar_53[5][156] , \_zy_simnet_tvar_53[5][155] , 
	\_zy_simnet_tvar_53[5][154] , \_zy_simnet_tvar_53[5][153] , 
	\_zy_simnet_tvar_53[5][152] , \_zy_simnet_tvar_53[5][151] , 
	\_zy_simnet_tvar_53[5][150] , \_zy_simnet_tvar_53[5][149] , 
	\_zy_simnet_tvar_53[5][148] , \_zy_simnet_tvar_53[5][147] , 
	\_zy_simnet_tvar_53[5][146] , \_zy_simnet_tvar_53[5][145] , 
	\_zy_simnet_tvar_53[5][144] , \_zy_simnet_tvar_53[5][143] , 
	\_zy_simnet_tvar_53[5][142] , \_zy_simnet_tvar_53[5][141] , 
	\_zy_simnet_tvar_53[5][140] , \_zy_simnet_tvar_53[5][139] , 
	\_zy_simnet_tvar_53[5][138] , \_zy_simnet_tvar_53[5][137] , 
	\_zy_simnet_tvar_53[5][136] , \_zy_simnet_tvar_53[5][135] , 
	\_zy_simnet_tvar_53[5][134] , \_zy_simnet_tvar_53[5][133] , 
	\_zy_simnet_tvar_53[5][132] , \_zy_simnet_tvar_53[5][131] , 
	\_zy_simnet_tvar_53[5][130] , \_zy_simnet_tvar_53[5][129] , 
	\_zy_simnet_tvar_53[5][128] , \_zy_simnet_tvar_53[5][127] , 
	\_zy_simnet_tvar_53[5][126] , \_zy_simnet_tvar_53[5][125] , 
	\_zy_simnet_tvar_53[5][124] , \_zy_simnet_tvar_53[5][123] , 
	\_zy_simnet_tvar_53[5][122] , \_zy_simnet_tvar_53[5][121] , 
	\_zy_simnet_tvar_53[5][120] , \_zy_simnet_tvar_53[5][119] , 
	\_zy_simnet_tvar_53[5][118] , \_zy_simnet_tvar_53[5][117] , 
	\_zy_simnet_tvar_53[5][116] , \_zy_simnet_tvar_53[5][115] , 
	\_zy_simnet_tvar_53[5][114] , \_zy_simnet_tvar_53[5][113] , 
	\_zy_simnet_tvar_53[5][112] , \_zy_simnet_tvar_53[5][111] , 
	\_zy_simnet_tvar_53[5][110] , \_zy_simnet_tvar_53[5][109] , 
	\_zy_simnet_tvar_53[5][108] , \_zy_simnet_tvar_53[5][107] , 
	\_zy_simnet_tvar_53[5][106] , \_zy_simnet_tvar_53[5][105] , 
	\_zy_simnet_tvar_53[5][104] , \_zy_simnet_tvar_53[5][103] , 
	\_zy_simnet_tvar_53[5][102] , \_zy_simnet_tvar_53[5][101] , 
	\_zy_simnet_tvar_53[5][100] , \_zy_simnet_tvar_53[5][99] , 
	\_zy_simnet_tvar_53[5][98] , \_zy_simnet_tvar_53[5][97] , 
	\_zy_simnet_tvar_53[5][96] , \_zy_simnet_tvar_53[5][95] , 
	\_zy_simnet_tvar_53[5][94] , \_zy_simnet_tvar_53[5][93] , 
	\_zy_simnet_tvar_53[5][92] , \_zy_simnet_tvar_53[5][91] , 
	\_zy_simnet_tvar_53[5][90] , \_zy_simnet_tvar_53[5][89] , 
	\_zy_simnet_tvar_53[5][88] , \_zy_simnet_tvar_53[5][87] , 
	\_zy_simnet_tvar_53[5][86] , \_zy_simnet_tvar_53[5][85] , 
	\_zy_simnet_tvar_53[5][84] , \_zy_simnet_tvar_53[5][83] , 
	\_zy_simnet_tvar_53[5][82] , \_zy_simnet_tvar_53[5][81] , 
	\_zy_simnet_tvar_53[5][80] , \_zy_simnet_tvar_53[5][79] , 
	\_zy_simnet_tvar_53[5][78] , \_zy_simnet_tvar_53[5][77] , 
	\_zy_simnet_tvar_53[5][76] , \_zy_simnet_tvar_53[5][75] , 
	\_zy_simnet_tvar_53[5][74] , \_zy_simnet_tvar_53[5][73] , 
	\_zy_simnet_tvar_53[5][72] , \_zy_simnet_tvar_53[5][71] , 
	\_zy_simnet_tvar_53[5][70] , \_zy_simnet_tvar_53[5][69] , 
	\_zy_simnet_tvar_53[5][68] , \_zy_simnet_tvar_53[5][67] , 
	\_zy_simnet_tvar_53[5][66] , \_zy_simnet_tvar_53[5][65] , 
	\_zy_simnet_tvar_53[5][64] , \_zy_simnet_tvar_53[5][63] , 
	\_zy_simnet_tvar_53[5][62] , \_zy_simnet_tvar_53[5][61] , 
	\_zy_simnet_tvar_53[5][60] , \_zy_simnet_tvar_53[5][59] , 
	\_zy_simnet_tvar_53[5][58] , \_zy_simnet_tvar_53[5][57] , 
	\_zy_simnet_tvar_53[5][56] , \_zy_simnet_tvar_53[5][55] , 
	\_zy_simnet_tvar_53[5][54] , \_zy_simnet_tvar_53[5][53] , 
	\_zy_simnet_tvar_53[5][52] , \_zy_simnet_tvar_53[5][51] , 
	\_zy_simnet_tvar_53[5][50] , \_zy_simnet_tvar_53[5][49] , 
	\_zy_simnet_tvar_53[5][48] , \_zy_simnet_tvar_53[5][47] , 
	\_zy_simnet_tvar_53[5][46] , \_zy_simnet_tvar_53[5][45] , 
	\_zy_simnet_tvar_53[5][44] , \_zy_simnet_tvar_53[5][43] , 
	\_zy_simnet_tvar_53[5][42] , \_zy_simnet_tvar_53[5][41] , 
	\_zy_simnet_tvar_53[5][40] , \_zy_simnet_tvar_53[5][39] , 
	\_zy_simnet_tvar_53[5][38] , \_zy_simnet_tvar_53[5][37] , 
	\_zy_simnet_tvar_53[5][36] , \_zy_simnet_tvar_53[5][35] , 
	\_zy_simnet_tvar_53[5][34] , \_zy_simnet_tvar_53[5][33] , 
	\_zy_simnet_tvar_53[5][32] , \_zy_simnet_tvar_53[5][31] , 
	\_zy_simnet_tvar_53[5][30] , \_zy_simnet_tvar_53[5][29] , 
	\_zy_simnet_tvar_53[5][28] , \_zy_simnet_tvar_53[5][27] , 
	\_zy_simnet_tvar_53[5][26] , \_zy_simnet_tvar_53[5][25] , 
	\_zy_simnet_tvar_53[5][24] , \_zy_simnet_tvar_53[5][23] , 
	\_zy_simnet_tvar_53[5][22] , \_zy_simnet_tvar_53[5][21] , 
	\_zy_simnet_tvar_53[5][20] , \_zy_simnet_tvar_53[5][19] , 
	\_zy_simnet_tvar_53[5][18] , \_zy_simnet_tvar_53[5][17] , 
	\_zy_simnet_tvar_53[5][16] , \_zy_simnet_tvar_53[5][15] , 
	\_zy_simnet_tvar_53[5][14] , \_zy_simnet_tvar_53[5][13] , 
	\_zy_simnet_tvar_53[5][12] , \_zy_simnet_tvar_53[5][11] , 
	\_zy_simnet_tvar_53[5][10] , \_zy_simnet_tvar_53[5][9] , 
	\_zy_simnet_tvar_53[5][8] , \_zy_simnet_tvar_53[5][7] , 
	\_zy_simnet_tvar_53[5][6] , \_zy_simnet_tvar_53[5][5] , 
	\_zy_simnet_tvar_53[5][4] , \_zy_simnet_tvar_53[5][3] , 
	\_zy_simnet_tvar_53[5][2] , \_zy_simnet_tvar_53[5][1] , 
	\_zy_simnet_tvar_53[5][0] , \_zy_simnet_tvar_53[4][271] , 
	\_zy_simnet_tvar_53[4][270] , \_zy_simnet_tvar_53[4][269] , 
	\_zy_simnet_tvar_53[4][268] , \_zy_simnet_tvar_53[4][267] , 
	\_zy_simnet_tvar_53[4][266] , \_zy_simnet_tvar_53[4][265] , 
	\_zy_simnet_tvar_53[4][264] , \_zy_simnet_tvar_53[4][263] , 
	\_zy_simnet_tvar_53[4][262] , \_zy_simnet_tvar_53[4][261] , 
	\_zy_simnet_tvar_53[4][260] , \_zy_simnet_tvar_53[4][259] , 
	\_zy_simnet_tvar_53[4][258] , \_zy_simnet_tvar_53[4][257] , 
	\_zy_simnet_tvar_53[4][256] , \_zy_simnet_tvar_53[4][255] , 
	\_zy_simnet_tvar_53[4][254] , \_zy_simnet_tvar_53[4][253] , 
	\_zy_simnet_tvar_53[4][252] , \_zy_simnet_tvar_53[4][251] , 
	\_zy_simnet_tvar_53[4][250] , \_zy_simnet_tvar_53[4][249] , 
	\_zy_simnet_tvar_53[4][248] , \_zy_simnet_tvar_53[4][247] , 
	\_zy_simnet_tvar_53[4][246] , \_zy_simnet_tvar_53[4][245] , 
	\_zy_simnet_tvar_53[4][244] , \_zy_simnet_tvar_53[4][243] , 
	\_zy_simnet_tvar_53[4][242] , \_zy_simnet_tvar_53[4][241] , 
	\_zy_simnet_tvar_53[4][240] , \_zy_simnet_tvar_53[4][239] , 
	\_zy_simnet_tvar_53[4][238] , \_zy_simnet_tvar_53[4][237] , 
	\_zy_simnet_tvar_53[4][236] , \_zy_simnet_tvar_53[4][235] , 
	\_zy_simnet_tvar_53[4][234] , \_zy_simnet_tvar_53[4][233] , 
	\_zy_simnet_tvar_53[4][232] , \_zy_simnet_tvar_53[4][231] , 
	\_zy_simnet_tvar_53[4][230] , \_zy_simnet_tvar_53[4][229] , 
	\_zy_simnet_tvar_53[4][228] , \_zy_simnet_tvar_53[4][227] , 
	\_zy_simnet_tvar_53[4][226] , \_zy_simnet_tvar_53[4][225] , 
	\_zy_simnet_tvar_53[4][224] , \_zy_simnet_tvar_53[4][223] , 
	\_zy_simnet_tvar_53[4][222] , \_zy_simnet_tvar_53[4][221] , 
	\_zy_simnet_tvar_53[4][220] , \_zy_simnet_tvar_53[4][219] , 
	\_zy_simnet_tvar_53[4][218] , \_zy_simnet_tvar_53[4][217] , 
	\_zy_simnet_tvar_53[4][216] , \_zy_simnet_tvar_53[4][215] , 
	\_zy_simnet_tvar_53[4][214] , \_zy_simnet_tvar_53[4][213] , 
	\_zy_simnet_tvar_53[4][212] , \_zy_simnet_tvar_53[4][211] , 
	\_zy_simnet_tvar_53[4][210] , \_zy_simnet_tvar_53[4][209] , 
	\_zy_simnet_tvar_53[4][208] , \_zy_simnet_tvar_53[4][207] , 
	\_zy_simnet_tvar_53[4][206] , \_zy_simnet_tvar_53[4][205] , 
	\_zy_simnet_tvar_53[4][204] , \_zy_simnet_tvar_53[4][203] , 
	\_zy_simnet_tvar_53[4][202] , \_zy_simnet_tvar_53[4][201] , 
	\_zy_simnet_tvar_53[4][200] , \_zy_simnet_tvar_53[4][199] , 
	\_zy_simnet_tvar_53[4][198] , \_zy_simnet_tvar_53[4][197] , 
	\_zy_simnet_tvar_53[4][196] , \_zy_simnet_tvar_53[4][195] , 
	\_zy_simnet_tvar_53[4][194] , \_zy_simnet_tvar_53[4][193] , 
	\_zy_simnet_tvar_53[4][192] , \_zy_simnet_tvar_53[4][191] , 
	\_zy_simnet_tvar_53[4][190] , \_zy_simnet_tvar_53[4][189] , 
	\_zy_simnet_tvar_53[4][188] , \_zy_simnet_tvar_53[4][187] , 
	\_zy_simnet_tvar_53[4][186] , \_zy_simnet_tvar_53[4][185] , 
	\_zy_simnet_tvar_53[4][184] , \_zy_simnet_tvar_53[4][183] , 
	\_zy_simnet_tvar_53[4][182] , \_zy_simnet_tvar_53[4][181] , 
	\_zy_simnet_tvar_53[4][180] , \_zy_simnet_tvar_53[4][179] , 
	\_zy_simnet_tvar_53[4][178] , \_zy_simnet_tvar_53[4][177] , 
	\_zy_simnet_tvar_53[4][176] , \_zy_simnet_tvar_53[4][175] , 
	\_zy_simnet_tvar_53[4][174] , \_zy_simnet_tvar_53[4][173] , 
	\_zy_simnet_tvar_53[4][172] , \_zy_simnet_tvar_53[4][171] , 
	\_zy_simnet_tvar_53[4][170] , \_zy_simnet_tvar_53[4][169] , 
	\_zy_simnet_tvar_53[4][168] , \_zy_simnet_tvar_53[4][167] , 
	\_zy_simnet_tvar_53[4][166] , \_zy_simnet_tvar_53[4][165] , 
	\_zy_simnet_tvar_53[4][164] , \_zy_simnet_tvar_53[4][163] , 
	\_zy_simnet_tvar_53[4][162] , \_zy_simnet_tvar_53[4][161] , 
	\_zy_simnet_tvar_53[4][160] , \_zy_simnet_tvar_53[4][159] , 
	\_zy_simnet_tvar_53[4][158] , \_zy_simnet_tvar_53[4][157] , 
	\_zy_simnet_tvar_53[4][156] , \_zy_simnet_tvar_53[4][155] , 
	\_zy_simnet_tvar_53[4][154] , \_zy_simnet_tvar_53[4][153] , 
	\_zy_simnet_tvar_53[4][152] , \_zy_simnet_tvar_53[4][151] , 
	\_zy_simnet_tvar_53[4][150] , \_zy_simnet_tvar_53[4][149] , 
	\_zy_simnet_tvar_53[4][148] , \_zy_simnet_tvar_53[4][147] , 
	\_zy_simnet_tvar_53[4][146] , \_zy_simnet_tvar_53[4][145] , 
	\_zy_simnet_tvar_53[4][144] , \_zy_simnet_tvar_53[4][143] , 
	\_zy_simnet_tvar_53[4][142] , \_zy_simnet_tvar_53[4][141] , 
	\_zy_simnet_tvar_53[4][140] , \_zy_simnet_tvar_53[4][139] , 
	\_zy_simnet_tvar_53[4][138] , \_zy_simnet_tvar_53[4][137] , 
	\_zy_simnet_tvar_53[4][136] , \_zy_simnet_tvar_53[4][135] , 
	\_zy_simnet_tvar_53[4][134] , \_zy_simnet_tvar_53[4][133] , 
	\_zy_simnet_tvar_53[4][132] , \_zy_simnet_tvar_53[4][131] , 
	\_zy_simnet_tvar_53[4][130] , \_zy_simnet_tvar_53[4][129] , 
	\_zy_simnet_tvar_53[4][128] , \_zy_simnet_tvar_53[4][127] , 
	\_zy_simnet_tvar_53[4][126] , \_zy_simnet_tvar_53[4][125] , 
	\_zy_simnet_tvar_53[4][124] , \_zy_simnet_tvar_53[4][123] , 
	\_zy_simnet_tvar_53[4][122] , \_zy_simnet_tvar_53[4][121] , 
	\_zy_simnet_tvar_53[4][120] , \_zy_simnet_tvar_53[4][119] , 
	\_zy_simnet_tvar_53[4][118] , \_zy_simnet_tvar_53[4][117] , 
	\_zy_simnet_tvar_53[4][116] , \_zy_simnet_tvar_53[4][115] , 
	\_zy_simnet_tvar_53[4][114] , \_zy_simnet_tvar_53[4][113] , 
	\_zy_simnet_tvar_53[4][112] , \_zy_simnet_tvar_53[4][111] , 
	\_zy_simnet_tvar_53[4][110] , \_zy_simnet_tvar_53[4][109] , 
	\_zy_simnet_tvar_53[4][108] , \_zy_simnet_tvar_53[4][107] , 
	\_zy_simnet_tvar_53[4][106] , \_zy_simnet_tvar_53[4][105] , 
	\_zy_simnet_tvar_53[4][104] , \_zy_simnet_tvar_53[4][103] , 
	\_zy_simnet_tvar_53[4][102] , \_zy_simnet_tvar_53[4][101] , 
	\_zy_simnet_tvar_53[4][100] , \_zy_simnet_tvar_53[4][99] , 
	\_zy_simnet_tvar_53[4][98] , \_zy_simnet_tvar_53[4][97] , 
	\_zy_simnet_tvar_53[4][96] , \_zy_simnet_tvar_53[4][95] , 
	\_zy_simnet_tvar_53[4][94] , \_zy_simnet_tvar_53[4][93] , 
	\_zy_simnet_tvar_53[4][92] , \_zy_simnet_tvar_53[4][91] , 
	\_zy_simnet_tvar_53[4][90] , \_zy_simnet_tvar_53[4][89] , 
	\_zy_simnet_tvar_53[4][88] , \_zy_simnet_tvar_53[4][87] , 
	\_zy_simnet_tvar_53[4][86] , \_zy_simnet_tvar_53[4][85] , 
	\_zy_simnet_tvar_53[4][84] , \_zy_simnet_tvar_53[4][83] , 
	\_zy_simnet_tvar_53[4][82] , \_zy_simnet_tvar_53[4][81] , 
	\_zy_simnet_tvar_53[4][80] , \_zy_simnet_tvar_53[4][79] , 
	\_zy_simnet_tvar_53[4][78] , \_zy_simnet_tvar_53[4][77] , 
	\_zy_simnet_tvar_53[4][76] , \_zy_simnet_tvar_53[4][75] , 
	\_zy_simnet_tvar_53[4][74] , \_zy_simnet_tvar_53[4][73] , 
	\_zy_simnet_tvar_53[4][72] , \_zy_simnet_tvar_53[4][71] , 
	\_zy_simnet_tvar_53[4][70] , \_zy_simnet_tvar_53[4][69] , 
	\_zy_simnet_tvar_53[4][68] , \_zy_simnet_tvar_53[4][67] , 
	\_zy_simnet_tvar_53[4][66] , \_zy_simnet_tvar_53[4][65] , 
	\_zy_simnet_tvar_53[4][64] , \_zy_simnet_tvar_53[4][63] , 
	\_zy_simnet_tvar_53[4][62] , \_zy_simnet_tvar_53[4][61] , 
	\_zy_simnet_tvar_53[4][60] , \_zy_simnet_tvar_53[4][59] , 
	\_zy_simnet_tvar_53[4][58] , \_zy_simnet_tvar_53[4][57] , 
	\_zy_simnet_tvar_53[4][56] , \_zy_simnet_tvar_53[4][55] , 
	\_zy_simnet_tvar_53[4][54] , \_zy_simnet_tvar_53[4][53] , 
	\_zy_simnet_tvar_53[4][52] , \_zy_simnet_tvar_53[4][51] , 
	\_zy_simnet_tvar_53[4][50] , \_zy_simnet_tvar_53[4][49] , 
	\_zy_simnet_tvar_53[4][48] , \_zy_simnet_tvar_53[4][47] , 
	\_zy_simnet_tvar_53[4][46] , \_zy_simnet_tvar_53[4][45] , 
	\_zy_simnet_tvar_53[4][44] , \_zy_simnet_tvar_53[4][43] , 
	\_zy_simnet_tvar_53[4][42] , \_zy_simnet_tvar_53[4][41] , 
	\_zy_simnet_tvar_53[4][40] , \_zy_simnet_tvar_53[4][39] , 
	\_zy_simnet_tvar_53[4][38] , \_zy_simnet_tvar_53[4][37] , 
	\_zy_simnet_tvar_53[4][36] , \_zy_simnet_tvar_53[4][35] , 
	\_zy_simnet_tvar_53[4][34] , \_zy_simnet_tvar_53[4][33] , 
	\_zy_simnet_tvar_53[4][32] , \_zy_simnet_tvar_53[4][31] , 
	\_zy_simnet_tvar_53[4][30] , \_zy_simnet_tvar_53[4][29] , 
	\_zy_simnet_tvar_53[4][28] , \_zy_simnet_tvar_53[4][27] , 
	\_zy_simnet_tvar_53[4][26] , \_zy_simnet_tvar_53[4][25] , 
	\_zy_simnet_tvar_53[4][24] , \_zy_simnet_tvar_53[4][23] , 
	\_zy_simnet_tvar_53[4][22] , \_zy_simnet_tvar_53[4][21] , 
	\_zy_simnet_tvar_53[4][20] , \_zy_simnet_tvar_53[4][19] , 
	\_zy_simnet_tvar_53[4][18] , \_zy_simnet_tvar_53[4][17] , 
	\_zy_simnet_tvar_53[4][16] , \_zy_simnet_tvar_53[4][15] , 
	\_zy_simnet_tvar_53[4][14] , \_zy_simnet_tvar_53[4][13] , 
	\_zy_simnet_tvar_53[4][12] , \_zy_simnet_tvar_53[4][11] , 
	\_zy_simnet_tvar_53[4][10] , \_zy_simnet_tvar_53[4][9] , 
	\_zy_simnet_tvar_53[4][8] , \_zy_simnet_tvar_53[4][7] , 
	\_zy_simnet_tvar_53[4][6] , \_zy_simnet_tvar_53[4][5] , 
	\_zy_simnet_tvar_53[4][4] , \_zy_simnet_tvar_53[4][3] , 
	\_zy_simnet_tvar_53[4][2] , \_zy_simnet_tvar_53[4][1] , 
	\_zy_simnet_tvar_53[4][0] , \_zy_simnet_tvar_53[3][271] , 
	\_zy_simnet_tvar_53[3][270] , \_zy_simnet_tvar_53[3][269] , 
	\_zy_simnet_tvar_53[3][268] , \_zy_simnet_tvar_53[3][267] , 
	\_zy_simnet_tvar_53[3][266] , \_zy_simnet_tvar_53[3][265] , 
	\_zy_simnet_tvar_53[3][264] , \_zy_simnet_tvar_53[3][263] , 
	\_zy_simnet_tvar_53[3][262] , \_zy_simnet_tvar_53[3][261] , 
	\_zy_simnet_tvar_53[3][260] , \_zy_simnet_tvar_53[3][259] , 
	\_zy_simnet_tvar_53[3][258] , \_zy_simnet_tvar_53[3][257] , 
	\_zy_simnet_tvar_53[3][256] , \_zy_simnet_tvar_53[3][255] , 
	\_zy_simnet_tvar_53[3][254] , \_zy_simnet_tvar_53[3][253] , 
	\_zy_simnet_tvar_53[3][252] , \_zy_simnet_tvar_53[3][251] , 
	\_zy_simnet_tvar_53[3][250] , \_zy_simnet_tvar_53[3][249] , 
	\_zy_simnet_tvar_53[3][248] , \_zy_simnet_tvar_53[3][247] , 
	\_zy_simnet_tvar_53[3][246] , \_zy_simnet_tvar_53[3][245] , 
	\_zy_simnet_tvar_53[3][244] , \_zy_simnet_tvar_53[3][243] , 
	\_zy_simnet_tvar_53[3][242] , \_zy_simnet_tvar_53[3][241] , 
	\_zy_simnet_tvar_53[3][240] , \_zy_simnet_tvar_53[3][239] , 
	\_zy_simnet_tvar_53[3][238] , \_zy_simnet_tvar_53[3][237] , 
	\_zy_simnet_tvar_53[3][236] , \_zy_simnet_tvar_53[3][235] , 
	\_zy_simnet_tvar_53[3][234] , \_zy_simnet_tvar_53[3][233] , 
	\_zy_simnet_tvar_53[3][232] , \_zy_simnet_tvar_53[3][231] , 
	\_zy_simnet_tvar_53[3][230] , \_zy_simnet_tvar_53[3][229] , 
	\_zy_simnet_tvar_53[3][228] , \_zy_simnet_tvar_53[3][227] , 
	\_zy_simnet_tvar_53[3][226] , \_zy_simnet_tvar_53[3][225] , 
	\_zy_simnet_tvar_53[3][224] , \_zy_simnet_tvar_53[3][223] , 
	\_zy_simnet_tvar_53[3][222] , \_zy_simnet_tvar_53[3][221] , 
	\_zy_simnet_tvar_53[3][220] , \_zy_simnet_tvar_53[3][219] , 
	\_zy_simnet_tvar_53[3][218] , \_zy_simnet_tvar_53[3][217] , 
	\_zy_simnet_tvar_53[3][216] , \_zy_simnet_tvar_53[3][215] , 
	\_zy_simnet_tvar_53[3][214] , \_zy_simnet_tvar_53[3][213] , 
	\_zy_simnet_tvar_53[3][212] , \_zy_simnet_tvar_53[3][211] , 
	\_zy_simnet_tvar_53[3][210] , \_zy_simnet_tvar_53[3][209] , 
	\_zy_simnet_tvar_53[3][208] , \_zy_simnet_tvar_53[3][207] , 
	\_zy_simnet_tvar_53[3][206] , \_zy_simnet_tvar_53[3][205] , 
	\_zy_simnet_tvar_53[3][204] , \_zy_simnet_tvar_53[3][203] , 
	\_zy_simnet_tvar_53[3][202] , \_zy_simnet_tvar_53[3][201] , 
	\_zy_simnet_tvar_53[3][200] , \_zy_simnet_tvar_53[3][199] , 
	\_zy_simnet_tvar_53[3][198] , \_zy_simnet_tvar_53[3][197] , 
	\_zy_simnet_tvar_53[3][196] , \_zy_simnet_tvar_53[3][195] , 
	\_zy_simnet_tvar_53[3][194] , \_zy_simnet_tvar_53[3][193] , 
	\_zy_simnet_tvar_53[3][192] , \_zy_simnet_tvar_53[3][191] , 
	\_zy_simnet_tvar_53[3][190] , \_zy_simnet_tvar_53[3][189] , 
	\_zy_simnet_tvar_53[3][188] , \_zy_simnet_tvar_53[3][187] , 
	\_zy_simnet_tvar_53[3][186] , \_zy_simnet_tvar_53[3][185] , 
	\_zy_simnet_tvar_53[3][184] , \_zy_simnet_tvar_53[3][183] , 
	\_zy_simnet_tvar_53[3][182] , \_zy_simnet_tvar_53[3][181] , 
	\_zy_simnet_tvar_53[3][180] , \_zy_simnet_tvar_53[3][179] , 
	\_zy_simnet_tvar_53[3][178] , \_zy_simnet_tvar_53[3][177] , 
	\_zy_simnet_tvar_53[3][176] , \_zy_simnet_tvar_53[3][175] , 
	\_zy_simnet_tvar_53[3][174] , \_zy_simnet_tvar_53[3][173] , 
	\_zy_simnet_tvar_53[3][172] , \_zy_simnet_tvar_53[3][171] , 
	\_zy_simnet_tvar_53[3][170] , \_zy_simnet_tvar_53[3][169] , 
	\_zy_simnet_tvar_53[3][168] , \_zy_simnet_tvar_53[3][167] , 
	\_zy_simnet_tvar_53[3][166] , \_zy_simnet_tvar_53[3][165] , 
	\_zy_simnet_tvar_53[3][164] , \_zy_simnet_tvar_53[3][163] , 
	\_zy_simnet_tvar_53[3][162] , \_zy_simnet_tvar_53[3][161] , 
	\_zy_simnet_tvar_53[3][160] , \_zy_simnet_tvar_53[3][159] , 
	\_zy_simnet_tvar_53[3][158] , \_zy_simnet_tvar_53[3][157] , 
	\_zy_simnet_tvar_53[3][156] , \_zy_simnet_tvar_53[3][155] , 
	\_zy_simnet_tvar_53[3][154] , \_zy_simnet_tvar_53[3][153] , 
	\_zy_simnet_tvar_53[3][152] , \_zy_simnet_tvar_53[3][151] , 
	\_zy_simnet_tvar_53[3][150] , \_zy_simnet_tvar_53[3][149] , 
	\_zy_simnet_tvar_53[3][148] , \_zy_simnet_tvar_53[3][147] , 
	\_zy_simnet_tvar_53[3][146] , \_zy_simnet_tvar_53[3][145] , 
	\_zy_simnet_tvar_53[3][144] , \_zy_simnet_tvar_53[3][143] , 
	\_zy_simnet_tvar_53[3][142] , \_zy_simnet_tvar_53[3][141] , 
	\_zy_simnet_tvar_53[3][140] , \_zy_simnet_tvar_53[3][139] , 
	\_zy_simnet_tvar_53[3][138] , \_zy_simnet_tvar_53[3][137] , 
	\_zy_simnet_tvar_53[3][136] , \_zy_simnet_tvar_53[3][135] , 
	\_zy_simnet_tvar_53[3][134] , \_zy_simnet_tvar_53[3][133] , 
	\_zy_simnet_tvar_53[3][132] , \_zy_simnet_tvar_53[3][131] , 
	\_zy_simnet_tvar_53[3][130] , \_zy_simnet_tvar_53[3][129] , 
	\_zy_simnet_tvar_53[3][128] , \_zy_simnet_tvar_53[3][127] , 
	\_zy_simnet_tvar_53[3][126] , \_zy_simnet_tvar_53[3][125] , 
	\_zy_simnet_tvar_53[3][124] , \_zy_simnet_tvar_53[3][123] , 
	\_zy_simnet_tvar_53[3][122] , \_zy_simnet_tvar_53[3][121] , 
	\_zy_simnet_tvar_53[3][120] , \_zy_simnet_tvar_53[3][119] , 
	\_zy_simnet_tvar_53[3][118] , \_zy_simnet_tvar_53[3][117] , 
	\_zy_simnet_tvar_53[3][116] , \_zy_simnet_tvar_53[3][115] , 
	\_zy_simnet_tvar_53[3][114] , \_zy_simnet_tvar_53[3][113] , 
	\_zy_simnet_tvar_53[3][112] , \_zy_simnet_tvar_53[3][111] , 
	\_zy_simnet_tvar_53[3][110] , \_zy_simnet_tvar_53[3][109] , 
	\_zy_simnet_tvar_53[3][108] , \_zy_simnet_tvar_53[3][107] , 
	\_zy_simnet_tvar_53[3][106] , \_zy_simnet_tvar_53[3][105] , 
	\_zy_simnet_tvar_53[3][104] , \_zy_simnet_tvar_53[3][103] , 
	\_zy_simnet_tvar_53[3][102] , \_zy_simnet_tvar_53[3][101] , 
	\_zy_simnet_tvar_53[3][100] , \_zy_simnet_tvar_53[3][99] , 
	\_zy_simnet_tvar_53[3][98] , \_zy_simnet_tvar_53[3][97] , 
	\_zy_simnet_tvar_53[3][96] , \_zy_simnet_tvar_53[3][95] , 
	\_zy_simnet_tvar_53[3][94] , \_zy_simnet_tvar_53[3][93] , 
	\_zy_simnet_tvar_53[3][92] , \_zy_simnet_tvar_53[3][91] , 
	\_zy_simnet_tvar_53[3][90] , \_zy_simnet_tvar_53[3][89] , 
	\_zy_simnet_tvar_53[3][88] , \_zy_simnet_tvar_53[3][87] , 
	\_zy_simnet_tvar_53[3][86] , \_zy_simnet_tvar_53[3][85] , 
	\_zy_simnet_tvar_53[3][84] , \_zy_simnet_tvar_53[3][83] , 
	\_zy_simnet_tvar_53[3][82] , \_zy_simnet_tvar_53[3][81] , 
	\_zy_simnet_tvar_53[3][80] , \_zy_simnet_tvar_53[3][79] , 
	\_zy_simnet_tvar_53[3][78] , \_zy_simnet_tvar_53[3][77] , 
	\_zy_simnet_tvar_53[3][76] , \_zy_simnet_tvar_53[3][75] , 
	\_zy_simnet_tvar_53[3][74] , \_zy_simnet_tvar_53[3][73] , 
	\_zy_simnet_tvar_53[3][72] , \_zy_simnet_tvar_53[3][71] , 
	\_zy_simnet_tvar_53[3][70] , \_zy_simnet_tvar_53[3][69] , 
	\_zy_simnet_tvar_53[3][68] , \_zy_simnet_tvar_53[3][67] , 
	\_zy_simnet_tvar_53[3][66] , \_zy_simnet_tvar_53[3][65] , 
	\_zy_simnet_tvar_53[3][64] , \_zy_simnet_tvar_53[3][63] , 
	\_zy_simnet_tvar_53[3][62] , \_zy_simnet_tvar_53[3][61] , 
	\_zy_simnet_tvar_53[3][60] , \_zy_simnet_tvar_53[3][59] , 
	\_zy_simnet_tvar_53[3][58] , \_zy_simnet_tvar_53[3][57] , 
	\_zy_simnet_tvar_53[3][56] , \_zy_simnet_tvar_53[3][55] , 
	\_zy_simnet_tvar_53[3][54] , \_zy_simnet_tvar_53[3][53] , 
	\_zy_simnet_tvar_53[3][52] , \_zy_simnet_tvar_53[3][51] , 
	\_zy_simnet_tvar_53[3][50] , \_zy_simnet_tvar_53[3][49] , 
	\_zy_simnet_tvar_53[3][48] , \_zy_simnet_tvar_53[3][47] , 
	\_zy_simnet_tvar_53[3][46] , \_zy_simnet_tvar_53[3][45] , 
	\_zy_simnet_tvar_53[3][44] , \_zy_simnet_tvar_53[3][43] , 
	\_zy_simnet_tvar_53[3][42] , \_zy_simnet_tvar_53[3][41] , 
	\_zy_simnet_tvar_53[3][40] , \_zy_simnet_tvar_53[3][39] , 
	\_zy_simnet_tvar_53[3][38] , \_zy_simnet_tvar_53[3][37] , 
	\_zy_simnet_tvar_53[3][36] , \_zy_simnet_tvar_53[3][35] , 
	\_zy_simnet_tvar_53[3][34] , \_zy_simnet_tvar_53[3][33] , 
	\_zy_simnet_tvar_53[3][32] , \_zy_simnet_tvar_53[3][31] , 
	\_zy_simnet_tvar_53[3][30] , \_zy_simnet_tvar_53[3][29] , 
	\_zy_simnet_tvar_53[3][28] , \_zy_simnet_tvar_53[3][27] , 
	\_zy_simnet_tvar_53[3][26] , \_zy_simnet_tvar_53[3][25] , 
	\_zy_simnet_tvar_53[3][24] , \_zy_simnet_tvar_53[3][23] , 
	\_zy_simnet_tvar_53[3][22] , \_zy_simnet_tvar_53[3][21] , 
	\_zy_simnet_tvar_53[3][20] , \_zy_simnet_tvar_53[3][19] , 
	\_zy_simnet_tvar_53[3][18] , \_zy_simnet_tvar_53[3][17] , 
	\_zy_simnet_tvar_53[3][16] , \_zy_simnet_tvar_53[3][15] , 
	\_zy_simnet_tvar_53[3][14] , \_zy_simnet_tvar_53[3][13] , 
	\_zy_simnet_tvar_53[3][12] , \_zy_simnet_tvar_53[3][11] , 
	\_zy_simnet_tvar_53[3][10] , \_zy_simnet_tvar_53[3][9] , 
	\_zy_simnet_tvar_53[3][8] , \_zy_simnet_tvar_53[3][7] , 
	\_zy_simnet_tvar_53[3][6] , \_zy_simnet_tvar_53[3][5] , 
	\_zy_simnet_tvar_53[3][4] , \_zy_simnet_tvar_53[3][3] , 
	\_zy_simnet_tvar_53[3][2] , \_zy_simnet_tvar_53[3][1] , 
	\_zy_simnet_tvar_53[3][0] , \_zy_simnet_tvar_53[2][271] , 
	\_zy_simnet_tvar_53[2][270] , \_zy_simnet_tvar_53[2][269] , 
	\_zy_simnet_tvar_53[2][268] , \_zy_simnet_tvar_53[2][267] , 
	\_zy_simnet_tvar_53[2][266] , \_zy_simnet_tvar_53[2][265] , 
	\_zy_simnet_tvar_53[2][264] , \_zy_simnet_tvar_53[2][263] , 
	\_zy_simnet_tvar_53[2][262] , \_zy_simnet_tvar_53[2][261] , 
	\_zy_simnet_tvar_53[2][260] , \_zy_simnet_tvar_53[2][259] , 
	\_zy_simnet_tvar_53[2][258] , \_zy_simnet_tvar_53[2][257] , 
	\_zy_simnet_tvar_53[2][256] , \_zy_simnet_tvar_53[2][255] , 
	\_zy_simnet_tvar_53[2][254] , \_zy_simnet_tvar_53[2][253] , 
	\_zy_simnet_tvar_53[2][252] , \_zy_simnet_tvar_53[2][251] , 
	\_zy_simnet_tvar_53[2][250] , \_zy_simnet_tvar_53[2][249] , 
	\_zy_simnet_tvar_53[2][248] , \_zy_simnet_tvar_53[2][247] , 
	\_zy_simnet_tvar_53[2][246] , \_zy_simnet_tvar_53[2][245] , 
	\_zy_simnet_tvar_53[2][244] , \_zy_simnet_tvar_53[2][243] , 
	\_zy_simnet_tvar_53[2][242] , \_zy_simnet_tvar_53[2][241] , 
	\_zy_simnet_tvar_53[2][240] , \_zy_simnet_tvar_53[2][239] , 
	\_zy_simnet_tvar_53[2][238] , \_zy_simnet_tvar_53[2][237] , 
	\_zy_simnet_tvar_53[2][236] , \_zy_simnet_tvar_53[2][235] , 
	\_zy_simnet_tvar_53[2][234] , \_zy_simnet_tvar_53[2][233] , 
	\_zy_simnet_tvar_53[2][232] , \_zy_simnet_tvar_53[2][231] , 
	\_zy_simnet_tvar_53[2][230] , \_zy_simnet_tvar_53[2][229] , 
	\_zy_simnet_tvar_53[2][228] , \_zy_simnet_tvar_53[2][227] , 
	\_zy_simnet_tvar_53[2][226] , \_zy_simnet_tvar_53[2][225] , 
	\_zy_simnet_tvar_53[2][224] , \_zy_simnet_tvar_53[2][223] , 
	\_zy_simnet_tvar_53[2][222] , \_zy_simnet_tvar_53[2][221] , 
	\_zy_simnet_tvar_53[2][220] , \_zy_simnet_tvar_53[2][219] , 
	\_zy_simnet_tvar_53[2][218] , \_zy_simnet_tvar_53[2][217] , 
	\_zy_simnet_tvar_53[2][216] , \_zy_simnet_tvar_53[2][215] , 
	\_zy_simnet_tvar_53[2][214] , \_zy_simnet_tvar_53[2][213] , 
	\_zy_simnet_tvar_53[2][212] , \_zy_simnet_tvar_53[2][211] , 
	\_zy_simnet_tvar_53[2][210] , \_zy_simnet_tvar_53[2][209] , 
	\_zy_simnet_tvar_53[2][208] , \_zy_simnet_tvar_53[2][207] , 
	\_zy_simnet_tvar_53[2][206] , \_zy_simnet_tvar_53[2][205] , 
	\_zy_simnet_tvar_53[2][204] , \_zy_simnet_tvar_53[2][203] , 
	\_zy_simnet_tvar_53[2][202] , \_zy_simnet_tvar_53[2][201] , 
	\_zy_simnet_tvar_53[2][200] , \_zy_simnet_tvar_53[2][199] , 
	\_zy_simnet_tvar_53[2][198] , \_zy_simnet_tvar_53[2][197] , 
	\_zy_simnet_tvar_53[2][196] , \_zy_simnet_tvar_53[2][195] , 
	\_zy_simnet_tvar_53[2][194] , \_zy_simnet_tvar_53[2][193] , 
	\_zy_simnet_tvar_53[2][192] , \_zy_simnet_tvar_53[2][191] , 
	\_zy_simnet_tvar_53[2][190] , \_zy_simnet_tvar_53[2][189] , 
	\_zy_simnet_tvar_53[2][188] , \_zy_simnet_tvar_53[2][187] , 
	\_zy_simnet_tvar_53[2][186] , \_zy_simnet_tvar_53[2][185] , 
	\_zy_simnet_tvar_53[2][184] , \_zy_simnet_tvar_53[2][183] , 
	\_zy_simnet_tvar_53[2][182] , \_zy_simnet_tvar_53[2][181] , 
	\_zy_simnet_tvar_53[2][180] , \_zy_simnet_tvar_53[2][179] , 
	\_zy_simnet_tvar_53[2][178] , \_zy_simnet_tvar_53[2][177] , 
	\_zy_simnet_tvar_53[2][176] , \_zy_simnet_tvar_53[2][175] , 
	\_zy_simnet_tvar_53[2][174] , \_zy_simnet_tvar_53[2][173] , 
	\_zy_simnet_tvar_53[2][172] , \_zy_simnet_tvar_53[2][171] , 
	\_zy_simnet_tvar_53[2][170] , \_zy_simnet_tvar_53[2][169] , 
	\_zy_simnet_tvar_53[2][168] , \_zy_simnet_tvar_53[2][167] , 
	\_zy_simnet_tvar_53[2][166] , \_zy_simnet_tvar_53[2][165] , 
	\_zy_simnet_tvar_53[2][164] , \_zy_simnet_tvar_53[2][163] , 
	\_zy_simnet_tvar_53[2][162] , \_zy_simnet_tvar_53[2][161] , 
	\_zy_simnet_tvar_53[2][160] , \_zy_simnet_tvar_53[2][159] , 
	\_zy_simnet_tvar_53[2][158] , \_zy_simnet_tvar_53[2][157] , 
	\_zy_simnet_tvar_53[2][156] , \_zy_simnet_tvar_53[2][155] , 
	\_zy_simnet_tvar_53[2][154] , \_zy_simnet_tvar_53[2][153] , 
	\_zy_simnet_tvar_53[2][152] , \_zy_simnet_tvar_53[2][151] , 
	\_zy_simnet_tvar_53[2][150] , \_zy_simnet_tvar_53[2][149] , 
	\_zy_simnet_tvar_53[2][148] , \_zy_simnet_tvar_53[2][147] , 
	\_zy_simnet_tvar_53[2][146] , \_zy_simnet_tvar_53[2][145] , 
	\_zy_simnet_tvar_53[2][144] , \_zy_simnet_tvar_53[2][143] , 
	\_zy_simnet_tvar_53[2][142] , \_zy_simnet_tvar_53[2][141] , 
	\_zy_simnet_tvar_53[2][140] , \_zy_simnet_tvar_53[2][139] , 
	\_zy_simnet_tvar_53[2][138] , \_zy_simnet_tvar_53[2][137] , 
	\_zy_simnet_tvar_53[2][136] , \_zy_simnet_tvar_53[2][135] , 
	\_zy_simnet_tvar_53[2][134] , \_zy_simnet_tvar_53[2][133] , 
	\_zy_simnet_tvar_53[2][132] , \_zy_simnet_tvar_53[2][131] , 
	\_zy_simnet_tvar_53[2][130] , \_zy_simnet_tvar_53[2][129] , 
	\_zy_simnet_tvar_53[2][128] , \_zy_simnet_tvar_53[2][127] , 
	\_zy_simnet_tvar_53[2][126] , \_zy_simnet_tvar_53[2][125] , 
	\_zy_simnet_tvar_53[2][124] , \_zy_simnet_tvar_53[2][123] , 
	\_zy_simnet_tvar_53[2][122] , \_zy_simnet_tvar_53[2][121] , 
	\_zy_simnet_tvar_53[2][120] , \_zy_simnet_tvar_53[2][119] , 
	\_zy_simnet_tvar_53[2][118] , \_zy_simnet_tvar_53[2][117] , 
	\_zy_simnet_tvar_53[2][116] , \_zy_simnet_tvar_53[2][115] , 
	\_zy_simnet_tvar_53[2][114] , \_zy_simnet_tvar_53[2][113] , 
	\_zy_simnet_tvar_53[2][112] , \_zy_simnet_tvar_53[2][111] , 
	\_zy_simnet_tvar_53[2][110] , \_zy_simnet_tvar_53[2][109] , 
	\_zy_simnet_tvar_53[2][108] , \_zy_simnet_tvar_53[2][107] , 
	\_zy_simnet_tvar_53[2][106] , \_zy_simnet_tvar_53[2][105] , 
	\_zy_simnet_tvar_53[2][104] , \_zy_simnet_tvar_53[2][103] , 
	\_zy_simnet_tvar_53[2][102] , \_zy_simnet_tvar_53[2][101] , 
	\_zy_simnet_tvar_53[2][100] , \_zy_simnet_tvar_53[2][99] , 
	\_zy_simnet_tvar_53[2][98] , \_zy_simnet_tvar_53[2][97] , 
	\_zy_simnet_tvar_53[2][96] , \_zy_simnet_tvar_53[2][95] , 
	\_zy_simnet_tvar_53[2][94] , \_zy_simnet_tvar_53[2][93] , 
	\_zy_simnet_tvar_53[2][92] , \_zy_simnet_tvar_53[2][91] , 
	\_zy_simnet_tvar_53[2][90] , \_zy_simnet_tvar_53[2][89] , 
	\_zy_simnet_tvar_53[2][88] , \_zy_simnet_tvar_53[2][87] , 
	\_zy_simnet_tvar_53[2][86] , \_zy_simnet_tvar_53[2][85] , 
	\_zy_simnet_tvar_53[2][84] , \_zy_simnet_tvar_53[2][83] , 
	\_zy_simnet_tvar_53[2][82] , \_zy_simnet_tvar_53[2][81] , 
	\_zy_simnet_tvar_53[2][80] , \_zy_simnet_tvar_53[2][79] , 
	\_zy_simnet_tvar_53[2][78] , \_zy_simnet_tvar_53[2][77] , 
	\_zy_simnet_tvar_53[2][76] , \_zy_simnet_tvar_53[2][75] , 
	\_zy_simnet_tvar_53[2][74] , \_zy_simnet_tvar_53[2][73] , 
	\_zy_simnet_tvar_53[2][72] , \_zy_simnet_tvar_53[2][71] , 
	\_zy_simnet_tvar_53[2][70] , \_zy_simnet_tvar_53[2][69] , 
	\_zy_simnet_tvar_53[2][68] , \_zy_simnet_tvar_53[2][67] , 
	\_zy_simnet_tvar_53[2][66] , \_zy_simnet_tvar_53[2][65] , 
	\_zy_simnet_tvar_53[2][64] , \_zy_simnet_tvar_53[2][63] , 
	\_zy_simnet_tvar_53[2][62] , \_zy_simnet_tvar_53[2][61] , 
	\_zy_simnet_tvar_53[2][60] , \_zy_simnet_tvar_53[2][59] , 
	\_zy_simnet_tvar_53[2][58] , \_zy_simnet_tvar_53[2][57] , 
	\_zy_simnet_tvar_53[2][56] , \_zy_simnet_tvar_53[2][55] , 
	\_zy_simnet_tvar_53[2][54] , \_zy_simnet_tvar_53[2][53] , 
	\_zy_simnet_tvar_53[2][52] , \_zy_simnet_tvar_53[2][51] , 
	\_zy_simnet_tvar_53[2][50] , \_zy_simnet_tvar_53[2][49] , 
	\_zy_simnet_tvar_53[2][48] , \_zy_simnet_tvar_53[2][47] , 
	\_zy_simnet_tvar_53[2][46] , \_zy_simnet_tvar_53[2][45] , 
	\_zy_simnet_tvar_53[2][44] , \_zy_simnet_tvar_53[2][43] , 
	\_zy_simnet_tvar_53[2][42] , \_zy_simnet_tvar_53[2][41] , 
	\_zy_simnet_tvar_53[2][40] , \_zy_simnet_tvar_53[2][39] , 
	\_zy_simnet_tvar_53[2][38] , \_zy_simnet_tvar_53[2][37] , 
	\_zy_simnet_tvar_53[2][36] , \_zy_simnet_tvar_53[2][35] , 
	\_zy_simnet_tvar_53[2][34] , \_zy_simnet_tvar_53[2][33] , 
	\_zy_simnet_tvar_53[2][32] , \_zy_simnet_tvar_53[2][31] , 
	\_zy_simnet_tvar_53[2][30] , \_zy_simnet_tvar_53[2][29] , 
	\_zy_simnet_tvar_53[2][28] , \_zy_simnet_tvar_53[2][27] , 
	\_zy_simnet_tvar_53[2][26] , \_zy_simnet_tvar_53[2][25] , 
	\_zy_simnet_tvar_53[2][24] , \_zy_simnet_tvar_53[2][23] , 
	\_zy_simnet_tvar_53[2][22] , \_zy_simnet_tvar_53[2][21] , 
	\_zy_simnet_tvar_53[2][20] , \_zy_simnet_tvar_53[2][19] , 
	\_zy_simnet_tvar_53[2][18] , \_zy_simnet_tvar_53[2][17] , 
	\_zy_simnet_tvar_53[2][16] , \_zy_simnet_tvar_53[2][15] , 
	\_zy_simnet_tvar_53[2][14] , \_zy_simnet_tvar_53[2][13] , 
	\_zy_simnet_tvar_53[2][12] , \_zy_simnet_tvar_53[2][11] , 
	\_zy_simnet_tvar_53[2][10] , \_zy_simnet_tvar_53[2][9] , 
	\_zy_simnet_tvar_53[2][8] , \_zy_simnet_tvar_53[2][7] , 
	\_zy_simnet_tvar_53[2][6] , \_zy_simnet_tvar_53[2][5] , 
	\_zy_simnet_tvar_53[2][4] , \_zy_simnet_tvar_53[2][3] , 
	\_zy_simnet_tvar_53[2][2] , \_zy_simnet_tvar_53[2][1] , 
	\_zy_simnet_tvar_53[2][0] , \_zy_simnet_tvar_53[1][271] , 
	\_zy_simnet_tvar_53[1][270] , \_zy_simnet_tvar_53[1][269] , 
	\_zy_simnet_tvar_53[1][268] , \_zy_simnet_tvar_53[1][267] , 
	\_zy_simnet_tvar_53[1][266] , \_zy_simnet_tvar_53[1][265] , 
	\_zy_simnet_tvar_53[1][264] , \_zy_simnet_tvar_53[1][263] , 
	\_zy_simnet_tvar_53[1][262] , \_zy_simnet_tvar_53[1][261] , 
	\_zy_simnet_tvar_53[1][260] , \_zy_simnet_tvar_53[1][259] , 
	\_zy_simnet_tvar_53[1][258] , \_zy_simnet_tvar_53[1][257] , 
	\_zy_simnet_tvar_53[1][256] , \_zy_simnet_tvar_53[1][255] , 
	\_zy_simnet_tvar_53[1][254] , \_zy_simnet_tvar_53[1][253] , 
	\_zy_simnet_tvar_53[1][252] , \_zy_simnet_tvar_53[1][251] , 
	\_zy_simnet_tvar_53[1][250] , \_zy_simnet_tvar_53[1][249] , 
	\_zy_simnet_tvar_53[1][248] , \_zy_simnet_tvar_53[1][247] , 
	\_zy_simnet_tvar_53[1][246] , \_zy_simnet_tvar_53[1][245] , 
	\_zy_simnet_tvar_53[1][244] , \_zy_simnet_tvar_53[1][243] , 
	\_zy_simnet_tvar_53[1][242] , \_zy_simnet_tvar_53[1][241] , 
	\_zy_simnet_tvar_53[1][240] , \_zy_simnet_tvar_53[1][239] , 
	\_zy_simnet_tvar_53[1][238] , \_zy_simnet_tvar_53[1][237] , 
	\_zy_simnet_tvar_53[1][236] , \_zy_simnet_tvar_53[1][235] , 
	\_zy_simnet_tvar_53[1][234] , \_zy_simnet_tvar_53[1][233] , 
	\_zy_simnet_tvar_53[1][232] , \_zy_simnet_tvar_53[1][231] , 
	\_zy_simnet_tvar_53[1][230] , \_zy_simnet_tvar_53[1][229] , 
	\_zy_simnet_tvar_53[1][228] , \_zy_simnet_tvar_53[1][227] , 
	\_zy_simnet_tvar_53[1][226] , \_zy_simnet_tvar_53[1][225] , 
	\_zy_simnet_tvar_53[1][224] , \_zy_simnet_tvar_53[1][223] , 
	\_zy_simnet_tvar_53[1][222] , \_zy_simnet_tvar_53[1][221] , 
	\_zy_simnet_tvar_53[1][220] , \_zy_simnet_tvar_53[1][219] , 
	\_zy_simnet_tvar_53[1][218] , \_zy_simnet_tvar_53[1][217] , 
	\_zy_simnet_tvar_53[1][216] , \_zy_simnet_tvar_53[1][215] , 
	\_zy_simnet_tvar_53[1][214] , \_zy_simnet_tvar_53[1][213] , 
	\_zy_simnet_tvar_53[1][212] , \_zy_simnet_tvar_53[1][211] , 
	\_zy_simnet_tvar_53[1][210] , \_zy_simnet_tvar_53[1][209] , 
	\_zy_simnet_tvar_53[1][208] , \_zy_simnet_tvar_53[1][207] , 
	\_zy_simnet_tvar_53[1][206] , \_zy_simnet_tvar_53[1][205] , 
	\_zy_simnet_tvar_53[1][204] , \_zy_simnet_tvar_53[1][203] , 
	\_zy_simnet_tvar_53[1][202] , \_zy_simnet_tvar_53[1][201] , 
	\_zy_simnet_tvar_53[1][200] , \_zy_simnet_tvar_53[1][199] , 
	\_zy_simnet_tvar_53[1][198] , \_zy_simnet_tvar_53[1][197] , 
	\_zy_simnet_tvar_53[1][196] , \_zy_simnet_tvar_53[1][195] , 
	\_zy_simnet_tvar_53[1][194] , \_zy_simnet_tvar_53[1][193] , 
	\_zy_simnet_tvar_53[1][192] , \_zy_simnet_tvar_53[1][191] , 
	\_zy_simnet_tvar_53[1][190] , \_zy_simnet_tvar_53[1][189] , 
	\_zy_simnet_tvar_53[1][188] , \_zy_simnet_tvar_53[1][187] , 
	\_zy_simnet_tvar_53[1][186] , \_zy_simnet_tvar_53[1][185] , 
	\_zy_simnet_tvar_53[1][184] , \_zy_simnet_tvar_53[1][183] , 
	\_zy_simnet_tvar_53[1][182] , \_zy_simnet_tvar_53[1][181] , 
	\_zy_simnet_tvar_53[1][180] , \_zy_simnet_tvar_53[1][179] , 
	\_zy_simnet_tvar_53[1][178] , \_zy_simnet_tvar_53[1][177] , 
	\_zy_simnet_tvar_53[1][176] , \_zy_simnet_tvar_53[1][175] , 
	\_zy_simnet_tvar_53[1][174] , \_zy_simnet_tvar_53[1][173] , 
	\_zy_simnet_tvar_53[1][172] , \_zy_simnet_tvar_53[1][171] , 
	\_zy_simnet_tvar_53[1][170] , \_zy_simnet_tvar_53[1][169] , 
	\_zy_simnet_tvar_53[1][168] , \_zy_simnet_tvar_53[1][167] , 
	\_zy_simnet_tvar_53[1][166] , \_zy_simnet_tvar_53[1][165] , 
	\_zy_simnet_tvar_53[1][164] , \_zy_simnet_tvar_53[1][163] , 
	\_zy_simnet_tvar_53[1][162] , \_zy_simnet_tvar_53[1][161] , 
	\_zy_simnet_tvar_53[1][160] , \_zy_simnet_tvar_53[1][159] , 
	\_zy_simnet_tvar_53[1][158] , \_zy_simnet_tvar_53[1][157] , 
	\_zy_simnet_tvar_53[1][156] , \_zy_simnet_tvar_53[1][155] , 
	\_zy_simnet_tvar_53[1][154] , \_zy_simnet_tvar_53[1][153] , 
	\_zy_simnet_tvar_53[1][152] , \_zy_simnet_tvar_53[1][151] , 
	\_zy_simnet_tvar_53[1][150] , \_zy_simnet_tvar_53[1][149] , 
	\_zy_simnet_tvar_53[1][148] , \_zy_simnet_tvar_53[1][147] , 
	\_zy_simnet_tvar_53[1][146] , \_zy_simnet_tvar_53[1][145] , 
	\_zy_simnet_tvar_53[1][144] , \_zy_simnet_tvar_53[1][143] , 
	\_zy_simnet_tvar_53[1][142] , \_zy_simnet_tvar_53[1][141] , 
	\_zy_simnet_tvar_53[1][140] , \_zy_simnet_tvar_53[1][139] , 
	\_zy_simnet_tvar_53[1][138] , \_zy_simnet_tvar_53[1][137] , 
	\_zy_simnet_tvar_53[1][136] , \_zy_simnet_tvar_53[1][135] , 
	\_zy_simnet_tvar_53[1][134] , \_zy_simnet_tvar_53[1][133] , 
	\_zy_simnet_tvar_53[1][132] , \_zy_simnet_tvar_53[1][131] , 
	\_zy_simnet_tvar_53[1][130] , \_zy_simnet_tvar_53[1][129] , 
	\_zy_simnet_tvar_53[1][128] , \_zy_simnet_tvar_53[1][127] , 
	\_zy_simnet_tvar_53[1][126] , \_zy_simnet_tvar_53[1][125] , 
	\_zy_simnet_tvar_53[1][124] , \_zy_simnet_tvar_53[1][123] , 
	\_zy_simnet_tvar_53[1][122] , \_zy_simnet_tvar_53[1][121] , 
	\_zy_simnet_tvar_53[1][120] , \_zy_simnet_tvar_53[1][119] , 
	\_zy_simnet_tvar_53[1][118] , \_zy_simnet_tvar_53[1][117] , 
	\_zy_simnet_tvar_53[1][116] , \_zy_simnet_tvar_53[1][115] , 
	\_zy_simnet_tvar_53[1][114] , \_zy_simnet_tvar_53[1][113] , 
	\_zy_simnet_tvar_53[1][112] , \_zy_simnet_tvar_53[1][111] , 
	\_zy_simnet_tvar_53[1][110] , \_zy_simnet_tvar_53[1][109] , 
	\_zy_simnet_tvar_53[1][108] , \_zy_simnet_tvar_53[1][107] , 
	\_zy_simnet_tvar_53[1][106] , \_zy_simnet_tvar_53[1][105] , 
	\_zy_simnet_tvar_53[1][104] , \_zy_simnet_tvar_53[1][103] , 
	\_zy_simnet_tvar_53[1][102] , \_zy_simnet_tvar_53[1][101] , 
	\_zy_simnet_tvar_53[1][100] , \_zy_simnet_tvar_53[1][99] , 
	\_zy_simnet_tvar_53[1][98] , \_zy_simnet_tvar_53[1][97] , 
	\_zy_simnet_tvar_53[1][96] , \_zy_simnet_tvar_53[1][95] , 
	\_zy_simnet_tvar_53[1][94] , \_zy_simnet_tvar_53[1][93] , 
	\_zy_simnet_tvar_53[1][92] , \_zy_simnet_tvar_53[1][91] , 
	\_zy_simnet_tvar_53[1][90] , \_zy_simnet_tvar_53[1][89] , 
	\_zy_simnet_tvar_53[1][88] , \_zy_simnet_tvar_53[1][87] , 
	\_zy_simnet_tvar_53[1][86] , \_zy_simnet_tvar_53[1][85] , 
	\_zy_simnet_tvar_53[1][84] , \_zy_simnet_tvar_53[1][83] , 
	\_zy_simnet_tvar_53[1][82] , \_zy_simnet_tvar_53[1][81] , 
	\_zy_simnet_tvar_53[1][80] , \_zy_simnet_tvar_53[1][79] , 
	\_zy_simnet_tvar_53[1][78] , \_zy_simnet_tvar_53[1][77] , 
	\_zy_simnet_tvar_53[1][76] , \_zy_simnet_tvar_53[1][75] , 
	\_zy_simnet_tvar_53[1][74] , \_zy_simnet_tvar_53[1][73] , 
	\_zy_simnet_tvar_53[1][72] , \_zy_simnet_tvar_53[1][71] , 
	\_zy_simnet_tvar_53[1][70] , \_zy_simnet_tvar_53[1][69] , 
	\_zy_simnet_tvar_53[1][68] , \_zy_simnet_tvar_53[1][67] , 
	\_zy_simnet_tvar_53[1][66] , \_zy_simnet_tvar_53[1][65] , 
	\_zy_simnet_tvar_53[1][64] , \_zy_simnet_tvar_53[1][63] , 
	\_zy_simnet_tvar_53[1][62] , \_zy_simnet_tvar_53[1][61] , 
	\_zy_simnet_tvar_53[1][60] , \_zy_simnet_tvar_53[1][59] , 
	\_zy_simnet_tvar_53[1][58] , \_zy_simnet_tvar_53[1][57] , 
	\_zy_simnet_tvar_53[1][56] , \_zy_simnet_tvar_53[1][55] , 
	\_zy_simnet_tvar_53[1][54] , \_zy_simnet_tvar_53[1][53] , 
	\_zy_simnet_tvar_53[1][52] , \_zy_simnet_tvar_53[1][51] , 
	\_zy_simnet_tvar_53[1][50] , \_zy_simnet_tvar_53[1][49] , 
	\_zy_simnet_tvar_53[1][48] , \_zy_simnet_tvar_53[1][47] , 
	\_zy_simnet_tvar_53[1][46] , \_zy_simnet_tvar_53[1][45] , 
	\_zy_simnet_tvar_53[1][44] , \_zy_simnet_tvar_53[1][43] , 
	\_zy_simnet_tvar_53[1][42] , \_zy_simnet_tvar_53[1][41] , 
	\_zy_simnet_tvar_53[1][40] , \_zy_simnet_tvar_53[1][39] , 
	\_zy_simnet_tvar_53[1][38] , \_zy_simnet_tvar_53[1][37] , 
	\_zy_simnet_tvar_53[1][36] , \_zy_simnet_tvar_53[1][35] , 
	\_zy_simnet_tvar_53[1][34] , \_zy_simnet_tvar_53[1][33] , 
	\_zy_simnet_tvar_53[1][32] , \_zy_simnet_tvar_53[1][31] , 
	\_zy_simnet_tvar_53[1][30] , \_zy_simnet_tvar_53[1][29] , 
	\_zy_simnet_tvar_53[1][28] , \_zy_simnet_tvar_53[1][27] , 
	\_zy_simnet_tvar_53[1][26] , \_zy_simnet_tvar_53[1][25] , 
	\_zy_simnet_tvar_53[1][24] , \_zy_simnet_tvar_53[1][23] , 
	\_zy_simnet_tvar_53[1][22] , \_zy_simnet_tvar_53[1][21] , 
	\_zy_simnet_tvar_53[1][20] , \_zy_simnet_tvar_53[1][19] , 
	\_zy_simnet_tvar_53[1][18] , \_zy_simnet_tvar_53[1][17] , 
	\_zy_simnet_tvar_53[1][16] , \_zy_simnet_tvar_53[1][15] , 
	\_zy_simnet_tvar_53[1][14] , \_zy_simnet_tvar_53[1][13] , 
	\_zy_simnet_tvar_53[1][12] , \_zy_simnet_tvar_53[1][11] , 
	\_zy_simnet_tvar_53[1][10] , \_zy_simnet_tvar_53[1][9] , 
	\_zy_simnet_tvar_53[1][8] , \_zy_simnet_tvar_53[1][7] , 
	\_zy_simnet_tvar_53[1][6] , \_zy_simnet_tvar_53[1][5] , 
	\_zy_simnet_tvar_53[1][4] , \_zy_simnet_tvar_53[1][3] , 
	\_zy_simnet_tvar_53[1][2] , \_zy_simnet_tvar_53[1][1] , 
	\_zy_simnet_tvar_53[1][0] , \_zy_simnet_tvar_53[0][271] , 
	\_zy_simnet_tvar_53[0][270] , \_zy_simnet_tvar_53[0][269] , 
	\_zy_simnet_tvar_53[0][268] , \_zy_simnet_tvar_53[0][267] , 
	\_zy_simnet_tvar_53[0][266] , \_zy_simnet_tvar_53[0][265] , 
	\_zy_simnet_tvar_53[0][264] , \_zy_simnet_tvar_53[0][263] , 
	\_zy_simnet_tvar_53[0][262] , \_zy_simnet_tvar_53[0][261] , 
	\_zy_simnet_tvar_53[0][260] , \_zy_simnet_tvar_53[0][259] , 
	\_zy_simnet_tvar_53[0][258] , \_zy_simnet_tvar_53[0][257] , 
	\_zy_simnet_tvar_53[0][256] , \_zy_simnet_tvar_53[0][255] , 
	\_zy_simnet_tvar_53[0][254] , \_zy_simnet_tvar_53[0][253] , 
	\_zy_simnet_tvar_53[0][252] , \_zy_simnet_tvar_53[0][251] , 
	\_zy_simnet_tvar_53[0][250] , \_zy_simnet_tvar_53[0][249] , 
	\_zy_simnet_tvar_53[0][248] , \_zy_simnet_tvar_53[0][247] , 
	\_zy_simnet_tvar_53[0][246] , \_zy_simnet_tvar_53[0][245] , 
	\_zy_simnet_tvar_53[0][244] , \_zy_simnet_tvar_53[0][243] , 
	\_zy_simnet_tvar_53[0][242] , \_zy_simnet_tvar_53[0][241] , 
	\_zy_simnet_tvar_53[0][240] , \_zy_simnet_tvar_53[0][239] , 
	\_zy_simnet_tvar_53[0][238] , \_zy_simnet_tvar_53[0][237] , 
	\_zy_simnet_tvar_53[0][236] , \_zy_simnet_tvar_53[0][235] , 
	\_zy_simnet_tvar_53[0][234] , \_zy_simnet_tvar_53[0][233] , 
	\_zy_simnet_tvar_53[0][232] , \_zy_simnet_tvar_53[0][231] , 
	\_zy_simnet_tvar_53[0][230] , \_zy_simnet_tvar_53[0][229] , 
	\_zy_simnet_tvar_53[0][228] , \_zy_simnet_tvar_53[0][227] , 
	\_zy_simnet_tvar_53[0][226] , \_zy_simnet_tvar_53[0][225] , 
	\_zy_simnet_tvar_53[0][224] , \_zy_simnet_tvar_53[0][223] , 
	\_zy_simnet_tvar_53[0][222] , \_zy_simnet_tvar_53[0][221] , 
	\_zy_simnet_tvar_53[0][220] , \_zy_simnet_tvar_53[0][219] , 
	\_zy_simnet_tvar_53[0][218] , \_zy_simnet_tvar_53[0][217] , 
	\_zy_simnet_tvar_53[0][216] , \_zy_simnet_tvar_53[0][215] , 
	\_zy_simnet_tvar_53[0][214] , \_zy_simnet_tvar_53[0][213] , 
	\_zy_simnet_tvar_53[0][212] , \_zy_simnet_tvar_53[0][211] , 
	\_zy_simnet_tvar_53[0][210] , \_zy_simnet_tvar_53[0][209] , 
	\_zy_simnet_tvar_53[0][208] , \_zy_simnet_tvar_53[0][207] , 
	\_zy_simnet_tvar_53[0][206] , \_zy_simnet_tvar_53[0][205] , 
	\_zy_simnet_tvar_53[0][204] , \_zy_simnet_tvar_53[0][203] , 
	\_zy_simnet_tvar_53[0][202] , \_zy_simnet_tvar_53[0][201] , 
	\_zy_simnet_tvar_53[0][200] , \_zy_simnet_tvar_53[0][199] , 
	\_zy_simnet_tvar_53[0][198] , \_zy_simnet_tvar_53[0][197] , 
	\_zy_simnet_tvar_53[0][196] , \_zy_simnet_tvar_53[0][195] , 
	\_zy_simnet_tvar_53[0][194] , \_zy_simnet_tvar_53[0][193] , 
	\_zy_simnet_tvar_53[0][192] , \_zy_simnet_tvar_53[0][191] , 
	\_zy_simnet_tvar_53[0][190] , \_zy_simnet_tvar_53[0][189] , 
	\_zy_simnet_tvar_53[0][188] , \_zy_simnet_tvar_53[0][187] , 
	\_zy_simnet_tvar_53[0][186] , \_zy_simnet_tvar_53[0][185] , 
	\_zy_simnet_tvar_53[0][184] , \_zy_simnet_tvar_53[0][183] , 
	\_zy_simnet_tvar_53[0][182] , \_zy_simnet_tvar_53[0][181] , 
	\_zy_simnet_tvar_53[0][180] , \_zy_simnet_tvar_53[0][179] , 
	\_zy_simnet_tvar_53[0][178] , \_zy_simnet_tvar_53[0][177] , 
	\_zy_simnet_tvar_53[0][176] , \_zy_simnet_tvar_53[0][175] , 
	\_zy_simnet_tvar_53[0][174] , \_zy_simnet_tvar_53[0][173] , 
	\_zy_simnet_tvar_53[0][172] , \_zy_simnet_tvar_53[0][171] , 
	\_zy_simnet_tvar_53[0][170] , \_zy_simnet_tvar_53[0][169] , 
	\_zy_simnet_tvar_53[0][168] , \_zy_simnet_tvar_53[0][167] , 
	\_zy_simnet_tvar_53[0][166] , \_zy_simnet_tvar_53[0][165] , 
	\_zy_simnet_tvar_53[0][164] , \_zy_simnet_tvar_53[0][163] , 
	\_zy_simnet_tvar_53[0][162] , \_zy_simnet_tvar_53[0][161] , 
	\_zy_simnet_tvar_53[0][160] , \_zy_simnet_tvar_53[0][159] , 
	\_zy_simnet_tvar_53[0][158] , \_zy_simnet_tvar_53[0][157] , 
	\_zy_simnet_tvar_53[0][156] , \_zy_simnet_tvar_53[0][155] , 
	\_zy_simnet_tvar_53[0][154] , \_zy_simnet_tvar_53[0][153] , 
	\_zy_simnet_tvar_53[0][152] , \_zy_simnet_tvar_53[0][151] , 
	\_zy_simnet_tvar_53[0][150] , \_zy_simnet_tvar_53[0][149] , 
	\_zy_simnet_tvar_53[0][148] , \_zy_simnet_tvar_53[0][147] , 
	\_zy_simnet_tvar_53[0][146] , \_zy_simnet_tvar_53[0][145] , 
	\_zy_simnet_tvar_53[0][144] , \_zy_simnet_tvar_53[0][143] , 
	\_zy_simnet_tvar_53[0][142] , \_zy_simnet_tvar_53[0][141] , 
	\_zy_simnet_tvar_53[0][140] , \_zy_simnet_tvar_53[0][139] , 
	\_zy_simnet_tvar_53[0][138] , \_zy_simnet_tvar_53[0][137] , 
	\_zy_simnet_tvar_53[0][136] , \_zy_simnet_tvar_53[0][135] , 
	\_zy_simnet_tvar_53[0][134] , \_zy_simnet_tvar_53[0][133] , 
	\_zy_simnet_tvar_53[0][132] , \_zy_simnet_tvar_53[0][131] , 
	\_zy_simnet_tvar_53[0][130] , \_zy_simnet_tvar_53[0][129] , 
	\_zy_simnet_tvar_53[0][128] , \_zy_simnet_tvar_53[0][127] , 
	\_zy_simnet_tvar_53[0][126] , \_zy_simnet_tvar_53[0][125] , 
	\_zy_simnet_tvar_53[0][124] , \_zy_simnet_tvar_53[0][123] , 
	\_zy_simnet_tvar_53[0][122] , \_zy_simnet_tvar_53[0][121] , 
	\_zy_simnet_tvar_53[0][120] , \_zy_simnet_tvar_53[0][119] , 
	\_zy_simnet_tvar_53[0][118] , \_zy_simnet_tvar_53[0][117] , 
	\_zy_simnet_tvar_53[0][116] , \_zy_simnet_tvar_53[0][115] , 
	\_zy_simnet_tvar_53[0][114] , \_zy_simnet_tvar_53[0][113] , 
	\_zy_simnet_tvar_53[0][112] , \_zy_simnet_tvar_53[0][111] , 
	\_zy_simnet_tvar_53[0][110] , \_zy_simnet_tvar_53[0][109] , 
	\_zy_simnet_tvar_53[0][108] , \_zy_simnet_tvar_53[0][107] , 
	\_zy_simnet_tvar_53[0][106] , \_zy_simnet_tvar_53[0][105] , 
	\_zy_simnet_tvar_53[0][104] , \_zy_simnet_tvar_53[0][103] , 
	\_zy_simnet_tvar_53[0][102] , \_zy_simnet_tvar_53[0][101] , 
	\_zy_simnet_tvar_53[0][100] , \_zy_simnet_tvar_53[0][99] , 
	\_zy_simnet_tvar_53[0][98] , \_zy_simnet_tvar_53[0][97] , 
	\_zy_simnet_tvar_53[0][96] , \_zy_simnet_tvar_53[0][95] , 
	\_zy_simnet_tvar_53[0][94] , \_zy_simnet_tvar_53[0][93] , 
	\_zy_simnet_tvar_53[0][92] , \_zy_simnet_tvar_53[0][91] , 
	\_zy_simnet_tvar_53[0][90] , \_zy_simnet_tvar_53[0][89] , 
	\_zy_simnet_tvar_53[0][88] , \_zy_simnet_tvar_53[0][87] , 
	\_zy_simnet_tvar_53[0][86] , \_zy_simnet_tvar_53[0][85] , 
	\_zy_simnet_tvar_53[0][84] , \_zy_simnet_tvar_53[0][83] , 
	\_zy_simnet_tvar_53[0][82] , \_zy_simnet_tvar_53[0][81] , 
	\_zy_simnet_tvar_53[0][80] , \_zy_simnet_tvar_53[0][79] , 
	\_zy_simnet_tvar_53[0][78] , \_zy_simnet_tvar_53[0][77] , 
	\_zy_simnet_tvar_53[0][76] , \_zy_simnet_tvar_53[0][75] , 
	\_zy_simnet_tvar_53[0][74] , \_zy_simnet_tvar_53[0][73] , 
	\_zy_simnet_tvar_53[0][72] , \_zy_simnet_tvar_53[0][71] , 
	\_zy_simnet_tvar_53[0][70] , \_zy_simnet_tvar_53[0][69] , 
	\_zy_simnet_tvar_53[0][68] , \_zy_simnet_tvar_53[0][67] , 
	\_zy_simnet_tvar_53[0][66] , \_zy_simnet_tvar_53[0][65] , 
	\_zy_simnet_tvar_53[0][64] , \_zy_simnet_tvar_53[0][63] , 
	\_zy_simnet_tvar_53[0][62] , \_zy_simnet_tvar_53[0][61] , 
	\_zy_simnet_tvar_53[0][60] , \_zy_simnet_tvar_53[0][59] , 
	\_zy_simnet_tvar_53[0][58] , \_zy_simnet_tvar_53[0][57] , 
	\_zy_simnet_tvar_53[0][56] , \_zy_simnet_tvar_53[0][55] , 
	\_zy_simnet_tvar_53[0][54] , \_zy_simnet_tvar_53[0][53] , 
	\_zy_simnet_tvar_53[0][52] , \_zy_simnet_tvar_53[0][51] , 
	\_zy_simnet_tvar_53[0][50] , \_zy_simnet_tvar_53[0][49] , 
	\_zy_simnet_tvar_53[0][48] , \_zy_simnet_tvar_53[0][47] , 
	\_zy_simnet_tvar_53[0][46] , \_zy_simnet_tvar_53[0][45] , 
	\_zy_simnet_tvar_53[0][44] , \_zy_simnet_tvar_53[0][43] , 
	\_zy_simnet_tvar_53[0][42] , \_zy_simnet_tvar_53[0][41] , 
	\_zy_simnet_tvar_53[0][40] , \_zy_simnet_tvar_53[0][39] , 
	\_zy_simnet_tvar_53[0][38] , \_zy_simnet_tvar_53[0][37] , 
	\_zy_simnet_tvar_53[0][36] , \_zy_simnet_tvar_53[0][35] , 
	\_zy_simnet_tvar_53[0][34] , \_zy_simnet_tvar_53[0][33] , 
	\_zy_simnet_tvar_53[0][32] , \_zy_simnet_tvar_53[0][31] , 
	\_zy_simnet_tvar_53[0][30] , \_zy_simnet_tvar_53[0][29] , 
	\_zy_simnet_tvar_53[0][28] , \_zy_simnet_tvar_53[0][27] , 
	\_zy_simnet_tvar_53[0][26] , \_zy_simnet_tvar_53[0][25] , 
	\_zy_simnet_tvar_53[0][24] , \_zy_simnet_tvar_53[0][23] , 
	\_zy_simnet_tvar_53[0][22] , \_zy_simnet_tvar_53[0][21] , 
	\_zy_simnet_tvar_53[0][20] , \_zy_simnet_tvar_53[0][19] , 
	\_zy_simnet_tvar_53[0][18] , \_zy_simnet_tvar_53[0][17] , 
	\_zy_simnet_tvar_53[0][16] , \_zy_simnet_tvar_53[0][15] , 
	\_zy_simnet_tvar_53[0][14] , \_zy_simnet_tvar_53[0][13] , 
	\_zy_simnet_tvar_53[0][12] , \_zy_simnet_tvar_53[0][11] , 
	\_zy_simnet_tvar_53[0][10] , \_zy_simnet_tvar_53[0][9] , 
	\_zy_simnet_tvar_53[0][8] , \_zy_simnet_tvar_53[0][7] , 
	\_zy_simnet_tvar_53[0][6] , \_zy_simnet_tvar_53[0][5] , 
	\_zy_simnet_tvar_53[0][4] , \_zy_simnet_tvar_53[0][3] , 
	\_zy_simnet_tvar_53[0][2] , \_zy_simnet_tvar_53[0][1] , 
	\_zy_simnet_tvar_53[0][0] });
ixc_assign_2176 _zz_strnp_29 ( { \_zy_simnet_tvar_20[7][271] , 
	\_zy_simnet_tvar_20[7][270] , \_zy_simnet_tvar_20[7][269] , 
	\_zy_simnet_tvar_20[7][268] , \_zy_simnet_tvar_20[7][267] , 
	\_zy_simnet_tvar_20[7][266] , \_zy_simnet_tvar_20[7][265] , 
	\_zy_simnet_tvar_20[7][264] , \_zy_simnet_tvar_20[7][263] , 
	\_zy_simnet_tvar_20[7][262] , \_zy_simnet_tvar_20[7][261] , 
	\_zy_simnet_tvar_20[7][260] , \_zy_simnet_tvar_20[7][259] , 
	\_zy_simnet_tvar_20[7][258] , \_zy_simnet_tvar_20[7][257] , 
	\_zy_simnet_tvar_20[7][256] , \_zy_simnet_tvar_20[7][255] , 
	\_zy_simnet_tvar_20[7][254] , \_zy_simnet_tvar_20[7][253] , 
	\_zy_simnet_tvar_20[7][252] , \_zy_simnet_tvar_20[7][251] , 
	\_zy_simnet_tvar_20[7][250] , \_zy_simnet_tvar_20[7][249] , 
	\_zy_simnet_tvar_20[7][248] , \_zy_simnet_tvar_20[7][247] , 
	\_zy_simnet_tvar_20[7][246] , \_zy_simnet_tvar_20[7][245] , 
	\_zy_simnet_tvar_20[7][244] , \_zy_simnet_tvar_20[7][243] , 
	\_zy_simnet_tvar_20[7][242] , \_zy_simnet_tvar_20[7][241] , 
	\_zy_simnet_tvar_20[7][240] , \_zy_simnet_tvar_20[7][239] , 
	\_zy_simnet_tvar_20[7][238] , \_zy_simnet_tvar_20[7][237] , 
	\_zy_simnet_tvar_20[7][236] , \_zy_simnet_tvar_20[7][235] , 
	\_zy_simnet_tvar_20[7][234] , \_zy_simnet_tvar_20[7][233] , 
	\_zy_simnet_tvar_20[7][232] , \_zy_simnet_tvar_20[7][231] , 
	\_zy_simnet_tvar_20[7][230] , \_zy_simnet_tvar_20[7][229] , 
	\_zy_simnet_tvar_20[7][228] , \_zy_simnet_tvar_20[7][227] , 
	\_zy_simnet_tvar_20[7][226] , \_zy_simnet_tvar_20[7][225] , 
	\_zy_simnet_tvar_20[7][224] , \_zy_simnet_tvar_20[7][223] , 
	\_zy_simnet_tvar_20[7][222] , \_zy_simnet_tvar_20[7][221] , 
	\_zy_simnet_tvar_20[7][220] , \_zy_simnet_tvar_20[7][219] , 
	\_zy_simnet_tvar_20[7][218] , \_zy_simnet_tvar_20[7][217] , 
	\_zy_simnet_tvar_20[7][216] , \_zy_simnet_tvar_20[7][215] , 
	\_zy_simnet_tvar_20[7][214] , \_zy_simnet_tvar_20[7][213] , 
	\_zy_simnet_tvar_20[7][212] , \_zy_simnet_tvar_20[7][211] , 
	\_zy_simnet_tvar_20[7][210] , \_zy_simnet_tvar_20[7][209] , 
	\_zy_simnet_tvar_20[7][208] , \_zy_simnet_tvar_20[7][207] , 
	\_zy_simnet_tvar_20[7][206] , \_zy_simnet_tvar_20[7][205] , 
	\_zy_simnet_tvar_20[7][204] , \_zy_simnet_tvar_20[7][203] , 
	\_zy_simnet_tvar_20[7][202] , \_zy_simnet_tvar_20[7][201] , 
	\_zy_simnet_tvar_20[7][200] , \_zy_simnet_tvar_20[7][199] , 
	\_zy_simnet_tvar_20[7][198] , \_zy_simnet_tvar_20[7][197] , 
	\_zy_simnet_tvar_20[7][196] , \_zy_simnet_tvar_20[7][195] , 
	\_zy_simnet_tvar_20[7][194] , \_zy_simnet_tvar_20[7][193] , 
	\_zy_simnet_tvar_20[7][192] , \_zy_simnet_tvar_20[7][191] , 
	\_zy_simnet_tvar_20[7][190] , \_zy_simnet_tvar_20[7][189] , 
	\_zy_simnet_tvar_20[7][188] , \_zy_simnet_tvar_20[7][187] , 
	\_zy_simnet_tvar_20[7][186] , \_zy_simnet_tvar_20[7][185] , 
	\_zy_simnet_tvar_20[7][184] , \_zy_simnet_tvar_20[7][183] , 
	\_zy_simnet_tvar_20[7][182] , \_zy_simnet_tvar_20[7][181] , 
	\_zy_simnet_tvar_20[7][180] , \_zy_simnet_tvar_20[7][179] , 
	\_zy_simnet_tvar_20[7][178] , \_zy_simnet_tvar_20[7][177] , 
	\_zy_simnet_tvar_20[7][176] , \_zy_simnet_tvar_20[7][175] , 
	\_zy_simnet_tvar_20[7][174] , \_zy_simnet_tvar_20[7][173] , 
	\_zy_simnet_tvar_20[7][172] , \_zy_simnet_tvar_20[7][171] , 
	\_zy_simnet_tvar_20[7][170] , \_zy_simnet_tvar_20[7][169] , 
	\_zy_simnet_tvar_20[7][168] , \_zy_simnet_tvar_20[7][167] , 
	\_zy_simnet_tvar_20[7][166] , \_zy_simnet_tvar_20[7][165] , 
	\_zy_simnet_tvar_20[7][164] , \_zy_simnet_tvar_20[7][163] , 
	\_zy_simnet_tvar_20[7][162] , \_zy_simnet_tvar_20[7][161] , 
	\_zy_simnet_tvar_20[7][160] , \_zy_simnet_tvar_20[7][159] , 
	\_zy_simnet_tvar_20[7][158] , \_zy_simnet_tvar_20[7][157] , 
	\_zy_simnet_tvar_20[7][156] , \_zy_simnet_tvar_20[7][155] , 
	\_zy_simnet_tvar_20[7][154] , \_zy_simnet_tvar_20[7][153] , 
	\_zy_simnet_tvar_20[7][152] , \_zy_simnet_tvar_20[7][151] , 
	\_zy_simnet_tvar_20[7][150] , \_zy_simnet_tvar_20[7][149] , 
	\_zy_simnet_tvar_20[7][148] , \_zy_simnet_tvar_20[7][147] , 
	\_zy_simnet_tvar_20[7][146] , \_zy_simnet_tvar_20[7][145] , 
	\_zy_simnet_tvar_20[7][144] , \_zy_simnet_tvar_20[7][143] , 
	\_zy_simnet_tvar_20[7][142] , \_zy_simnet_tvar_20[7][141] , 
	\_zy_simnet_tvar_20[7][140] , \_zy_simnet_tvar_20[7][139] , 
	\_zy_simnet_tvar_20[7][138] , \_zy_simnet_tvar_20[7][137] , 
	\_zy_simnet_tvar_20[7][136] , \_zy_simnet_tvar_20[7][135] , 
	\_zy_simnet_tvar_20[7][134] , \_zy_simnet_tvar_20[7][133] , 
	\_zy_simnet_tvar_20[7][132] , \_zy_simnet_tvar_20[7][131] , 
	\_zy_simnet_tvar_20[7][130] , \_zy_simnet_tvar_20[7][129] , 
	\_zy_simnet_tvar_20[7][128] , \_zy_simnet_tvar_20[7][127] , 
	\_zy_simnet_tvar_20[7][126] , \_zy_simnet_tvar_20[7][125] , 
	\_zy_simnet_tvar_20[7][124] , \_zy_simnet_tvar_20[7][123] , 
	\_zy_simnet_tvar_20[7][122] , \_zy_simnet_tvar_20[7][121] , 
	\_zy_simnet_tvar_20[7][120] , \_zy_simnet_tvar_20[7][119] , 
	\_zy_simnet_tvar_20[7][118] , \_zy_simnet_tvar_20[7][117] , 
	\_zy_simnet_tvar_20[7][116] , \_zy_simnet_tvar_20[7][115] , 
	\_zy_simnet_tvar_20[7][114] , \_zy_simnet_tvar_20[7][113] , 
	\_zy_simnet_tvar_20[7][112] , \_zy_simnet_tvar_20[7][111] , 
	\_zy_simnet_tvar_20[7][110] , \_zy_simnet_tvar_20[7][109] , 
	\_zy_simnet_tvar_20[7][108] , \_zy_simnet_tvar_20[7][107] , 
	\_zy_simnet_tvar_20[7][106] , \_zy_simnet_tvar_20[7][105] , 
	\_zy_simnet_tvar_20[7][104] , \_zy_simnet_tvar_20[7][103] , 
	\_zy_simnet_tvar_20[7][102] , \_zy_simnet_tvar_20[7][101] , 
	\_zy_simnet_tvar_20[7][100] , \_zy_simnet_tvar_20[7][99] , 
	\_zy_simnet_tvar_20[7][98] , \_zy_simnet_tvar_20[7][97] , 
	\_zy_simnet_tvar_20[7][96] , \_zy_simnet_tvar_20[7][95] , 
	\_zy_simnet_tvar_20[7][94] , \_zy_simnet_tvar_20[7][93] , 
	\_zy_simnet_tvar_20[7][92] , \_zy_simnet_tvar_20[7][91] , 
	\_zy_simnet_tvar_20[7][90] , \_zy_simnet_tvar_20[7][89] , 
	\_zy_simnet_tvar_20[7][88] , \_zy_simnet_tvar_20[7][87] , 
	\_zy_simnet_tvar_20[7][86] , \_zy_simnet_tvar_20[7][85] , 
	\_zy_simnet_tvar_20[7][84] , \_zy_simnet_tvar_20[7][83] , 
	\_zy_simnet_tvar_20[7][82] , \_zy_simnet_tvar_20[7][81] , 
	\_zy_simnet_tvar_20[7][80] , \_zy_simnet_tvar_20[7][79] , 
	\_zy_simnet_tvar_20[7][78] , \_zy_simnet_tvar_20[7][77] , 
	\_zy_simnet_tvar_20[7][76] , \_zy_simnet_tvar_20[7][75] , 
	\_zy_simnet_tvar_20[7][74] , \_zy_simnet_tvar_20[7][73] , 
	\_zy_simnet_tvar_20[7][72] , \_zy_simnet_tvar_20[7][71] , 
	\_zy_simnet_tvar_20[7][70] , \_zy_simnet_tvar_20[7][69] , 
	\_zy_simnet_tvar_20[7][68] , \_zy_simnet_tvar_20[7][67] , 
	\_zy_simnet_tvar_20[7][66] , \_zy_simnet_tvar_20[7][65] , 
	\_zy_simnet_tvar_20[7][64] , \_zy_simnet_tvar_20[7][63] , 
	\_zy_simnet_tvar_20[7][62] , \_zy_simnet_tvar_20[7][61] , 
	\_zy_simnet_tvar_20[7][60] , \_zy_simnet_tvar_20[7][59] , 
	\_zy_simnet_tvar_20[7][58] , \_zy_simnet_tvar_20[7][57] , 
	\_zy_simnet_tvar_20[7][56] , \_zy_simnet_tvar_20[7][55] , 
	\_zy_simnet_tvar_20[7][54] , \_zy_simnet_tvar_20[7][53] , 
	\_zy_simnet_tvar_20[7][52] , \_zy_simnet_tvar_20[7][51] , 
	\_zy_simnet_tvar_20[7][50] , \_zy_simnet_tvar_20[7][49] , 
	\_zy_simnet_tvar_20[7][48] , \_zy_simnet_tvar_20[7][47] , 
	\_zy_simnet_tvar_20[7][46] , \_zy_simnet_tvar_20[7][45] , 
	\_zy_simnet_tvar_20[7][44] , \_zy_simnet_tvar_20[7][43] , 
	\_zy_simnet_tvar_20[7][42] , \_zy_simnet_tvar_20[7][41] , 
	\_zy_simnet_tvar_20[7][40] , \_zy_simnet_tvar_20[7][39] , 
	\_zy_simnet_tvar_20[7][38] , \_zy_simnet_tvar_20[7][37] , 
	\_zy_simnet_tvar_20[7][36] , \_zy_simnet_tvar_20[7][35] , 
	\_zy_simnet_tvar_20[7][34] , \_zy_simnet_tvar_20[7][33] , 
	\_zy_simnet_tvar_20[7][32] , \_zy_simnet_tvar_20[7][31] , 
	\_zy_simnet_tvar_20[7][30] , \_zy_simnet_tvar_20[7][29] , 
	\_zy_simnet_tvar_20[7][28] , \_zy_simnet_tvar_20[7][27] , 
	\_zy_simnet_tvar_20[7][26] , \_zy_simnet_tvar_20[7][25] , 
	\_zy_simnet_tvar_20[7][24] , \_zy_simnet_tvar_20[7][23] , 
	\_zy_simnet_tvar_20[7][22] , \_zy_simnet_tvar_20[7][21] , 
	\_zy_simnet_tvar_20[7][20] , \_zy_simnet_tvar_20[7][19] , 
	\_zy_simnet_tvar_20[7][18] , \_zy_simnet_tvar_20[7][17] , 
	\_zy_simnet_tvar_20[7][16] , \_zy_simnet_tvar_20[7][15] , 
	\_zy_simnet_tvar_20[7][14] , \_zy_simnet_tvar_20[7][13] , 
	\_zy_simnet_tvar_20[7][12] , \_zy_simnet_tvar_20[7][11] , 
	\_zy_simnet_tvar_20[7][10] , \_zy_simnet_tvar_20[7][9] , 
	\_zy_simnet_tvar_20[7][8] , \_zy_simnet_tvar_20[7][7] , 
	\_zy_simnet_tvar_20[7][6] , \_zy_simnet_tvar_20[7][5] , 
	\_zy_simnet_tvar_20[7][4] , \_zy_simnet_tvar_20[7][3] , 
	\_zy_simnet_tvar_20[7][2] , \_zy_simnet_tvar_20[7][1] , 
	\_zy_simnet_tvar_20[7][0] , \_zy_simnet_tvar_20[6][271] , 
	\_zy_simnet_tvar_20[6][270] , \_zy_simnet_tvar_20[6][269] , 
	\_zy_simnet_tvar_20[6][268] , \_zy_simnet_tvar_20[6][267] , 
	\_zy_simnet_tvar_20[6][266] , \_zy_simnet_tvar_20[6][265] , 
	\_zy_simnet_tvar_20[6][264] , \_zy_simnet_tvar_20[6][263] , 
	\_zy_simnet_tvar_20[6][262] , \_zy_simnet_tvar_20[6][261] , 
	\_zy_simnet_tvar_20[6][260] , \_zy_simnet_tvar_20[6][259] , 
	\_zy_simnet_tvar_20[6][258] , \_zy_simnet_tvar_20[6][257] , 
	\_zy_simnet_tvar_20[6][256] , \_zy_simnet_tvar_20[6][255] , 
	\_zy_simnet_tvar_20[6][254] , \_zy_simnet_tvar_20[6][253] , 
	\_zy_simnet_tvar_20[6][252] , \_zy_simnet_tvar_20[6][251] , 
	\_zy_simnet_tvar_20[6][250] , \_zy_simnet_tvar_20[6][249] , 
	\_zy_simnet_tvar_20[6][248] , \_zy_simnet_tvar_20[6][247] , 
	\_zy_simnet_tvar_20[6][246] , \_zy_simnet_tvar_20[6][245] , 
	\_zy_simnet_tvar_20[6][244] , \_zy_simnet_tvar_20[6][243] , 
	\_zy_simnet_tvar_20[6][242] , \_zy_simnet_tvar_20[6][241] , 
	\_zy_simnet_tvar_20[6][240] , \_zy_simnet_tvar_20[6][239] , 
	\_zy_simnet_tvar_20[6][238] , \_zy_simnet_tvar_20[6][237] , 
	\_zy_simnet_tvar_20[6][236] , \_zy_simnet_tvar_20[6][235] , 
	\_zy_simnet_tvar_20[6][234] , \_zy_simnet_tvar_20[6][233] , 
	\_zy_simnet_tvar_20[6][232] , \_zy_simnet_tvar_20[6][231] , 
	\_zy_simnet_tvar_20[6][230] , \_zy_simnet_tvar_20[6][229] , 
	\_zy_simnet_tvar_20[6][228] , \_zy_simnet_tvar_20[6][227] , 
	\_zy_simnet_tvar_20[6][226] , \_zy_simnet_tvar_20[6][225] , 
	\_zy_simnet_tvar_20[6][224] , \_zy_simnet_tvar_20[6][223] , 
	\_zy_simnet_tvar_20[6][222] , \_zy_simnet_tvar_20[6][221] , 
	\_zy_simnet_tvar_20[6][220] , \_zy_simnet_tvar_20[6][219] , 
	\_zy_simnet_tvar_20[6][218] , \_zy_simnet_tvar_20[6][217] , 
	\_zy_simnet_tvar_20[6][216] , \_zy_simnet_tvar_20[6][215] , 
	\_zy_simnet_tvar_20[6][214] , \_zy_simnet_tvar_20[6][213] , 
	\_zy_simnet_tvar_20[6][212] , \_zy_simnet_tvar_20[6][211] , 
	\_zy_simnet_tvar_20[6][210] , \_zy_simnet_tvar_20[6][209] , 
	\_zy_simnet_tvar_20[6][208] , \_zy_simnet_tvar_20[6][207] , 
	\_zy_simnet_tvar_20[6][206] , \_zy_simnet_tvar_20[6][205] , 
	\_zy_simnet_tvar_20[6][204] , \_zy_simnet_tvar_20[6][203] , 
	\_zy_simnet_tvar_20[6][202] , \_zy_simnet_tvar_20[6][201] , 
	\_zy_simnet_tvar_20[6][200] , \_zy_simnet_tvar_20[6][199] , 
	\_zy_simnet_tvar_20[6][198] , \_zy_simnet_tvar_20[6][197] , 
	\_zy_simnet_tvar_20[6][196] , \_zy_simnet_tvar_20[6][195] , 
	\_zy_simnet_tvar_20[6][194] , \_zy_simnet_tvar_20[6][193] , 
	\_zy_simnet_tvar_20[6][192] , \_zy_simnet_tvar_20[6][191] , 
	\_zy_simnet_tvar_20[6][190] , \_zy_simnet_tvar_20[6][189] , 
	\_zy_simnet_tvar_20[6][188] , \_zy_simnet_tvar_20[6][187] , 
	\_zy_simnet_tvar_20[6][186] , \_zy_simnet_tvar_20[6][185] , 
	\_zy_simnet_tvar_20[6][184] , \_zy_simnet_tvar_20[6][183] , 
	\_zy_simnet_tvar_20[6][182] , \_zy_simnet_tvar_20[6][181] , 
	\_zy_simnet_tvar_20[6][180] , \_zy_simnet_tvar_20[6][179] , 
	\_zy_simnet_tvar_20[6][178] , \_zy_simnet_tvar_20[6][177] , 
	\_zy_simnet_tvar_20[6][176] , \_zy_simnet_tvar_20[6][175] , 
	\_zy_simnet_tvar_20[6][174] , \_zy_simnet_tvar_20[6][173] , 
	\_zy_simnet_tvar_20[6][172] , \_zy_simnet_tvar_20[6][171] , 
	\_zy_simnet_tvar_20[6][170] , \_zy_simnet_tvar_20[6][169] , 
	\_zy_simnet_tvar_20[6][168] , \_zy_simnet_tvar_20[6][167] , 
	\_zy_simnet_tvar_20[6][166] , \_zy_simnet_tvar_20[6][165] , 
	\_zy_simnet_tvar_20[6][164] , \_zy_simnet_tvar_20[6][163] , 
	\_zy_simnet_tvar_20[6][162] , \_zy_simnet_tvar_20[6][161] , 
	\_zy_simnet_tvar_20[6][160] , \_zy_simnet_tvar_20[6][159] , 
	\_zy_simnet_tvar_20[6][158] , \_zy_simnet_tvar_20[6][157] , 
	\_zy_simnet_tvar_20[6][156] , \_zy_simnet_tvar_20[6][155] , 
	\_zy_simnet_tvar_20[6][154] , \_zy_simnet_tvar_20[6][153] , 
	\_zy_simnet_tvar_20[6][152] , \_zy_simnet_tvar_20[6][151] , 
	\_zy_simnet_tvar_20[6][150] , \_zy_simnet_tvar_20[6][149] , 
	\_zy_simnet_tvar_20[6][148] , \_zy_simnet_tvar_20[6][147] , 
	\_zy_simnet_tvar_20[6][146] , \_zy_simnet_tvar_20[6][145] , 
	\_zy_simnet_tvar_20[6][144] , \_zy_simnet_tvar_20[6][143] , 
	\_zy_simnet_tvar_20[6][142] , \_zy_simnet_tvar_20[6][141] , 
	\_zy_simnet_tvar_20[6][140] , \_zy_simnet_tvar_20[6][139] , 
	\_zy_simnet_tvar_20[6][138] , \_zy_simnet_tvar_20[6][137] , 
	\_zy_simnet_tvar_20[6][136] , \_zy_simnet_tvar_20[6][135] , 
	\_zy_simnet_tvar_20[6][134] , \_zy_simnet_tvar_20[6][133] , 
	\_zy_simnet_tvar_20[6][132] , \_zy_simnet_tvar_20[6][131] , 
	\_zy_simnet_tvar_20[6][130] , \_zy_simnet_tvar_20[6][129] , 
	\_zy_simnet_tvar_20[6][128] , \_zy_simnet_tvar_20[6][127] , 
	\_zy_simnet_tvar_20[6][126] , \_zy_simnet_tvar_20[6][125] , 
	\_zy_simnet_tvar_20[6][124] , \_zy_simnet_tvar_20[6][123] , 
	\_zy_simnet_tvar_20[6][122] , \_zy_simnet_tvar_20[6][121] , 
	\_zy_simnet_tvar_20[6][120] , \_zy_simnet_tvar_20[6][119] , 
	\_zy_simnet_tvar_20[6][118] , \_zy_simnet_tvar_20[6][117] , 
	\_zy_simnet_tvar_20[6][116] , \_zy_simnet_tvar_20[6][115] , 
	\_zy_simnet_tvar_20[6][114] , \_zy_simnet_tvar_20[6][113] , 
	\_zy_simnet_tvar_20[6][112] , \_zy_simnet_tvar_20[6][111] , 
	\_zy_simnet_tvar_20[6][110] , \_zy_simnet_tvar_20[6][109] , 
	\_zy_simnet_tvar_20[6][108] , \_zy_simnet_tvar_20[6][107] , 
	\_zy_simnet_tvar_20[6][106] , \_zy_simnet_tvar_20[6][105] , 
	\_zy_simnet_tvar_20[6][104] , \_zy_simnet_tvar_20[6][103] , 
	\_zy_simnet_tvar_20[6][102] , \_zy_simnet_tvar_20[6][101] , 
	\_zy_simnet_tvar_20[6][100] , \_zy_simnet_tvar_20[6][99] , 
	\_zy_simnet_tvar_20[6][98] , \_zy_simnet_tvar_20[6][97] , 
	\_zy_simnet_tvar_20[6][96] , \_zy_simnet_tvar_20[6][95] , 
	\_zy_simnet_tvar_20[6][94] , \_zy_simnet_tvar_20[6][93] , 
	\_zy_simnet_tvar_20[6][92] , \_zy_simnet_tvar_20[6][91] , 
	\_zy_simnet_tvar_20[6][90] , \_zy_simnet_tvar_20[6][89] , 
	\_zy_simnet_tvar_20[6][88] , \_zy_simnet_tvar_20[6][87] , 
	\_zy_simnet_tvar_20[6][86] , \_zy_simnet_tvar_20[6][85] , 
	\_zy_simnet_tvar_20[6][84] , \_zy_simnet_tvar_20[6][83] , 
	\_zy_simnet_tvar_20[6][82] , \_zy_simnet_tvar_20[6][81] , 
	\_zy_simnet_tvar_20[6][80] , \_zy_simnet_tvar_20[6][79] , 
	\_zy_simnet_tvar_20[6][78] , \_zy_simnet_tvar_20[6][77] , 
	\_zy_simnet_tvar_20[6][76] , \_zy_simnet_tvar_20[6][75] , 
	\_zy_simnet_tvar_20[6][74] , \_zy_simnet_tvar_20[6][73] , 
	\_zy_simnet_tvar_20[6][72] , \_zy_simnet_tvar_20[6][71] , 
	\_zy_simnet_tvar_20[6][70] , \_zy_simnet_tvar_20[6][69] , 
	\_zy_simnet_tvar_20[6][68] , \_zy_simnet_tvar_20[6][67] , 
	\_zy_simnet_tvar_20[6][66] , \_zy_simnet_tvar_20[6][65] , 
	\_zy_simnet_tvar_20[6][64] , \_zy_simnet_tvar_20[6][63] , 
	\_zy_simnet_tvar_20[6][62] , \_zy_simnet_tvar_20[6][61] , 
	\_zy_simnet_tvar_20[6][60] , \_zy_simnet_tvar_20[6][59] , 
	\_zy_simnet_tvar_20[6][58] , \_zy_simnet_tvar_20[6][57] , 
	\_zy_simnet_tvar_20[6][56] , \_zy_simnet_tvar_20[6][55] , 
	\_zy_simnet_tvar_20[6][54] , \_zy_simnet_tvar_20[6][53] , 
	\_zy_simnet_tvar_20[6][52] , \_zy_simnet_tvar_20[6][51] , 
	\_zy_simnet_tvar_20[6][50] , \_zy_simnet_tvar_20[6][49] , 
	\_zy_simnet_tvar_20[6][48] , \_zy_simnet_tvar_20[6][47] , 
	\_zy_simnet_tvar_20[6][46] , \_zy_simnet_tvar_20[6][45] , 
	\_zy_simnet_tvar_20[6][44] , \_zy_simnet_tvar_20[6][43] , 
	\_zy_simnet_tvar_20[6][42] , \_zy_simnet_tvar_20[6][41] , 
	\_zy_simnet_tvar_20[6][40] , \_zy_simnet_tvar_20[6][39] , 
	\_zy_simnet_tvar_20[6][38] , \_zy_simnet_tvar_20[6][37] , 
	\_zy_simnet_tvar_20[6][36] , \_zy_simnet_tvar_20[6][35] , 
	\_zy_simnet_tvar_20[6][34] , \_zy_simnet_tvar_20[6][33] , 
	\_zy_simnet_tvar_20[6][32] , \_zy_simnet_tvar_20[6][31] , 
	\_zy_simnet_tvar_20[6][30] , \_zy_simnet_tvar_20[6][29] , 
	\_zy_simnet_tvar_20[6][28] , \_zy_simnet_tvar_20[6][27] , 
	\_zy_simnet_tvar_20[6][26] , \_zy_simnet_tvar_20[6][25] , 
	\_zy_simnet_tvar_20[6][24] , \_zy_simnet_tvar_20[6][23] , 
	\_zy_simnet_tvar_20[6][22] , \_zy_simnet_tvar_20[6][21] , 
	\_zy_simnet_tvar_20[6][20] , \_zy_simnet_tvar_20[6][19] , 
	\_zy_simnet_tvar_20[6][18] , \_zy_simnet_tvar_20[6][17] , 
	\_zy_simnet_tvar_20[6][16] , \_zy_simnet_tvar_20[6][15] , 
	\_zy_simnet_tvar_20[6][14] , \_zy_simnet_tvar_20[6][13] , 
	\_zy_simnet_tvar_20[6][12] , \_zy_simnet_tvar_20[6][11] , 
	\_zy_simnet_tvar_20[6][10] , \_zy_simnet_tvar_20[6][9] , 
	\_zy_simnet_tvar_20[6][8] , \_zy_simnet_tvar_20[6][7] , 
	\_zy_simnet_tvar_20[6][6] , \_zy_simnet_tvar_20[6][5] , 
	\_zy_simnet_tvar_20[6][4] , \_zy_simnet_tvar_20[6][3] , 
	\_zy_simnet_tvar_20[6][2] , \_zy_simnet_tvar_20[6][1] , 
	\_zy_simnet_tvar_20[6][0] , \_zy_simnet_tvar_20[5][271] , 
	\_zy_simnet_tvar_20[5][270] , \_zy_simnet_tvar_20[5][269] , 
	\_zy_simnet_tvar_20[5][268] , \_zy_simnet_tvar_20[5][267] , 
	\_zy_simnet_tvar_20[5][266] , \_zy_simnet_tvar_20[5][265] , 
	\_zy_simnet_tvar_20[5][264] , \_zy_simnet_tvar_20[5][263] , 
	\_zy_simnet_tvar_20[5][262] , \_zy_simnet_tvar_20[5][261] , 
	\_zy_simnet_tvar_20[5][260] , \_zy_simnet_tvar_20[5][259] , 
	\_zy_simnet_tvar_20[5][258] , \_zy_simnet_tvar_20[5][257] , 
	\_zy_simnet_tvar_20[5][256] , \_zy_simnet_tvar_20[5][255] , 
	\_zy_simnet_tvar_20[5][254] , \_zy_simnet_tvar_20[5][253] , 
	\_zy_simnet_tvar_20[5][252] , \_zy_simnet_tvar_20[5][251] , 
	\_zy_simnet_tvar_20[5][250] , \_zy_simnet_tvar_20[5][249] , 
	\_zy_simnet_tvar_20[5][248] , \_zy_simnet_tvar_20[5][247] , 
	\_zy_simnet_tvar_20[5][246] , \_zy_simnet_tvar_20[5][245] , 
	\_zy_simnet_tvar_20[5][244] , \_zy_simnet_tvar_20[5][243] , 
	\_zy_simnet_tvar_20[5][242] , \_zy_simnet_tvar_20[5][241] , 
	\_zy_simnet_tvar_20[5][240] , \_zy_simnet_tvar_20[5][239] , 
	\_zy_simnet_tvar_20[5][238] , \_zy_simnet_tvar_20[5][237] , 
	\_zy_simnet_tvar_20[5][236] , \_zy_simnet_tvar_20[5][235] , 
	\_zy_simnet_tvar_20[5][234] , \_zy_simnet_tvar_20[5][233] , 
	\_zy_simnet_tvar_20[5][232] , \_zy_simnet_tvar_20[5][231] , 
	\_zy_simnet_tvar_20[5][230] , \_zy_simnet_tvar_20[5][229] , 
	\_zy_simnet_tvar_20[5][228] , \_zy_simnet_tvar_20[5][227] , 
	\_zy_simnet_tvar_20[5][226] , \_zy_simnet_tvar_20[5][225] , 
	\_zy_simnet_tvar_20[5][224] , \_zy_simnet_tvar_20[5][223] , 
	\_zy_simnet_tvar_20[5][222] , \_zy_simnet_tvar_20[5][221] , 
	\_zy_simnet_tvar_20[5][220] , \_zy_simnet_tvar_20[5][219] , 
	\_zy_simnet_tvar_20[5][218] , \_zy_simnet_tvar_20[5][217] , 
	\_zy_simnet_tvar_20[5][216] , \_zy_simnet_tvar_20[5][215] , 
	\_zy_simnet_tvar_20[5][214] , \_zy_simnet_tvar_20[5][213] , 
	\_zy_simnet_tvar_20[5][212] , \_zy_simnet_tvar_20[5][211] , 
	\_zy_simnet_tvar_20[5][210] , \_zy_simnet_tvar_20[5][209] , 
	\_zy_simnet_tvar_20[5][208] , \_zy_simnet_tvar_20[5][207] , 
	\_zy_simnet_tvar_20[5][206] , \_zy_simnet_tvar_20[5][205] , 
	\_zy_simnet_tvar_20[5][204] , \_zy_simnet_tvar_20[5][203] , 
	\_zy_simnet_tvar_20[5][202] , \_zy_simnet_tvar_20[5][201] , 
	\_zy_simnet_tvar_20[5][200] , \_zy_simnet_tvar_20[5][199] , 
	\_zy_simnet_tvar_20[5][198] , \_zy_simnet_tvar_20[5][197] , 
	\_zy_simnet_tvar_20[5][196] , \_zy_simnet_tvar_20[5][195] , 
	\_zy_simnet_tvar_20[5][194] , \_zy_simnet_tvar_20[5][193] , 
	\_zy_simnet_tvar_20[5][192] , \_zy_simnet_tvar_20[5][191] , 
	\_zy_simnet_tvar_20[5][190] , \_zy_simnet_tvar_20[5][189] , 
	\_zy_simnet_tvar_20[5][188] , \_zy_simnet_tvar_20[5][187] , 
	\_zy_simnet_tvar_20[5][186] , \_zy_simnet_tvar_20[5][185] , 
	\_zy_simnet_tvar_20[5][184] , \_zy_simnet_tvar_20[5][183] , 
	\_zy_simnet_tvar_20[5][182] , \_zy_simnet_tvar_20[5][181] , 
	\_zy_simnet_tvar_20[5][180] , \_zy_simnet_tvar_20[5][179] , 
	\_zy_simnet_tvar_20[5][178] , \_zy_simnet_tvar_20[5][177] , 
	\_zy_simnet_tvar_20[5][176] , \_zy_simnet_tvar_20[5][175] , 
	\_zy_simnet_tvar_20[5][174] , \_zy_simnet_tvar_20[5][173] , 
	\_zy_simnet_tvar_20[5][172] , \_zy_simnet_tvar_20[5][171] , 
	\_zy_simnet_tvar_20[5][170] , \_zy_simnet_tvar_20[5][169] , 
	\_zy_simnet_tvar_20[5][168] , \_zy_simnet_tvar_20[5][167] , 
	\_zy_simnet_tvar_20[5][166] , \_zy_simnet_tvar_20[5][165] , 
	\_zy_simnet_tvar_20[5][164] , \_zy_simnet_tvar_20[5][163] , 
	\_zy_simnet_tvar_20[5][162] , \_zy_simnet_tvar_20[5][161] , 
	\_zy_simnet_tvar_20[5][160] , \_zy_simnet_tvar_20[5][159] , 
	\_zy_simnet_tvar_20[5][158] , \_zy_simnet_tvar_20[5][157] , 
	\_zy_simnet_tvar_20[5][156] , \_zy_simnet_tvar_20[5][155] , 
	\_zy_simnet_tvar_20[5][154] , \_zy_simnet_tvar_20[5][153] , 
	\_zy_simnet_tvar_20[5][152] , \_zy_simnet_tvar_20[5][151] , 
	\_zy_simnet_tvar_20[5][150] , \_zy_simnet_tvar_20[5][149] , 
	\_zy_simnet_tvar_20[5][148] , \_zy_simnet_tvar_20[5][147] , 
	\_zy_simnet_tvar_20[5][146] , \_zy_simnet_tvar_20[5][145] , 
	\_zy_simnet_tvar_20[5][144] , \_zy_simnet_tvar_20[5][143] , 
	\_zy_simnet_tvar_20[5][142] , \_zy_simnet_tvar_20[5][141] , 
	\_zy_simnet_tvar_20[5][140] , \_zy_simnet_tvar_20[5][139] , 
	\_zy_simnet_tvar_20[5][138] , \_zy_simnet_tvar_20[5][137] , 
	\_zy_simnet_tvar_20[5][136] , \_zy_simnet_tvar_20[5][135] , 
	\_zy_simnet_tvar_20[5][134] , \_zy_simnet_tvar_20[5][133] , 
	\_zy_simnet_tvar_20[5][132] , \_zy_simnet_tvar_20[5][131] , 
	\_zy_simnet_tvar_20[5][130] , \_zy_simnet_tvar_20[5][129] , 
	\_zy_simnet_tvar_20[5][128] , \_zy_simnet_tvar_20[5][127] , 
	\_zy_simnet_tvar_20[5][126] , \_zy_simnet_tvar_20[5][125] , 
	\_zy_simnet_tvar_20[5][124] , \_zy_simnet_tvar_20[5][123] , 
	\_zy_simnet_tvar_20[5][122] , \_zy_simnet_tvar_20[5][121] , 
	\_zy_simnet_tvar_20[5][120] , \_zy_simnet_tvar_20[5][119] , 
	\_zy_simnet_tvar_20[5][118] , \_zy_simnet_tvar_20[5][117] , 
	\_zy_simnet_tvar_20[5][116] , \_zy_simnet_tvar_20[5][115] , 
	\_zy_simnet_tvar_20[5][114] , \_zy_simnet_tvar_20[5][113] , 
	\_zy_simnet_tvar_20[5][112] , \_zy_simnet_tvar_20[5][111] , 
	\_zy_simnet_tvar_20[5][110] , \_zy_simnet_tvar_20[5][109] , 
	\_zy_simnet_tvar_20[5][108] , \_zy_simnet_tvar_20[5][107] , 
	\_zy_simnet_tvar_20[5][106] , \_zy_simnet_tvar_20[5][105] , 
	\_zy_simnet_tvar_20[5][104] , \_zy_simnet_tvar_20[5][103] , 
	\_zy_simnet_tvar_20[5][102] , \_zy_simnet_tvar_20[5][101] , 
	\_zy_simnet_tvar_20[5][100] , \_zy_simnet_tvar_20[5][99] , 
	\_zy_simnet_tvar_20[5][98] , \_zy_simnet_tvar_20[5][97] , 
	\_zy_simnet_tvar_20[5][96] , \_zy_simnet_tvar_20[5][95] , 
	\_zy_simnet_tvar_20[5][94] , \_zy_simnet_tvar_20[5][93] , 
	\_zy_simnet_tvar_20[5][92] , \_zy_simnet_tvar_20[5][91] , 
	\_zy_simnet_tvar_20[5][90] , \_zy_simnet_tvar_20[5][89] , 
	\_zy_simnet_tvar_20[5][88] , \_zy_simnet_tvar_20[5][87] , 
	\_zy_simnet_tvar_20[5][86] , \_zy_simnet_tvar_20[5][85] , 
	\_zy_simnet_tvar_20[5][84] , \_zy_simnet_tvar_20[5][83] , 
	\_zy_simnet_tvar_20[5][82] , \_zy_simnet_tvar_20[5][81] , 
	\_zy_simnet_tvar_20[5][80] , \_zy_simnet_tvar_20[5][79] , 
	\_zy_simnet_tvar_20[5][78] , \_zy_simnet_tvar_20[5][77] , 
	\_zy_simnet_tvar_20[5][76] , \_zy_simnet_tvar_20[5][75] , 
	\_zy_simnet_tvar_20[5][74] , \_zy_simnet_tvar_20[5][73] , 
	\_zy_simnet_tvar_20[5][72] , \_zy_simnet_tvar_20[5][71] , 
	\_zy_simnet_tvar_20[5][70] , \_zy_simnet_tvar_20[5][69] , 
	\_zy_simnet_tvar_20[5][68] , \_zy_simnet_tvar_20[5][67] , 
	\_zy_simnet_tvar_20[5][66] , \_zy_simnet_tvar_20[5][65] , 
	\_zy_simnet_tvar_20[5][64] , \_zy_simnet_tvar_20[5][63] , 
	\_zy_simnet_tvar_20[5][62] , \_zy_simnet_tvar_20[5][61] , 
	\_zy_simnet_tvar_20[5][60] , \_zy_simnet_tvar_20[5][59] , 
	\_zy_simnet_tvar_20[5][58] , \_zy_simnet_tvar_20[5][57] , 
	\_zy_simnet_tvar_20[5][56] , \_zy_simnet_tvar_20[5][55] , 
	\_zy_simnet_tvar_20[5][54] , \_zy_simnet_tvar_20[5][53] , 
	\_zy_simnet_tvar_20[5][52] , \_zy_simnet_tvar_20[5][51] , 
	\_zy_simnet_tvar_20[5][50] , \_zy_simnet_tvar_20[5][49] , 
	\_zy_simnet_tvar_20[5][48] , \_zy_simnet_tvar_20[5][47] , 
	\_zy_simnet_tvar_20[5][46] , \_zy_simnet_tvar_20[5][45] , 
	\_zy_simnet_tvar_20[5][44] , \_zy_simnet_tvar_20[5][43] , 
	\_zy_simnet_tvar_20[5][42] , \_zy_simnet_tvar_20[5][41] , 
	\_zy_simnet_tvar_20[5][40] , \_zy_simnet_tvar_20[5][39] , 
	\_zy_simnet_tvar_20[5][38] , \_zy_simnet_tvar_20[5][37] , 
	\_zy_simnet_tvar_20[5][36] , \_zy_simnet_tvar_20[5][35] , 
	\_zy_simnet_tvar_20[5][34] , \_zy_simnet_tvar_20[5][33] , 
	\_zy_simnet_tvar_20[5][32] , \_zy_simnet_tvar_20[5][31] , 
	\_zy_simnet_tvar_20[5][30] , \_zy_simnet_tvar_20[5][29] , 
	\_zy_simnet_tvar_20[5][28] , \_zy_simnet_tvar_20[5][27] , 
	\_zy_simnet_tvar_20[5][26] , \_zy_simnet_tvar_20[5][25] , 
	\_zy_simnet_tvar_20[5][24] , \_zy_simnet_tvar_20[5][23] , 
	\_zy_simnet_tvar_20[5][22] , \_zy_simnet_tvar_20[5][21] , 
	\_zy_simnet_tvar_20[5][20] , \_zy_simnet_tvar_20[5][19] , 
	\_zy_simnet_tvar_20[5][18] , \_zy_simnet_tvar_20[5][17] , 
	\_zy_simnet_tvar_20[5][16] , \_zy_simnet_tvar_20[5][15] , 
	\_zy_simnet_tvar_20[5][14] , \_zy_simnet_tvar_20[5][13] , 
	\_zy_simnet_tvar_20[5][12] , \_zy_simnet_tvar_20[5][11] , 
	\_zy_simnet_tvar_20[5][10] , \_zy_simnet_tvar_20[5][9] , 
	\_zy_simnet_tvar_20[5][8] , \_zy_simnet_tvar_20[5][7] , 
	\_zy_simnet_tvar_20[5][6] , \_zy_simnet_tvar_20[5][5] , 
	\_zy_simnet_tvar_20[5][4] , \_zy_simnet_tvar_20[5][3] , 
	\_zy_simnet_tvar_20[5][2] , \_zy_simnet_tvar_20[5][1] , 
	\_zy_simnet_tvar_20[5][0] , \_zy_simnet_tvar_20[4][271] , 
	\_zy_simnet_tvar_20[4][270] , \_zy_simnet_tvar_20[4][269] , 
	\_zy_simnet_tvar_20[4][268] , \_zy_simnet_tvar_20[4][267] , 
	\_zy_simnet_tvar_20[4][266] , \_zy_simnet_tvar_20[4][265] , 
	\_zy_simnet_tvar_20[4][264] , \_zy_simnet_tvar_20[4][263] , 
	\_zy_simnet_tvar_20[4][262] , \_zy_simnet_tvar_20[4][261] , 
	\_zy_simnet_tvar_20[4][260] , \_zy_simnet_tvar_20[4][259] , 
	\_zy_simnet_tvar_20[4][258] , \_zy_simnet_tvar_20[4][257] , 
	\_zy_simnet_tvar_20[4][256] , \_zy_simnet_tvar_20[4][255] , 
	\_zy_simnet_tvar_20[4][254] , \_zy_simnet_tvar_20[4][253] , 
	\_zy_simnet_tvar_20[4][252] , \_zy_simnet_tvar_20[4][251] , 
	\_zy_simnet_tvar_20[4][250] , \_zy_simnet_tvar_20[4][249] , 
	\_zy_simnet_tvar_20[4][248] , \_zy_simnet_tvar_20[4][247] , 
	\_zy_simnet_tvar_20[4][246] , \_zy_simnet_tvar_20[4][245] , 
	\_zy_simnet_tvar_20[4][244] , \_zy_simnet_tvar_20[4][243] , 
	\_zy_simnet_tvar_20[4][242] , \_zy_simnet_tvar_20[4][241] , 
	\_zy_simnet_tvar_20[4][240] , \_zy_simnet_tvar_20[4][239] , 
	\_zy_simnet_tvar_20[4][238] , \_zy_simnet_tvar_20[4][237] , 
	\_zy_simnet_tvar_20[4][236] , \_zy_simnet_tvar_20[4][235] , 
	\_zy_simnet_tvar_20[4][234] , \_zy_simnet_tvar_20[4][233] , 
	\_zy_simnet_tvar_20[4][232] , \_zy_simnet_tvar_20[4][231] , 
	\_zy_simnet_tvar_20[4][230] , \_zy_simnet_tvar_20[4][229] , 
	\_zy_simnet_tvar_20[4][228] , \_zy_simnet_tvar_20[4][227] , 
	\_zy_simnet_tvar_20[4][226] , \_zy_simnet_tvar_20[4][225] , 
	\_zy_simnet_tvar_20[4][224] , \_zy_simnet_tvar_20[4][223] , 
	\_zy_simnet_tvar_20[4][222] , \_zy_simnet_tvar_20[4][221] , 
	\_zy_simnet_tvar_20[4][220] , \_zy_simnet_tvar_20[4][219] , 
	\_zy_simnet_tvar_20[4][218] , \_zy_simnet_tvar_20[4][217] , 
	\_zy_simnet_tvar_20[4][216] , \_zy_simnet_tvar_20[4][215] , 
	\_zy_simnet_tvar_20[4][214] , \_zy_simnet_tvar_20[4][213] , 
	\_zy_simnet_tvar_20[4][212] , \_zy_simnet_tvar_20[4][211] , 
	\_zy_simnet_tvar_20[4][210] , \_zy_simnet_tvar_20[4][209] , 
	\_zy_simnet_tvar_20[4][208] , \_zy_simnet_tvar_20[4][207] , 
	\_zy_simnet_tvar_20[4][206] , \_zy_simnet_tvar_20[4][205] , 
	\_zy_simnet_tvar_20[4][204] , \_zy_simnet_tvar_20[4][203] , 
	\_zy_simnet_tvar_20[4][202] , \_zy_simnet_tvar_20[4][201] , 
	\_zy_simnet_tvar_20[4][200] , \_zy_simnet_tvar_20[4][199] , 
	\_zy_simnet_tvar_20[4][198] , \_zy_simnet_tvar_20[4][197] , 
	\_zy_simnet_tvar_20[4][196] , \_zy_simnet_tvar_20[4][195] , 
	\_zy_simnet_tvar_20[4][194] , \_zy_simnet_tvar_20[4][193] , 
	\_zy_simnet_tvar_20[4][192] , \_zy_simnet_tvar_20[4][191] , 
	\_zy_simnet_tvar_20[4][190] , \_zy_simnet_tvar_20[4][189] , 
	\_zy_simnet_tvar_20[4][188] , \_zy_simnet_tvar_20[4][187] , 
	\_zy_simnet_tvar_20[4][186] , \_zy_simnet_tvar_20[4][185] , 
	\_zy_simnet_tvar_20[4][184] , \_zy_simnet_tvar_20[4][183] , 
	\_zy_simnet_tvar_20[4][182] , \_zy_simnet_tvar_20[4][181] , 
	\_zy_simnet_tvar_20[4][180] , \_zy_simnet_tvar_20[4][179] , 
	\_zy_simnet_tvar_20[4][178] , \_zy_simnet_tvar_20[4][177] , 
	\_zy_simnet_tvar_20[4][176] , \_zy_simnet_tvar_20[4][175] , 
	\_zy_simnet_tvar_20[4][174] , \_zy_simnet_tvar_20[4][173] , 
	\_zy_simnet_tvar_20[4][172] , \_zy_simnet_tvar_20[4][171] , 
	\_zy_simnet_tvar_20[4][170] , \_zy_simnet_tvar_20[4][169] , 
	\_zy_simnet_tvar_20[4][168] , \_zy_simnet_tvar_20[4][167] , 
	\_zy_simnet_tvar_20[4][166] , \_zy_simnet_tvar_20[4][165] , 
	\_zy_simnet_tvar_20[4][164] , \_zy_simnet_tvar_20[4][163] , 
	\_zy_simnet_tvar_20[4][162] , \_zy_simnet_tvar_20[4][161] , 
	\_zy_simnet_tvar_20[4][160] , \_zy_simnet_tvar_20[4][159] , 
	\_zy_simnet_tvar_20[4][158] , \_zy_simnet_tvar_20[4][157] , 
	\_zy_simnet_tvar_20[4][156] , \_zy_simnet_tvar_20[4][155] , 
	\_zy_simnet_tvar_20[4][154] , \_zy_simnet_tvar_20[4][153] , 
	\_zy_simnet_tvar_20[4][152] , \_zy_simnet_tvar_20[4][151] , 
	\_zy_simnet_tvar_20[4][150] , \_zy_simnet_tvar_20[4][149] , 
	\_zy_simnet_tvar_20[4][148] , \_zy_simnet_tvar_20[4][147] , 
	\_zy_simnet_tvar_20[4][146] , \_zy_simnet_tvar_20[4][145] , 
	\_zy_simnet_tvar_20[4][144] , \_zy_simnet_tvar_20[4][143] , 
	\_zy_simnet_tvar_20[4][142] , \_zy_simnet_tvar_20[4][141] , 
	\_zy_simnet_tvar_20[4][140] , \_zy_simnet_tvar_20[4][139] , 
	\_zy_simnet_tvar_20[4][138] , \_zy_simnet_tvar_20[4][137] , 
	\_zy_simnet_tvar_20[4][136] , \_zy_simnet_tvar_20[4][135] , 
	\_zy_simnet_tvar_20[4][134] , \_zy_simnet_tvar_20[4][133] , 
	\_zy_simnet_tvar_20[4][132] , \_zy_simnet_tvar_20[4][131] , 
	\_zy_simnet_tvar_20[4][130] , \_zy_simnet_tvar_20[4][129] , 
	\_zy_simnet_tvar_20[4][128] , \_zy_simnet_tvar_20[4][127] , 
	\_zy_simnet_tvar_20[4][126] , \_zy_simnet_tvar_20[4][125] , 
	\_zy_simnet_tvar_20[4][124] , \_zy_simnet_tvar_20[4][123] , 
	\_zy_simnet_tvar_20[4][122] , \_zy_simnet_tvar_20[4][121] , 
	\_zy_simnet_tvar_20[4][120] , \_zy_simnet_tvar_20[4][119] , 
	\_zy_simnet_tvar_20[4][118] , \_zy_simnet_tvar_20[4][117] , 
	\_zy_simnet_tvar_20[4][116] , \_zy_simnet_tvar_20[4][115] , 
	\_zy_simnet_tvar_20[4][114] , \_zy_simnet_tvar_20[4][113] , 
	\_zy_simnet_tvar_20[4][112] , \_zy_simnet_tvar_20[4][111] , 
	\_zy_simnet_tvar_20[4][110] , \_zy_simnet_tvar_20[4][109] , 
	\_zy_simnet_tvar_20[4][108] , \_zy_simnet_tvar_20[4][107] , 
	\_zy_simnet_tvar_20[4][106] , \_zy_simnet_tvar_20[4][105] , 
	\_zy_simnet_tvar_20[4][104] , \_zy_simnet_tvar_20[4][103] , 
	\_zy_simnet_tvar_20[4][102] , \_zy_simnet_tvar_20[4][101] , 
	\_zy_simnet_tvar_20[4][100] , \_zy_simnet_tvar_20[4][99] , 
	\_zy_simnet_tvar_20[4][98] , \_zy_simnet_tvar_20[4][97] , 
	\_zy_simnet_tvar_20[4][96] , \_zy_simnet_tvar_20[4][95] , 
	\_zy_simnet_tvar_20[4][94] , \_zy_simnet_tvar_20[4][93] , 
	\_zy_simnet_tvar_20[4][92] , \_zy_simnet_tvar_20[4][91] , 
	\_zy_simnet_tvar_20[4][90] , \_zy_simnet_tvar_20[4][89] , 
	\_zy_simnet_tvar_20[4][88] , \_zy_simnet_tvar_20[4][87] , 
	\_zy_simnet_tvar_20[4][86] , \_zy_simnet_tvar_20[4][85] , 
	\_zy_simnet_tvar_20[4][84] , \_zy_simnet_tvar_20[4][83] , 
	\_zy_simnet_tvar_20[4][82] , \_zy_simnet_tvar_20[4][81] , 
	\_zy_simnet_tvar_20[4][80] , \_zy_simnet_tvar_20[4][79] , 
	\_zy_simnet_tvar_20[4][78] , \_zy_simnet_tvar_20[4][77] , 
	\_zy_simnet_tvar_20[4][76] , \_zy_simnet_tvar_20[4][75] , 
	\_zy_simnet_tvar_20[4][74] , \_zy_simnet_tvar_20[4][73] , 
	\_zy_simnet_tvar_20[4][72] , \_zy_simnet_tvar_20[4][71] , 
	\_zy_simnet_tvar_20[4][70] , \_zy_simnet_tvar_20[4][69] , 
	\_zy_simnet_tvar_20[4][68] , \_zy_simnet_tvar_20[4][67] , 
	\_zy_simnet_tvar_20[4][66] , \_zy_simnet_tvar_20[4][65] , 
	\_zy_simnet_tvar_20[4][64] , \_zy_simnet_tvar_20[4][63] , 
	\_zy_simnet_tvar_20[4][62] , \_zy_simnet_tvar_20[4][61] , 
	\_zy_simnet_tvar_20[4][60] , \_zy_simnet_tvar_20[4][59] , 
	\_zy_simnet_tvar_20[4][58] , \_zy_simnet_tvar_20[4][57] , 
	\_zy_simnet_tvar_20[4][56] , \_zy_simnet_tvar_20[4][55] , 
	\_zy_simnet_tvar_20[4][54] , \_zy_simnet_tvar_20[4][53] , 
	\_zy_simnet_tvar_20[4][52] , \_zy_simnet_tvar_20[4][51] , 
	\_zy_simnet_tvar_20[4][50] , \_zy_simnet_tvar_20[4][49] , 
	\_zy_simnet_tvar_20[4][48] , \_zy_simnet_tvar_20[4][47] , 
	\_zy_simnet_tvar_20[4][46] , \_zy_simnet_tvar_20[4][45] , 
	\_zy_simnet_tvar_20[4][44] , \_zy_simnet_tvar_20[4][43] , 
	\_zy_simnet_tvar_20[4][42] , \_zy_simnet_tvar_20[4][41] , 
	\_zy_simnet_tvar_20[4][40] , \_zy_simnet_tvar_20[4][39] , 
	\_zy_simnet_tvar_20[4][38] , \_zy_simnet_tvar_20[4][37] , 
	\_zy_simnet_tvar_20[4][36] , \_zy_simnet_tvar_20[4][35] , 
	\_zy_simnet_tvar_20[4][34] , \_zy_simnet_tvar_20[4][33] , 
	\_zy_simnet_tvar_20[4][32] , \_zy_simnet_tvar_20[4][31] , 
	\_zy_simnet_tvar_20[4][30] , \_zy_simnet_tvar_20[4][29] , 
	\_zy_simnet_tvar_20[4][28] , \_zy_simnet_tvar_20[4][27] , 
	\_zy_simnet_tvar_20[4][26] , \_zy_simnet_tvar_20[4][25] , 
	\_zy_simnet_tvar_20[4][24] , \_zy_simnet_tvar_20[4][23] , 
	\_zy_simnet_tvar_20[4][22] , \_zy_simnet_tvar_20[4][21] , 
	\_zy_simnet_tvar_20[4][20] , \_zy_simnet_tvar_20[4][19] , 
	\_zy_simnet_tvar_20[4][18] , \_zy_simnet_tvar_20[4][17] , 
	\_zy_simnet_tvar_20[4][16] , \_zy_simnet_tvar_20[4][15] , 
	\_zy_simnet_tvar_20[4][14] , \_zy_simnet_tvar_20[4][13] , 
	\_zy_simnet_tvar_20[4][12] , \_zy_simnet_tvar_20[4][11] , 
	\_zy_simnet_tvar_20[4][10] , \_zy_simnet_tvar_20[4][9] , 
	\_zy_simnet_tvar_20[4][8] , \_zy_simnet_tvar_20[4][7] , 
	\_zy_simnet_tvar_20[4][6] , \_zy_simnet_tvar_20[4][5] , 
	\_zy_simnet_tvar_20[4][4] , \_zy_simnet_tvar_20[4][3] , 
	\_zy_simnet_tvar_20[4][2] , \_zy_simnet_tvar_20[4][1] , 
	\_zy_simnet_tvar_20[4][0] , \_zy_simnet_tvar_20[3][271] , 
	\_zy_simnet_tvar_20[3][270] , \_zy_simnet_tvar_20[3][269] , 
	\_zy_simnet_tvar_20[3][268] , \_zy_simnet_tvar_20[3][267] , 
	\_zy_simnet_tvar_20[3][266] , \_zy_simnet_tvar_20[3][265] , 
	\_zy_simnet_tvar_20[3][264] , \_zy_simnet_tvar_20[3][263] , 
	\_zy_simnet_tvar_20[3][262] , \_zy_simnet_tvar_20[3][261] , 
	\_zy_simnet_tvar_20[3][260] , \_zy_simnet_tvar_20[3][259] , 
	\_zy_simnet_tvar_20[3][258] , \_zy_simnet_tvar_20[3][257] , 
	\_zy_simnet_tvar_20[3][256] , \_zy_simnet_tvar_20[3][255] , 
	\_zy_simnet_tvar_20[3][254] , \_zy_simnet_tvar_20[3][253] , 
	\_zy_simnet_tvar_20[3][252] , \_zy_simnet_tvar_20[3][251] , 
	\_zy_simnet_tvar_20[3][250] , \_zy_simnet_tvar_20[3][249] , 
	\_zy_simnet_tvar_20[3][248] , \_zy_simnet_tvar_20[3][247] , 
	\_zy_simnet_tvar_20[3][246] , \_zy_simnet_tvar_20[3][245] , 
	\_zy_simnet_tvar_20[3][244] , \_zy_simnet_tvar_20[3][243] , 
	\_zy_simnet_tvar_20[3][242] , \_zy_simnet_tvar_20[3][241] , 
	\_zy_simnet_tvar_20[3][240] , \_zy_simnet_tvar_20[3][239] , 
	\_zy_simnet_tvar_20[3][238] , \_zy_simnet_tvar_20[3][237] , 
	\_zy_simnet_tvar_20[3][236] , \_zy_simnet_tvar_20[3][235] , 
	\_zy_simnet_tvar_20[3][234] , \_zy_simnet_tvar_20[3][233] , 
	\_zy_simnet_tvar_20[3][232] , \_zy_simnet_tvar_20[3][231] , 
	\_zy_simnet_tvar_20[3][230] , \_zy_simnet_tvar_20[3][229] , 
	\_zy_simnet_tvar_20[3][228] , \_zy_simnet_tvar_20[3][227] , 
	\_zy_simnet_tvar_20[3][226] , \_zy_simnet_tvar_20[3][225] , 
	\_zy_simnet_tvar_20[3][224] , \_zy_simnet_tvar_20[3][223] , 
	\_zy_simnet_tvar_20[3][222] , \_zy_simnet_tvar_20[3][221] , 
	\_zy_simnet_tvar_20[3][220] , \_zy_simnet_tvar_20[3][219] , 
	\_zy_simnet_tvar_20[3][218] , \_zy_simnet_tvar_20[3][217] , 
	\_zy_simnet_tvar_20[3][216] , \_zy_simnet_tvar_20[3][215] , 
	\_zy_simnet_tvar_20[3][214] , \_zy_simnet_tvar_20[3][213] , 
	\_zy_simnet_tvar_20[3][212] , \_zy_simnet_tvar_20[3][211] , 
	\_zy_simnet_tvar_20[3][210] , \_zy_simnet_tvar_20[3][209] , 
	\_zy_simnet_tvar_20[3][208] , \_zy_simnet_tvar_20[3][207] , 
	\_zy_simnet_tvar_20[3][206] , \_zy_simnet_tvar_20[3][205] , 
	\_zy_simnet_tvar_20[3][204] , \_zy_simnet_tvar_20[3][203] , 
	\_zy_simnet_tvar_20[3][202] , \_zy_simnet_tvar_20[3][201] , 
	\_zy_simnet_tvar_20[3][200] , \_zy_simnet_tvar_20[3][199] , 
	\_zy_simnet_tvar_20[3][198] , \_zy_simnet_tvar_20[3][197] , 
	\_zy_simnet_tvar_20[3][196] , \_zy_simnet_tvar_20[3][195] , 
	\_zy_simnet_tvar_20[3][194] , \_zy_simnet_tvar_20[3][193] , 
	\_zy_simnet_tvar_20[3][192] , \_zy_simnet_tvar_20[3][191] , 
	\_zy_simnet_tvar_20[3][190] , \_zy_simnet_tvar_20[3][189] , 
	\_zy_simnet_tvar_20[3][188] , \_zy_simnet_tvar_20[3][187] , 
	\_zy_simnet_tvar_20[3][186] , \_zy_simnet_tvar_20[3][185] , 
	\_zy_simnet_tvar_20[3][184] , \_zy_simnet_tvar_20[3][183] , 
	\_zy_simnet_tvar_20[3][182] , \_zy_simnet_tvar_20[3][181] , 
	\_zy_simnet_tvar_20[3][180] , \_zy_simnet_tvar_20[3][179] , 
	\_zy_simnet_tvar_20[3][178] , \_zy_simnet_tvar_20[3][177] , 
	\_zy_simnet_tvar_20[3][176] , \_zy_simnet_tvar_20[3][175] , 
	\_zy_simnet_tvar_20[3][174] , \_zy_simnet_tvar_20[3][173] , 
	\_zy_simnet_tvar_20[3][172] , \_zy_simnet_tvar_20[3][171] , 
	\_zy_simnet_tvar_20[3][170] , \_zy_simnet_tvar_20[3][169] , 
	\_zy_simnet_tvar_20[3][168] , \_zy_simnet_tvar_20[3][167] , 
	\_zy_simnet_tvar_20[3][166] , \_zy_simnet_tvar_20[3][165] , 
	\_zy_simnet_tvar_20[3][164] , \_zy_simnet_tvar_20[3][163] , 
	\_zy_simnet_tvar_20[3][162] , \_zy_simnet_tvar_20[3][161] , 
	\_zy_simnet_tvar_20[3][160] , \_zy_simnet_tvar_20[3][159] , 
	\_zy_simnet_tvar_20[3][158] , \_zy_simnet_tvar_20[3][157] , 
	\_zy_simnet_tvar_20[3][156] , \_zy_simnet_tvar_20[3][155] , 
	\_zy_simnet_tvar_20[3][154] , \_zy_simnet_tvar_20[3][153] , 
	\_zy_simnet_tvar_20[3][152] , \_zy_simnet_tvar_20[3][151] , 
	\_zy_simnet_tvar_20[3][150] , \_zy_simnet_tvar_20[3][149] , 
	\_zy_simnet_tvar_20[3][148] , \_zy_simnet_tvar_20[3][147] , 
	\_zy_simnet_tvar_20[3][146] , \_zy_simnet_tvar_20[3][145] , 
	\_zy_simnet_tvar_20[3][144] , \_zy_simnet_tvar_20[3][143] , 
	\_zy_simnet_tvar_20[3][142] , \_zy_simnet_tvar_20[3][141] , 
	\_zy_simnet_tvar_20[3][140] , \_zy_simnet_tvar_20[3][139] , 
	\_zy_simnet_tvar_20[3][138] , \_zy_simnet_tvar_20[3][137] , 
	\_zy_simnet_tvar_20[3][136] , \_zy_simnet_tvar_20[3][135] , 
	\_zy_simnet_tvar_20[3][134] , \_zy_simnet_tvar_20[3][133] , 
	\_zy_simnet_tvar_20[3][132] , \_zy_simnet_tvar_20[3][131] , 
	\_zy_simnet_tvar_20[3][130] , \_zy_simnet_tvar_20[3][129] , 
	\_zy_simnet_tvar_20[3][128] , \_zy_simnet_tvar_20[3][127] , 
	\_zy_simnet_tvar_20[3][126] , \_zy_simnet_tvar_20[3][125] , 
	\_zy_simnet_tvar_20[3][124] , \_zy_simnet_tvar_20[3][123] , 
	\_zy_simnet_tvar_20[3][122] , \_zy_simnet_tvar_20[3][121] , 
	\_zy_simnet_tvar_20[3][120] , \_zy_simnet_tvar_20[3][119] , 
	\_zy_simnet_tvar_20[3][118] , \_zy_simnet_tvar_20[3][117] , 
	\_zy_simnet_tvar_20[3][116] , \_zy_simnet_tvar_20[3][115] , 
	\_zy_simnet_tvar_20[3][114] , \_zy_simnet_tvar_20[3][113] , 
	\_zy_simnet_tvar_20[3][112] , \_zy_simnet_tvar_20[3][111] , 
	\_zy_simnet_tvar_20[3][110] , \_zy_simnet_tvar_20[3][109] , 
	\_zy_simnet_tvar_20[3][108] , \_zy_simnet_tvar_20[3][107] , 
	\_zy_simnet_tvar_20[3][106] , \_zy_simnet_tvar_20[3][105] , 
	\_zy_simnet_tvar_20[3][104] , \_zy_simnet_tvar_20[3][103] , 
	\_zy_simnet_tvar_20[3][102] , \_zy_simnet_tvar_20[3][101] , 
	\_zy_simnet_tvar_20[3][100] , \_zy_simnet_tvar_20[3][99] , 
	\_zy_simnet_tvar_20[3][98] , \_zy_simnet_tvar_20[3][97] , 
	\_zy_simnet_tvar_20[3][96] , \_zy_simnet_tvar_20[3][95] , 
	\_zy_simnet_tvar_20[3][94] , \_zy_simnet_tvar_20[3][93] , 
	\_zy_simnet_tvar_20[3][92] , \_zy_simnet_tvar_20[3][91] , 
	\_zy_simnet_tvar_20[3][90] , \_zy_simnet_tvar_20[3][89] , 
	\_zy_simnet_tvar_20[3][88] , \_zy_simnet_tvar_20[3][87] , 
	\_zy_simnet_tvar_20[3][86] , \_zy_simnet_tvar_20[3][85] , 
	\_zy_simnet_tvar_20[3][84] , \_zy_simnet_tvar_20[3][83] , 
	\_zy_simnet_tvar_20[3][82] , \_zy_simnet_tvar_20[3][81] , 
	\_zy_simnet_tvar_20[3][80] , \_zy_simnet_tvar_20[3][79] , 
	\_zy_simnet_tvar_20[3][78] , \_zy_simnet_tvar_20[3][77] , 
	\_zy_simnet_tvar_20[3][76] , \_zy_simnet_tvar_20[3][75] , 
	\_zy_simnet_tvar_20[3][74] , \_zy_simnet_tvar_20[3][73] , 
	\_zy_simnet_tvar_20[3][72] , \_zy_simnet_tvar_20[3][71] , 
	\_zy_simnet_tvar_20[3][70] , \_zy_simnet_tvar_20[3][69] , 
	\_zy_simnet_tvar_20[3][68] , \_zy_simnet_tvar_20[3][67] , 
	\_zy_simnet_tvar_20[3][66] , \_zy_simnet_tvar_20[3][65] , 
	\_zy_simnet_tvar_20[3][64] , \_zy_simnet_tvar_20[3][63] , 
	\_zy_simnet_tvar_20[3][62] , \_zy_simnet_tvar_20[3][61] , 
	\_zy_simnet_tvar_20[3][60] , \_zy_simnet_tvar_20[3][59] , 
	\_zy_simnet_tvar_20[3][58] , \_zy_simnet_tvar_20[3][57] , 
	\_zy_simnet_tvar_20[3][56] , \_zy_simnet_tvar_20[3][55] , 
	\_zy_simnet_tvar_20[3][54] , \_zy_simnet_tvar_20[3][53] , 
	\_zy_simnet_tvar_20[3][52] , \_zy_simnet_tvar_20[3][51] , 
	\_zy_simnet_tvar_20[3][50] , \_zy_simnet_tvar_20[3][49] , 
	\_zy_simnet_tvar_20[3][48] , \_zy_simnet_tvar_20[3][47] , 
	\_zy_simnet_tvar_20[3][46] , \_zy_simnet_tvar_20[3][45] , 
	\_zy_simnet_tvar_20[3][44] , \_zy_simnet_tvar_20[3][43] , 
	\_zy_simnet_tvar_20[3][42] , \_zy_simnet_tvar_20[3][41] , 
	\_zy_simnet_tvar_20[3][40] , \_zy_simnet_tvar_20[3][39] , 
	\_zy_simnet_tvar_20[3][38] , \_zy_simnet_tvar_20[3][37] , 
	\_zy_simnet_tvar_20[3][36] , \_zy_simnet_tvar_20[3][35] , 
	\_zy_simnet_tvar_20[3][34] , \_zy_simnet_tvar_20[3][33] , 
	\_zy_simnet_tvar_20[3][32] , \_zy_simnet_tvar_20[3][31] , 
	\_zy_simnet_tvar_20[3][30] , \_zy_simnet_tvar_20[3][29] , 
	\_zy_simnet_tvar_20[3][28] , \_zy_simnet_tvar_20[3][27] , 
	\_zy_simnet_tvar_20[3][26] , \_zy_simnet_tvar_20[3][25] , 
	\_zy_simnet_tvar_20[3][24] , \_zy_simnet_tvar_20[3][23] , 
	\_zy_simnet_tvar_20[3][22] , \_zy_simnet_tvar_20[3][21] , 
	\_zy_simnet_tvar_20[3][20] , \_zy_simnet_tvar_20[3][19] , 
	\_zy_simnet_tvar_20[3][18] , \_zy_simnet_tvar_20[3][17] , 
	\_zy_simnet_tvar_20[3][16] , \_zy_simnet_tvar_20[3][15] , 
	\_zy_simnet_tvar_20[3][14] , \_zy_simnet_tvar_20[3][13] , 
	\_zy_simnet_tvar_20[3][12] , \_zy_simnet_tvar_20[3][11] , 
	\_zy_simnet_tvar_20[3][10] , \_zy_simnet_tvar_20[3][9] , 
	\_zy_simnet_tvar_20[3][8] , \_zy_simnet_tvar_20[3][7] , 
	\_zy_simnet_tvar_20[3][6] , \_zy_simnet_tvar_20[3][5] , 
	\_zy_simnet_tvar_20[3][4] , \_zy_simnet_tvar_20[3][3] , 
	\_zy_simnet_tvar_20[3][2] , \_zy_simnet_tvar_20[3][1] , 
	\_zy_simnet_tvar_20[3][0] , \_zy_simnet_tvar_20[2][271] , 
	\_zy_simnet_tvar_20[2][270] , \_zy_simnet_tvar_20[2][269] , 
	\_zy_simnet_tvar_20[2][268] , \_zy_simnet_tvar_20[2][267] , 
	\_zy_simnet_tvar_20[2][266] , \_zy_simnet_tvar_20[2][265] , 
	\_zy_simnet_tvar_20[2][264] , \_zy_simnet_tvar_20[2][263] , 
	\_zy_simnet_tvar_20[2][262] , \_zy_simnet_tvar_20[2][261] , 
	\_zy_simnet_tvar_20[2][260] , \_zy_simnet_tvar_20[2][259] , 
	\_zy_simnet_tvar_20[2][258] , \_zy_simnet_tvar_20[2][257] , 
	\_zy_simnet_tvar_20[2][256] , \_zy_simnet_tvar_20[2][255] , 
	\_zy_simnet_tvar_20[2][254] , \_zy_simnet_tvar_20[2][253] , 
	\_zy_simnet_tvar_20[2][252] , \_zy_simnet_tvar_20[2][251] , 
	\_zy_simnet_tvar_20[2][250] , \_zy_simnet_tvar_20[2][249] , 
	\_zy_simnet_tvar_20[2][248] , \_zy_simnet_tvar_20[2][247] , 
	\_zy_simnet_tvar_20[2][246] , \_zy_simnet_tvar_20[2][245] , 
	\_zy_simnet_tvar_20[2][244] , \_zy_simnet_tvar_20[2][243] , 
	\_zy_simnet_tvar_20[2][242] , \_zy_simnet_tvar_20[2][241] , 
	\_zy_simnet_tvar_20[2][240] , \_zy_simnet_tvar_20[2][239] , 
	\_zy_simnet_tvar_20[2][238] , \_zy_simnet_tvar_20[2][237] , 
	\_zy_simnet_tvar_20[2][236] , \_zy_simnet_tvar_20[2][235] , 
	\_zy_simnet_tvar_20[2][234] , \_zy_simnet_tvar_20[2][233] , 
	\_zy_simnet_tvar_20[2][232] , \_zy_simnet_tvar_20[2][231] , 
	\_zy_simnet_tvar_20[2][230] , \_zy_simnet_tvar_20[2][229] , 
	\_zy_simnet_tvar_20[2][228] , \_zy_simnet_tvar_20[2][227] , 
	\_zy_simnet_tvar_20[2][226] , \_zy_simnet_tvar_20[2][225] , 
	\_zy_simnet_tvar_20[2][224] , \_zy_simnet_tvar_20[2][223] , 
	\_zy_simnet_tvar_20[2][222] , \_zy_simnet_tvar_20[2][221] , 
	\_zy_simnet_tvar_20[2][220] , \_zy_simnet_tvar_20[2][219] , 
	\_zy_simnet_tvar_20[2][218] , \_zy_simnet_tvar_20[2][217] , 
	\_zy_simnet_tvar_20[2][216] , \_zy_simnet_tvar_20[2][215] , 
	\_zy_simnet_tvar_20[2][214] , \_zy_simnet_tvar_20[2][213] , 
	\_zy_simnet_tvar_20[2][212] , \_zy_simnet_tvar_20[2][211] , 
	\_zy_simnet_tvar_20[2][210] , \_zy_simnet_tvar_20[2][209] , 
	\_zy_simnet_tvar_20[2][208] , \_zy_simnet_tvar_20[2][207] , 
	\_zy_simnet_tvar_20[2][206] , \_zy_simnet_tvar_20[2][205] , 
	\_zy_simnet_tvar_20[2][204] , \_zy_simnet_tvar_20[2][203] , 
	\_zy_simnet_tvar_20[2][202] , \_zy_simnet_tvar_20[2][201] , 
	\_zy_simnet_tvar_20[2][200] , \_zy_simnet_tvar_20[2][199] , 
	\_zy_simnet_tvar_20[2][198] , \_zy_simnet_tvar_20[2][197] , 
	\_zy_simnet_tvar_20[2][196] , \_zy_simnet_tvar_20[2][195] , 
	\_zy_simnet_tvar_20[2][194] , \_zy_simnet_tvar_20[2][193] , 
	\_zy_simnet_tvar_20[2][192] , \_zy_simnet_tvar_20[2][191] , 
	\_zy_simnet_tvar_20[2][190] , \_zy_simnet_tvar_20[2][189] , 
	\_zy_simnet_tvar_20[2][188] , \_zy_simnet_tvar_20[2][187] , 
	\_zy_simnet_tvar_20[2][186] , \_zy_simnet_tvar_20[2][185] , 
	\_zy_simnet_tvar_20[2][184] , \_zy_simnet_tvar_20[2][183] , 
	\_zy_simnet_tvar_20[2][182] , \_zy_simnet_tvar_20[2][181] , 
	\_zy_simnet_tvar_20[2][180] , \_zy_simnet_tvar_20[2][179] , 
	\_zy_simnet_tvar_20[2][178] , \_zy_simnet_tvar_20[2][177] , 
	\_zy_simnet_tvar_20[2][176] , \_zy_simnet_tvar_20[2][175] , 
	\_zy_simnet_tvar_20[2][174] , \_zy_simnet_tvar_20[2][173] , 
	\_zy_simnet_tvar_20[2][172] , \_zy_simnet_tvar_20[2][171] , 
	\_zy_simnet_tvar_20[2][170] , \_zy_simnet_tvar_20[2][169] , 
	\_zy_simnet_tvar_20[2][168] , \_zy_simnet_tvar_20[2][167] , 
	\_zy_simnet_tvar_20[2][166] , \_zy_simnet_tvar_20[2][165] , 
	\_zy_simnet_tvar_20[2][164] , \_zy_simnet_tvar_20[2][163] , 
	\_zy_simnet_tvar_20[2][162] , \_zy_simnet_tvar_20[2][161] , 
	\_zy_simnet_tvar_20[2][160] , \_zy_simnet_tvar_20[2][159] , 
	\_zy_simnet_tvar_20[2][158] , \_zy_simnet_tvar_20[2][157] , 
	\_zy_simnet_tvar_20[2][156] , \_zy_simnet_tvar_20[2][155] , 
	\_zy_simnet_tvar_20[2][154] , \_zy_simnet_tvar_20[2][153] , 
	\_zy_simnet_tvar_20[2][152] , \_zy_simnet_tvar_20[2][151] , 
	\_zy_simnet_tvar_20[2][150] , \_zy_simnet_tvar_20[2][149] , 
	\_zy_simnet_tvar_20[2][148] , \_zy_simnet_tvar_20[2][147] , 
	\_zy_simnet_tvar_20[2][146] , \_zy_simnet_tvar_20[2][145] , 
	\_zy_simnet_tvar_20[2][144] , \_zy_simnet_tvar_20[2][143] , 
	\_zy_simnet_tvar_20[2][142] , \_zy_simnet_tvar_20[2][141] , 
	\_zy_simnet_tvar_20[2][140] , \_zy_simnet_tvar_20[2][139] , 
	\_zy_simnet_tvar_20[2][138] , \_zy_simnet_tvar_20[2][137] , 
	\_zy_simnet_tvar_20[2][136] , \_zy_simnet_tvar_20[2][135] , 
	\_zy_simnet_tvar_20[2][134] , \_zy_simnet_tvar_20[2][133] , 
	\_zy_simnet_tvar_20[2][132] , \_zy_simnet_tvar_20[2][131] , 
	\_zy_simnet_tvar_20[2][130] , \_zy_simnet_tvar_20[2][129] , 
	\_zy_simnet_tvar_20[2][128] , \_zy_simnet_tvar_20[2][127] , 
	\_zy_simnet_tvar_20[2][126] , \_zy_simnet_tvar_20[2][125] , 
	\_zy_simnet_tvar_20[2][124] , \_zy_simnet_tvar_20[2][123] , 
	\_zy_simnet_tvar_20[2][122] , \_zy_simnet_tvar_20[2][121] , 
	\_zy_simnet_tvar_20[2][120] , \_zy_simnet_tvar_20[2][119] , 
	\_zy_simnet_tvar_20[2][118] , \_zy_simnet_tvar_20[2][117] , 
	\_zy_simnet_tvar_20[2][116] , \_zy_simnet_tvar_20[2][115] , 
	\_zy_simnet_tvar_20[2][114] , \_zy_simnet_tvar_20[2][113] , 
	\_zy_simnet_tvar_20[2][112] , \_zy_simnet_tvar_20[2][111] , 
	\_zy_simnet_tvar_20[2][110] , \_zy_simnet_tvar_20[2][109] , 
	\_zy_simnet_tvar_20[2][108] , \_zy_simnet_tvar_20[2][107] , 
	\_zy_simnet_tvar_20[2][106] , \_zy_simnet_tvar_20[2][105] , 
	\_zy_simnet_tvar_20[2][104] , \_zy_simnet_tvar_20[2][103] , 
	\_zy_simnet_tvar_20[2][102] , \_zy_simnet_tvar_20[2][101] , 
	\_zy_simnet_tvar_20[2][100] , \_zy_simnet_tvar_20[2][99] , 
	\_zy_simnet_tvar_20[2][98] , \_zy_simnet_tvar_20[2][97] , 
	\_zy_simnet_tvar_20[2][96] , \_zy_simnet_tvar_20[2][95] , 
	\_zy_simnet_tvar_20[2][94] , \_zy_simnet_tvar_20[2][93] , 
	\_zy_simnet_tvar_20[2][92] , \_zy_simnet_tvar_20[2][91] , 
	\_zy_simnet_tvar_20[2][90] , \_zy_simnet_tvar_20[2][89] , 
	\_zy_simnet_tvar_20[2][88] , \_zy_simnet_tvar_20[2][87] , 
	\_zy_simnet_tvar_20[2][86] , \_zy_simnet_tvar_20[2][85] , 
	\_zy_simnet_tvar_20[2][84] , \_zy_simnet_tvar_20[2][83] , 
	\_zy_simnet_tvar_20[2][82] , \_zy_simnet_tvar_20[2][81] , 
	\_zy_simnet_tvar_20[2][80] , \_zy_simnet_tvar_20[2][79] , 
	\_zy_simnet_tvar_20[2][78] , \_zy_simnet_tvar_20[2][77] , 
	\_zy_simnet_tvar_20[2][76] , \_zy_simnet_tvar_20[2][75] , 
	\_zy_simnet_tvar_20[2][74] , \_zy_simnet_tvar_20[2][73] , 
	\_zy_simnet_tvar_20[2][72] , \_zy_simnet_tvar_20[2][71] , 
	\_zy_simnet_tvar_20[2][70] , \_zy_simnet_tvar_20[2][69] , 
	\_zy_simnet_tvar_20[2][68] , \_zy_simnet_tvar_20[2][67] , 
	\_zy_simnet_tvar_20[2][66] , \_zy_simnet_tvar_20[2][65] , 
	\_zy_simnet_tvar_20[2][64] , \_zy_simnet_tvar_20[2][63] , 
	\_zy_simnet_tvar_20[2][62] , \_zy_simnet_tvar_20[2][61] , 
	\_zy_simnet_tvar_20[2][60] , \_zy_simnet_tvar_20[2][59] , 
	\_zy_simnet_tvar_20[2][58] , \_zy_simnet_tvar_20[2][57] , 
	\_zy_simnet_tvar_20[2][56] , \_zy_simnet_tvar_20[2][55] , 
	\_zy_simnet_tvar_20[2][54] , \_zy_simnet_tvar_20[2][53] , 
	\_zy_simnet_tvar_20[2][52] , \_zy_simnet_tvar_20[2][51] , 
	\_zy_simnet_tvar_20[2][50] , \_zy_simnet_tvar_20[2][49] , 
	\_zy_simnet_tvar_20[2][48] , \_zy_simnet_tvar_20[2][47] , 
	\_zy_simnet_tvar_20[2][46] , \_zy_simnet_tvar_20[2][45] , 
	\_zy_simnet_tvar_20[2][44] , \_zy_simnet_tvar_20[2][43] , 
	\_zy_simnet_tvar_20[2][42] , \_zy_simnet_tvar_20[2][41] , 
	\_zy_simnet_tvar_20[2][40] , \_zy_simnet_tvar_20[2][39] , 
	\_zy_simnet_tvar_20[2][38] , \_zy_simnet_tvar_20[2][37] , 
	\_zy_simnet_tvar_20[2][36] , \_zy_simnet_tvar_20[2][35] , 
	\_zy_simnet_tvar_20[2][34] , \_zy_simnet_tvar_20[2][33] , 
	\_zy_simnet_tvar_20[2][32] , \_zy_simnet_tvar_20[2][31] , 
	\_zy_simnet_tvar_20[2][30] , \_zy_simnet_tvar_20[2][29] , 
	\_zy_simnet_tvar_20[2][28] , \_zy_simnet_tvar_20[2][27] , 
	\_zy_simnet_tvar_20[2][26] , \_zy_simnet_tvar_20[2][25] , 
	\_zy_simnet_tvar_20[2][24] , \_zy_simnet_tvar_20[2][23] , 
	\_zy_simnet_tvar_20[2][22] , \_zy_simnet_tvar_20[2][21] , 
	\_zy_simnet_tvar_20[2][20] , \_zy_simnet_tvar_20[2][19] , 
	\_zy_simnet_tvar_20[2][18] , \_zy_simnet_tvar_20[2][17] , 
	\_zy_simnet_tvar_20[2][16] , \_zy_simnet_tvar_20[2][15] , 
	\_zy_simnet_tvar_20[2][14] , \_zy_simnet_tvar_20[2][13] , 
	\_zy_simnet_tvar_20[2][12] , \_zy_simnet_tvar_20[2][11] , 
	\_zy_simnet_tvar_20[2][10] , \_zy_simnet_tvar_20[2][9] , 
	\_zy_simnet_tvar_20[2][8] , \_zy_simnet_tvar_20[2][7] , 
	\_zy_simnet_tvar_20[2][6] , \_zy_simnet_tvar_20[2][5] , 
	\_zy_simnet_tvar_20[2][4] , \_zy_simnet_tvar_20[2][3] , 
	\_zy_simnet_tvar_20[2][2] , \_zy_simnet_tvar_20[2][1] , 
	\_zy_simnet_tvar_20[2][0] , \_zy_simnet_tvar_20[1][271] , 
	\_zy_simnet_tvar_20[1][270] , \_zy_simnet_tvar_20[1][269] , 
	\_zy_simnet_tvar_20[1][268] , \_zy_simnet_tvar_20[1][267] , 
	\_zy_simnet_tvar_20[1][266] , \_zy_simnet_tvar_20[1][265] , 
	\_zy_simnet_tvar_20[1][264] , \_zy_simnet_tvar_20[1][263] , 
	\_zy_simnet_tvar_20[1][262] , \_zy_simnet_tvar_20[1][261] , 
	\_zy_simnet_tvar_20[1][260] , \_zy_simnet_tvar_20[1][259] , 
	\_zy_simnet_tvar_20[1][258] , \_zy_simnet_tvar_20[1][257] , 
	\_zy_simnet_tvar_20[1][256] , \_zy_simnet_tvar_20[1][255] , 
	\_zy_simnet_tvar_20[1][254] , \_zy_simnet_tvar_20[1][253] , 
	\_zy_simnet_tvar_20[1][252] , \_zy_simnet_tvar_20[1][251] , 
	\_zy_simnet_tvar_20[1][250] , \_zy_simnet_tvar_20[1][249] , 
	\_zy_simnet_tvar_20[1][248] , \_zy_simnet_tvar_20[1][247] , 
	\_zy_simnet_tvar_20[1][246] , \_zy_simnet_tvar_20[1][245] , 
	\_zy_simnet_tvar_20[1][244] , \_zy_simnet_tvar_20[1][243] , 
	\_zy_simnet_tvar_20[1][242] , \_zy_simnet_tvar_20[1][241] , 
	\_zy_simnet_tvar_20[1][240] , \_zy_simnet_tvar_20[1][239] , 
	\_zy_simnet_tvar_20[1][238] , \_zy_simnet_tvar_20[1][237] , 
	\_zy_simnet_tvar_20[1][236] , \_zy_simnet_tvar_20[1][235] , 
	\_zy_simnet_tvar_20[1][234] , \_zy_simnet_tvar_20[1][233] , 
	\_zy_simnet_tvar_20[1][232] , \_zy_simnet_tvar_20[1][231] , 
	\_zy_simnet_tvar_20[1][230] , \_zy_simnet_tvar_20[1][229] , 
	\_zy_simnet_tvar_20[1][228] , \_zy_simnet_tvar_20[1][227] , 
	\_zy_simnet_tvar_20[1][226] , \_zy_simnet_tvar_20[1][225] , 
	\_zy_simnet_tvar_20[1][224] , \_zy_simnet_tvar_20[1][223] , 
	\_zy_simnet_tvar_20[1][222] , \_zy_simnet_tvar_20[1][221] , 
	\_zy_simnet_tvar_20[1][220] , \_zy_simnet_tvar_20[1][219] , 
	\_zy_simnet_tvar_20[1][218] , \_zy_simnet_tvar_20[1][217] , 
	\_zy_simnet_tvar_20[1][216] , \_zy_simnet_tvar_20[1][215] , 
	\_zy_simnet_tvar_20[1][214] , \_zy_simnet_tvar_20[1][213] , 
	\_zy_simnet_tvar_20[1][212] , \_zy_simnet_tvar_20[1][211] , 
	\_zy_simnet_tvar_20[1][210] , \_zy_simnet_tvar_20[1][209] , 
	\_zy_simnet_tvar_20[1][208] , \_zy_simnet_tvar_20[1][207] , 
	\_zy_simnet_tvar_20[1][206] , \_zy_simnet_tvar_20[1][205] , 
	\_zy_simnet_tvar_20[1][204] , \_zy_simnet_tvar_20[1][203] , 
	\_zy_simnet_tvar_20[1][202] , \_zy_simnet_tvar_20[1][201] , 
	\_zy_simnet_tvar_20[1][200] , \_zy_simnet_tvar_20[1][199] , 
	\_zy_simnet_tvar_20[1][198] , \_zy_simnet_tvar_20[1][197] , 
	\_zy_simnet_tvar_20[1][196] , \_zy_simnet_tvar_20[1][195] , 
	\_zy_simnet_tvar_20[1][194] , \_zy_simnet_tvar_20[1][193] , 
	\_zy_simnet_tvar_20[1][192] , \_zy_simnet_tvar_20[1][191] , 
	\_zy_simnet_tvar_20[1][190] , \_zy_simnet_tvar_20[1][189] , 
	\_zy_simnet_tvar_20[1][188] , \_zy_simnet_tvar_20[1][187] , 
	\_zy_simnet_tvar_20[1][186] , \_zy_simnet_tvar_20[1][185] , 
	\_zy_simnet_tvar_20[1][184] , \_zy_simnet_tvar_20[1][183] , 
	\_zy_simnet_tvar_20[1][182] , \_zy_simnet_tvar_20[1][181] , 
	\_zy_simnet_tvar_20[1][180] , \_zy_simnet_tvar_20[1][179] , 
	\_zy_simnet_tvar_20[1][178] , \_zy_simnet_tvar_20[1][177] , 
	\_zy_simnet_tvar_20[1][176] , \_zy_simnet_tvar_20[1][175] , 
	\_zy_simnet_tvar_20[1][174] , \_zy_simnet_tvar_20[1][173] , 
	\_zy_simnet_tvar_20[1][172] , \_zy_simnet_tvar_20[1][171] , 
	\_zy_simnet_tvar_20[1][170] , \_zy_simnet_tvar_20[1][169] , 
	\_zy_simnet_tvar_20[1][168] , \_zy_simnet_tvar_20[1][167] , 
	\_zy_simnet_tvar_20[1][166] , \_zy_simnet_tvar_20[1][165] , 
	\_zy_simnet_tvar_20[1][164] , \_zy_simnet_tvar_20[1][163] , 
	\_zy_simnet_tvar_20[1][162] , \_zy_simnet_tvar_20[1][161] , 
	\_zy_simnet_tvar_20[1][160] , \_zy_simnet_tvar_20[1][159] , 
	\_zy_simnet_tvar_20[1][158] , \_zy_simnet_tvar_20[1][157] , 
	\_zy_simnet_tvar_20[1][156] , \_zy_simnet_tvar_20[1][155] , 
	\_zy_simnet_tvar_20[1][154] , \_zy_simnet_tvar_20[1][153] , 
	\_zy_simnet_tvar_20[1][152] , \_zy_simnet_tvar_20[1][151] , 
	\_zy_simnet_tvar_20[1][150] , \_zy_simnet_tvar_20[1][149] , 
	\_zy_simnet_tvar_20[1][148] , \_zy_simnet_tvar_20[1][147] , 
	\_zy_simnet_tvar_20[1][146] , \_zy_simnet_tvar_20[1][145] , 
	\_zy_simnet_tvar_20[1][144] , \_zy_simnet_tvar_20[1][143] , 
	\_zy_simnet_tvar_20[1][142] , \_zy_simnet_tvar_20[1][141] , 
	\_zy_simnet_tvar_20[1][140] , \_zy_simnet_tvar_20[1][139] , 
	\_zy_simnet_tvar_20[1][138] , \_zy_simnet_tvar_20[1][137] , 
	\_zy_simnet_tvar_20[1][136] , \_zy_simnet_tvar_20[1][135] , 
	\_zy_simnet_tvar_20[1][134] , \_zy_simnet_tvar_20[1][133] , 
	\_zy_simnet_tvar_20[1][132] , \_zy_simnet_tvar_20[1][131] , 
	\_zy_simnet_tvar_20[1][130] , \_zy_simnet_tvar_20[1][129] , 
	\_zy_simnet_tvar_20[1][128] , \_zy_simnet_tvar_20[1][127] , 
	\_zy_simnet_tvar_20[1][126] , \_zy_simnet_tvar_20[1][125] , 
	\_zy_simnet_tvar_20[1][124] , \_zy_simnet_tvar_20[1][123] , 
	\_zy_simnet_tvar_20[1][122] , \_zy_simnet_tvar_20[1][121] , 
	\_zy_simnet_tvar_20[1][120] , \_zy_simnet_tvar_20[1][119] , 
	\_zy_simnet_tvar_20[1][118] , \_zy_simnet_tvar_20[1][117] , 
	\_zy_simnet_tvar_20[1][116] , \_zy_simnet_tvar_20[1][115] , 
	\_zy_simnet_tvar_20[1][114] , \_zy_simnet_tvar_20[1][113] , 
	\_zy_simnet_tvar_20[1][112] , \_zy_simnet_tvar_20[1][111] , 
	\_zy_simnet_tvar_20[1][110] , \_zy_simnet_tvar_20[1][109] , 
	\_zy_simnet_tvar_20[1][108] , \_zy_simnet_tvar_20[1][107] , 
	\_zy_simnet_tvar_20[1][106] , \_zy_simnet_tvar_20[1][105] , 
	\_zy_simnet_tvar_20[1][104] , \_zy_simnet_tvar_20[1][103] , 
	\_zy_simnet_tvar_20[1][102] , \_zy_simnet_tvar_20[1][101] , 
	\_zy_simnet_tvar_20[1][100] , \_zy_simnet_tvar_20[1][99] , 
	\_zy_simnet_tvar_20[1][98] , \_zy_simnet_tvar_20[1][97] , 
	\_zy_simnet_tvar_20[1][96] , \_zy_simnet_tvar_20[1][95] , 
	\_zy_simnet_tvar_20[1][94] , \_zy_simnet_tvar_20[1][93] , 
	\_zy_simnet_tvar_20[1][92] , \_zy_simnet_tvar_20[1][91] , 
	\_zy_simnet_tvar_20[1][90] , \_zy_simnet_tvar_20[1][89] , 
	\_zy_simnet_tvar_20[1][88] , \_zy_simnet_tvar_20[1][87] , 
	\_zy_simnet_tvar_20[1][86] , \_zy_simnet_tvar_20[1][85] , 
	\_zy_simnet_tvar_20[1][84] , \_zy_simnet_tvar_20[1][83] , 
	\_zy_simnet_tvar_20[1][82] , \_zy_simnet_tvar_20[1][81] , 
	\_zy_simnet_tvar_20[1][80] , \_zy_simnet_tvar_20[1][79] , 
	\_zy_simnet_tvar_20[1][78] , \_zy_simnet_tvar_20[1][77] , 
	\_zy_simnet_tvar_20[1][76] , \_zy_simnet_tvar_20[1][75] , 
	\_zy_simnet_tvar_20[1][74] , \_zy_simnet_tvar_20[1][73] , 
	\_zy_simnet_tvar_20[1][72] , \_zy_simnet_tvar_20[1][71] , 
	\_zy_simnet_tvar_20[1][70] , \_zy_simnet_tvar_20[1][69] , 
	\_zy_simnet_tvar_20[1][68] , \_zy_simnet_tvar_20[1][67] , 
	\_zy_simnet_tvar_20[1][66] , \_zy_simnet_tvar_20[1][65] , 
	\_zy_simnet_tvar_20[1][64] , \_zy_simnet_tvar_20[1][63] , 
	\_zy_simnet_tvar_20[1][62] , \_zy_simnet_tvar_20[1][61] , 
	\_zy_simnet_tvar_20[1][60] , \_zy_simnet_tvar_20[1][59] , 
	\_zy_simnet_tvar_20[1][58] , \_zy_simnet_tvar_20[1][57] , 
	\_zy_simnet_tvar_20[1][56] , \_zy_simnet_tvar_20[1][55] , 
	\_zy_simnet_tvar_20[1][54] , \_zy_simnet_tvar_20[1][53] , 
	\_zy_simnet_tvar_20[1][52] , \_zy_simnet_tvar_20[1][51] , 
	\_zy_simnet_tvar_20[1][50] , \_zy_simnet_tvar_20[1][49] , 
	\_zy_simnet_tvar_20[1][48] , \_zy_simnet_tvar_20[1][47] , 
	\_zy_simnet_tvar_20[1][46] , \_zy_simnet_tvar_20[1][45] , 
	\_zy_simnet_tvar_20[1][44] , \_zy_simnet_tvar_20[1][43] , 
	\_zy_simnet_tvar_20[1][42] , \_zy_simnet_tvar_20[1][41] , 
	\_zy_simnet_tvar_20[1][40] , \_zy_simnet_tvar_20[1][39] , 
	\_zy_simnet_tvar_20[1][38] , \_zy_simnet_tvar_20[1][37] , 
	\_zy_simnet_tvar_20[1][36] , \_zy_simnet_tvar_20[1][35] , 
	\_zy_simnet_tvar_20[1][34] , \_zy_simnet_tvar_20[1][33] , 
	\_zy_simnet_tvar_20[1][32] , \_zy_simnet_tvar_20[1][31] , 
	\_zy_simnet_tvar_20[1][30] , \_zy_simnet_tvar_20[1][29] , 
	\_zy_simnet_tvar_20[1][28] , \_zy_simnet_tvar_20[1][27] , 
	\_zy_simnet_tvar_20[1][26] , \_zy_simnet_tvar_20[1][25] , 
	\_zy_simnet_tvar_20[1][24] , \_zy_simnet_tvar_20[1][23] , 
	\_zy_simnet_tvar_20[1][22] , \_zy_simnet_tvar_20[1][21] , 
	\_zy_simnet_tvar_20[1][20] , \_zy_simnet_tvar_20[1][19] , 
	\_zy_simnet_tvar_20[1][18] , \_zy_simnet_tvar_20[1][17] , 
	\_zy_simnet_tvar_20[1][16] , \_zy_simnet_tvar_20[1][15] , 
	\_zy_simnet_tvar_20[1][14] , \_zy_simnet_tvar_20[1][13] , 
	\_zy_simnet_tvar_20[1][12] , \_zy_simnet_tvar_20[1][11] , 
	\_zy_simnet_tvar_20[1][10] , \_zy_simnet_tvar_20[1][9] , 
	\_zy_simnet_tvar_20[1][8] , \_zy_simnet_tvar_20[1][7] , 
	\_zy_simnet_tvar_20[1][6] , \_zy_simnet_tvar_20[1][5] , 
	\_zy_simnet_tvar_20[1][4] , \_zy_simnet_tvar_20[1][3] , 
	\_zy_simnet_tvar_20[1][2] , \_zy_simnet_tvar_20[1][1] , 
	\_zy_simnet_tvar_20[1][0] , \_zy_simnet_tvar_20[0][271] , 
	\_zy_simnet_tvar_20[0][270] , \_zy_simnet_tvar_20[0][269] , 
	\_zy_simnet_tvar_20[0][268] , \_zy_simnet_tvar_20[0][267] , 
	\_zy_simnet_tvar_20[0][266] , \_zy_simnet_tvar_20[0][265] , 
	\_zy_simnet_tvar_20[0][264] , \_zy_simnet_tvar_20[0][263] , 
	\_zy_simnet_tvar_20[0][262] , \_zy_simnet_tvar_20[0][261] , 
	\_zy_simnet_tvar_20[0][260] , \_zy_simnet_tvar_20[0][259] , 
	\_zy_simnet_tvar_20[0][258] , \_zy_simnet_tvar_20[0][257] , 
	\_zy_simnet_tvar_20[0][256] , \_zy_simnet_tvar_20[0][255] , 
	\_zy_simnet_tvar_20[0][254] , \_zy_simnet_tvar_20[0][253] , 
	\_zy_simnet_tvar_20[0][252] , \_zy_simnet_tvar_20[0][251] , 
	\_zy_simnet_tvar_20[0][250] , \_zy_simnet_tvar_20[0][249] , 
	\_zy_simnet_tvar_20[0][248] , \_zy_simnet_tvar_20[0][247] , 
	\_zy_simnet_tvar_20[0][246] , \_zy_simnet_tvar_20[0][245] , 
	\_zy_simnet_tvar_20[0][244] , \_zy_simnet_tvar_20[0][243] , 
	\_zy_simnet_tvar_20[0][242] , \_zy_simnet_tvar_20[0][241] , 
	\_zy_simnet_tvar_20[0][240] , \_zy_simnet_tvar_20[0][239] , 
	\_zy_simnet_tvar_20[0][238] , \_zy_simnet_tvar_20[0][237] , 
	\_zy_simnet_tvar_20[0][236] , \_zy_simnet_tvar_20[0][235] , 
	\_zy_simnet_tvar_20[0][234] , \_zy_simnet_tvar_20[0][233] , 
	\_zy_simnet_tvar_20[0][232] , \_zy_simnet_tvar_20[0][231] , 
	\_zy_simnet_tvar_20[0][230] , \_zy_simnet_tvar_20[0][229] , 
	\_zy_simnet_tvar_20[0][228] , \_zy_simnet_tvar_20[0][227] , 
	\_zy_simnet_tvar_20[0][226] , \_zy_simnet_tvar_20[0][225] , 
	\_zy_simnet_tvar_20[0][224] , \_zy_simnet_tvar_20[0][223] , 
	\_zy_simnet_tvar_20[0][222] , \_zy_simnet_tvar_20[0][221] , 
	\_zy_simnet_tvar_20[0][220] , \_zy_simnet_tvar_20[0][219] , 
	\_zy_simnet_tvar_20[0][218] , \_zy_simnet_tvar_20[0][217] , 
	\_zy_simnet_tvar_20[0][216] , \_zy_simnet_tvar_20[0][215] , 
	\_zy_simnet_tvar_20[0][214] , \_zy_simnet_tvar_20[0][213] , 
	\_zy_simnet_tvar_20[0][212] , \_zy_simnet_tvar_20[0][211] , 
	\_zy_simnet_tvar_20[0][210] , \_zy_simnet_tvar_20[0][209] , 
	\_zy_simnet_tvar_20[0][208] , \_zy_simnet_tvar_20[0][207] , 
	\_zy_simnet_tvar_20[0][206] , \_zy_simnet_tvar_20[0][205] , 
	\_zy_simnet_tvar_20[0][204] , \_zy_simnet_tvar_20[0][203] , 
	\_zy_simnet_tvar_20[0][202] , \_zy_simnet_tvar_20[0][201] , 
	\_zy_simnet_tvar_20[0][200] , \_zy_simnet_tvar_20[0][199] , 
	\_zy_simnet_tvar_20[0][198] , \_zy_simnet_tvar_20[0][197] , 
	\_zy_simnet_tvar_20[0][196] , \_zy_simnet_tvar_20[0][195] , 
	\_zy_simnet_tvar_20[0][194] , \_zy_simnet_tvar_20[0][193] , 
	\_zy_simnet_tvar_20[0][192] , \_zy_simnet_tvar_20[0][191] , 
	\_zy_simnet_tvar_20[0][190] , \_zy_simnet_tvar_20[0][189] , 
	\_zy_simnet_tvar_20[0][188] , \_zy_simnet_tvar_20[0][187] , 
	\_zy_simnet_tvar_20[0][186] , \_zy_simnet_tvar_20[0][185] , 
	\_zy_simnet_tvar_20[0][184] , \_zy_simnet_tvar_20[0][183] , 
	\_zy_simnet_tvar_20[0][182] , \_zy_simnet_tvar_20[0][181] , 
	\_zy_simnet_tvar_20[0][180] , \_zy_simnet_tvar_20[0][179] , 
	\_zy_simnet_tvar_20[0][178] , \_zy_simnet_tvar_20[0][177] , 
	\_zy_simnet_tvar_20[0][176] , \_zy_simnet_tvar_20[0][175] , 
	\_zy_simnet_tvar_20[0][174] , \_zy_simnet_tvar_20[0][173] , 
	\_zy_simnet_tvar_20[0][172] , \_zy_simnet_tvar_20[0][171] , 
	\_zy_simnet_tvar_20[0][170] , \_zy_simnet_tvar_20[0][169] , 
	\_zy_simnet_tvar_20[0][168] , \_zy_simnet_tvar_20[0][167] , 
	\_zy_simnet_tvar_20[0][166] , \_zy_simnet_tvar_20[0][165] , 
	\_zy_simnet_tvar_20[0][164] , \_zy_simnet_tvar_20[0][163] , 
	\_zy_simnet_tvar_20[0][162] , \_zy_simnet_tvar_20[0][161] , 
	\_zy_simnet_tvar_20[0][160] , \_zy_simnet_tvar_20[0][159] , 
	\_zy_simnet_tvar_20[0][158] , \_zy_simnet_tvar_20[0][157] , 
	\_zy_simnet_tvar_20[0][156] , \_zy_simnet_tvar_20[0][155] , 
	\_zy_simnet_tvar_20[0][154] , \_zy_simnet_tvar_20[0][153] , 
	\_zy_simnet_tvar_20[0][152] , \_zy_simnet_tvar_20[0][151] , 
	\_zy_simnet_tvar_20[0][150] , \_zy_simnet_tvar_20[0][149] , 
	\_zy_simnet_tvar_20[0][148] , \_zy_simnet_tvar_20[0][147] , 
	\_zy_simnet_tvar_20[0][146] , \_zy_simnet_tvar_20[0][145] , 
	\_zy_simnet_tvar_20[0][144] , \_zy_simnet_tvar_20[0][143] , 
	\_zy_simnet_tvar_20[0][142] , \_zy_simnet_tvar_20[0][141] , 
	\_zy_simnet_tvar_20[0][140] , \_zy_simnet_tvar_20[0][139] , 
	\_zy_simnet_tvar_20[0][138] , \_zy_simnet_tvar_20[0][137] , 
	\_zy_simnet_tvar_20[0][136] , \_zy_simnet_tvar_20[0][135] , 
	\_zy_simnet_tvar_20[0][134] , \_zy_simnet_tvar_20[0][133] , 
	\_zy_simnet_tvar_20[0][132] , \_zy_simnet_tvar_20[0][131] , 
	\_zy_simnet_tvar_20[0][130] , \_zy_simnet_tvar_20[0][129] , 
	\_zy_simnet_tvar_20[0][128] , \_zy_simnet_tvar_20[0][127] , 
	\_zy_simnet_tvar_20[0][126] , \_zy_simnet_tvar_20[0][125] , 
	\_zy_simnet_tvar_20[0][124] , \_zy_simnet_tvar_20[0][123] , 
	\_zy_simnet_tvar_20[0][122] , \_zy_simnet_tvar_20[0][121] , 
	\_zy_simnet_tvar_20[0][120] , \_zy_simnet_tvar_20[0][119] , 
	\_zy_simnet_tvar_20[0][118] , \_zy_simnet_tvar_20[0][117] , 
	\_zy_simnet_tvar_20[0][116] , \_zy_simnet_tvar_20[0][115] , 
	\_zy_simnet_tvar_20[0][114] , \_zy_simnet_tvar_20[0][113] , 
	\_zy_simnet_tvar_20[0][112] , \_zy_simnet_tvar_20[0][111] , 
	\_zy_simnet_tvar_20[0][110] , \_zy_simnet_tvar_20[0][109] , 
	\_zy_simnet_tvar_20[0][108] , \_zy_simnet_tvar_20[0][107] , 
	\_zy_simnet_tvar_20[0][106] , \_zy_simnet_tvar_20[0][105] , 
	\_zy_simnet_tvar_20[0][104] , \_zy_simnet_tvar_20[0][103] , 
	\_zy_simnet_tvar_20[0][102] , \_zy_simnet_tvar_20[0][101] , 
	\_zy_simnet_tvar_20[0][100] , \_zy_simnet_tvar_20[0][99] , 
	\_zy_simnet_tvar_20[0][98] , \_zy_simnet_tvar_20[0][97] , 
	\_zy_simnet_tvar_20[0][96] , \_zy_simnet_tvar_20[0][95] , 
	\_zy_simnet_tvar_20[0][94] , \_zy_simnet_tvar_20[0][93] , 
	\_zy_simnet_tvar_20[0][92] , \_zy_simnet_tvar_20[0][91] , 
	\_zy_simnet_tvar_20[0][90] , \_zy_simnet_tvar_20[0][89] , 
	\_zy_simnet_tvar_20[0][88] , \_zy_simnet_tvar_20[0][87] , 
	\_zy_simnet_tvar_20[0][86] , \_zy_simnet_tvar_20[0][85] , 
	\_zy_simnet_tvar_20[0][84] , \_zy_simnet_tvar_20[0][83] , 
	\_zy_simnet_tvar_20[0][82] , \_zy_simnet_tvar_20[0][81] , 
	\_zy_simnet_tvar_20[0][80] , \_zy_simnet_tvar_20[0][79] , 
	\_zy_simnet_tvar_20[0][78] , \_zy_simnet_tvar_20[0][77] , 
	\_zy_simnet_tvar_20[0][76] , \_zy_simnet_tvar_20[0][75] , 
	\_zy_simnet_tvar_20[0][74] , \_zy_simnet_tvar_20[0][73] , 
	\_zy_simnet_tvar_20[0][72] , \_zy_simnet_tvar_20[0][71] , 
	\_zy_simnet_tvar_20[0][70] , \_zy_simnet_tvar_20[0][69] , 
	\_zy_simnet_tvar_20[0][68] , \_zy_simnet_tvar_20[0][67] , 
	\_zy_simnet_tvar_20[0][66] , \_zy_simnet_tvar_20[0][65] , 
	\_zy_simnet_tvar_20[0][64] , \_zy_simnet_tvar_20[0][63] , 
	\_zy_simnet_tvar_20[0][62] , \_zy_simnet_tvar_20[0][61] , 
	\_zy_simnet_tvar_20[0][60] , \_zy_simnet_tvar_20[0][59] , 
	\_zy_simnet_tvar_20[0][58] , \_zy_simnet_tvar_20[0][57] , 
	\_zy_simnet_tvar_20[0][56] , \_zy_simnet_tvar_20[0][55] , 
	\_zy_simnet_tvar_20[0][54] , \_zy_simnet_tvar_20[0][53] , 
	\_zy_simnet_tvar_20[0][52] , \_zy_simnet_tvar_20[0][51] , 
	\_zy_simnet_tvar_20[0][50] , \_zy_simnet_tvar_20[0][49] , 
	\_zy_simnet_tvar_20[0][48] , \_zy_simnet_tvar_20[0][47] , 
	\_zy_simnet_tvar_20[0][46] , \_zy_simnet_tvar_20[0][45] , 
	\_zy_simnet_tvar_20[0][44] , \_zy_simnet_tvar_20[0][43] , 
	\_zy_simnet_tvar_20[0][42] , \_zy_simnet_tvar_20[0][41] , 
	\_zy_simnet_tvar_20[0][40] , \_zy_simnet_tvar_20[0][39] , 
	\_zy_simnet_tvar_20[0][38] , \_zy_simnet_tvar_20[0][37] , 
	\_zy_simnet_tvar_20[0][36] , \_zy_simnet_tvar_20[0][35] , 
	\_zy_simnet_tvar_20[0][34] , \_zy_simnet_tvar_20[0][33] , 
	\_zy_simnet_tvar_20[0][32] , \_zy_simnet_tvar_20[0][31] , 
	\_zy_simnet_tvar_20[0][30] , \_zy_simnet_tvar_20[0][29] , 
	\_zy_simnet_tvar_20[0][28] , \_zy_simnet_tvar_20[0][27] , 
	\_zy_simnet_tvar_20[0][26] , \_zy_simnet_tvar_20[0][25] , 
	\_zy_simnet_tvar_20[0][24] , \_zy_simnet_tvar_20[0][23] , 
	\_zy_simnet_tvar_20[0][22] , \_zy_simnet_tvar_20[0][21] , 
	\_zy_simnet_tvar_20[0][20] , \_zy_simnet_tvar_20[0][19] , 
	\_zy_simnet_tvar_20[0][18] , \_zy_simnet_tvar_20[0][17] , 
	\_zy_simnet_tvar_20[0][16] , \_zy_simnet_tvar_20[0][15] , 
	\_zy_simnet_tvar_20[0][14] , \_zy_simnet_tvar_20[0][13] , 
	\_zy_simnet_tvar_20[0][12] , \_zy_simnet_tvar_20[0][11] , 
	\_zy_simnet_tvar_20[0][10] , \_zy_simnet_tvar_20[0][9] , 
	\_zy_simnet_tvar_20[0][8] , \_zy_simnet_tvar_20[0][7] , 
	\_zy_simnet_tvar_20[0][6] , \_zy_simnet_tvar_20[0][5] , 
	\_zy_simnet_tvar_20[0][4] , \_zy_simnet_tvar_20[0][3] , 
	\_zy_simnet_tvar_20[0][2] , \_zy_simnet_tvar_20[0][1] , 
	\_zy_simnet_tvar_20[0][0] }, { \labels[7][271] , \labels[7][270] , 
	\labels[7][269] , \labels[7][268] , \labels[7][267] , 
	\labels[7][266] , \labels[7][265] , \labels[7][264] , 
	\labels[7][263] , \labels[7][262] , \labels[7][261] , 
	\labels[7][260] , \labels[7][259] , \labels[7][258] , 
	\labels[7][257] , \labels[7][256] , \labels[7][255] , 
	\labels[7][254] , \labels[7][253] , \labels[7][252] , 
	\labels[7][251] , \labels[7][250] , \labels[7][249] , 
	\labels[7][248] , \labels[7][247] , \labels[7][246] , 
	\labels[7][245] , \labels[7][244] , \labels[7][243] , 
	\labels[7][242] , \labels[7][241] , \labels[7][240] , 
	\labels[7][239] , \labels[7][238] , \labels[7][237] , 
	\labels[7][236] , \labels[7][235] , \labels[7][234] , 
	\labels[7][233] , \labels[7][232] , \labels[7][231] , 
	\labels[7][230] , \labels[7][229] , \labels[7][228] , 
	\labels[7][227] , \labels[7][226] , \labels[7][225] , 
	\labels[7][224] , \labels[7][223] , \labels[7][222] , 
	\labels[7][221] , \labels[7][220] , \labels[7][219] , 
	\labels[7][218] , \labels[7][217] , \labels[7][216] , 
	\labels[7][215] , \labels[7][214] , \labels[7][213] , 
	\labels[7][212] , \labels[7][211] , \labels[7][210] , 
	\labels[7][209] , \labels[7][208] , \labels[7][207] , 
	\labels[7][206] , \labels[7][205] , \labels[7][204] , 
	\labels[7][203] , \labels[7][202] , \labels[7][201] , 
	\labels[7][200] , \labels[7][199] , \labels[7][198] , 
	\labels[7][197] , \labels[7][196] , \labels[7][195] , 
	\labels[7][194] , \labels[7][193] , \labels[7][192] , 
	\labels[7][191] , \labels[7][190] , \labels[7][189] , 
	\labels[7][188] , \labels[7][187] , \labels[7][186] , 
	\labels[7][185] , \labels[7][184] , \labels[7][183] , 
	\labels[7][182] , \labels[7][181] , \labels[7][180] , 
	\labels[7][179] , \labels[7][178] , \labels[7][177] , 
	\labels[7][176] , \labels[7][175] , \labels[7][174] , 
	\labels[7][173] , \labels[7][172] , \labels[7][171] , 
	\labels[7][170] , \labels[7][169] , \labels[7][168] , 
	\labels[7][167] , \labels[7][166] , \labels[7][165] , 
	\labels[7][164] , \labels[7][163] , \labels[7][162] , 
	\labels[7][161] , \labels[7][160] , \labels[7][159] , 
	\labels[7][158] , \labels[7][157] , \labels[7][156] , 
	\labels[7][155] , \labels[7][154] , \labels[7][153] , 
	\labels[7][152] , \labels[7][151] , \labels[7][150] , 
	\labels[7][149] , \labels[7][148] , \labels[7][147] , 
	\labels[7][146] , \labels[7][145] , \labels[7][144] , 
	\labels[7][143] , \labels[7][142] , \labels[7][141] , 
	\labels[7][140] , \labels[7][139] , \labels[7][138] , 
	\labels[7][137] , \labels[7][136] , \labels[7][135] , 
	\labels[7][134] , \labels[7][133] , \labels[7][132] , 
	\labels[7][131] , \labels[7][130] , \labels[7][129] , 
	\labels[7][128] , \labels[7][127] , \labels[7][126] , 
	\labels[7][125] , \labels[7][124] , \labels[7][123] , 
	\labels[7][122] , \labels[7][121] , \labels[7][120] , 
	\labels[7][119] , \labels[7][118] , \labels[7][117] , 
	\labels[7][116] , \labels[7][115] , \labels[7][114] , 
	\labels[7][113] , \labels[7][112] , \labels[7][111] , 
	\labels[7][110] , \labels[7][109] , \labels[7][108] , 
	\labels[7][107] , \labels[7][106] , \labels[7][105] , 
	\labels[7][104] , \labels[7][103] , \labels[7][102] , 
	\labels[7][101] , \labels[7][100] , \labels[7][99] , \labels[7][98] , 
	\labels[7][97] , \labels[7][96] , \labels[7][95] , \labels[7][94] , 
	\labels[7][93] , \labels[7][92] , \labels[7][91] , \labels[7][90] , 
	\labels[7][89] , \labels[7][88] , \labels[7][87] , \labels[7][86] , 
	\labels[7][85] , \labels[7][84] , \labels[7][83] , \labels[7][82] , 
	\labels[7][81] , \labels[7][80] , \labels[7][79] , \labels[7][78] , 
	\labels[7][77] , \labels[7][76] , \labels[7][75] , \labels[7][74] , 
	\labels[7][73] , \labels[7][72] , \labels[7][71] , \labels[7][70] , 
	\labels[7][69] , \labels[7][68] , \labels[7][67] , \labels[7][66] , 
	\labels[7][65] , \labels[7][64] , \labels[7][63] , \labels[7][62] , 
	\labels[7][61] , \labels[7][60] , \labels[7][59] , \labels[7][58] , 
	\labels[7][57] , \labels[7][56] , \labels[7][55] , \labels[7][54] , 
	\labels[7][53] , \labels[7][52] , \labels[7][51] , \labels[7][50] , 
	\labels[7][49] , \labels[7][48] , \labels[7][47] , \labels[7][46] , 
	\labels[7][45] , \labels[7][44] , \labels[7][43] , \labels[7][42] , 
	\labels[7][41] , \labels[7][40] , \labels[7][39] , \labels[7][38] , 
	\labels[7][37] , \labels[7][36] , \labels[7][35] , \labels[7][34] , 
	\labels[7][33] , \labels[7][32] , \labels[7][31] , \labels[7][30] , 
	\labels[7][29] , \labels[7][28] , \labels[7][27] , \labels[7][26] , 
	\labels[7][25] , \labels[7][24] , \labels[7][23] , \labels[7][22] , 
	\labels[7][21] , \labels[7][20] , \labels[7][19] , \labels[7][18] , 
	\labels[7][17] , \labels[7][16] , \labels[7][15] , \labels[7][14] , 
	\labels[7][13] , \labels[7][12] , \labels[7][11] , \labels[7][10] , 
	\labels[7][9] , \labels[7][8] , \labels[7][7] , \labels[7][6] , 
	\labels[7][5] , \labels[7][4] , \labels[7][3] , \labels[7][2] , 
	\labels[7][1] , \labels[7][0] , \labels[6][271] , \labels[6][270] , 
	\labels[6][269] , \labels[6][268] , \labels[6][267] , 
	\labels[6][266] , \labels[6][265] , \labels[6][264] , 
	\labels[6][263] , \labels[6][262] , \labels[6][261] , 
	\labels[6][260] , \labels[6][259] , \labels[6][258] , 
	\labels[6][257] , \labels[6][256] , \labels[6][255] , 
	\labels[6][254] , \labels[6][253] , \labels[6][252] , 
	\labels[6][251] , \labels[6][250] , \labels[6][249] , 
	\labels[6][248] , \labels[6][247] , \labels[6][246] , 
	\labels[6][245] , \labels[6][244] , \labels[6][243] , 
	\labels[6][242] , \labels[6][241] , \labels[6][240] , 
	\labels[6][239] , \labels[6][238] , \labels[6][237] , 
	\labels[6][236] , \labels[6][235] , \labels[6][234] , 
	\labels[6][233] , \labels[6][232] , \labels[6][231] , 
	\labels[6][230] , \labels[6][229] , \labels[6][228] , 
	\labels[6][227] , \labels[6][226] , \labels[6][225] , 
	\labels[6][224] , \labels[6][223] , \labels[6][222] , 
	\labels[6][221] , \labels[6][220] , \labels[6][219] , 
	\labels[6][218] , \labels[6][217] , \labels[6][216] , 
	\labels[6][215] , \labels[6][214] , \labels[6][213] , 
	\labels[6][212] , \labels[6][211] , \labels[6][210] , 
	\labels[6][209] , \labels[6][208] , \labels[6][207] , 
	\labels[6][206] , \labels[6][205] , \labels[6][204] , 
	\labels[6][203] , \labels[6][202] , \labels[6][201] , 
	\labels[6][200] , \labels[6][199] , \labels[6][198] , 
	\labels[6][197] , \labels[6][196] , \labels[6][195] , 
	\labels[6][194] , \labels[6][193] , \labels[6][192] , 
	\labels[6][191] , \labels[6][190] , \labels[6][189] , 
	\labels[6][188] , \labels[6][187] , \labels[6][186] , 
	\labels[6][185] , \labels[6][184] , \labels[6][183] , 
	\labels[6][182] , \labels[6][181] , \labels[6][180] , 
	\labels[6][179] , \labels[6][178] , \labels[6][177] , 
	\labels[6][176] , \labels[6][175] , \labels[6][174] , 
	\labels[6][173] , \labels[6][172] , \labels[6][171] , 
	\labels[6][170] , \labels[6][169] , \labels[6][168] , 
	\labels[6][167] , \labels[6][166] , \labels[6][165] , 
	\labels[6][164] , \labels[6][163] , \labels[6][162] , 
	\labels[6][161] , \labels[6][160] , \labels[6][159] , 
	\labels[6][158] , \labels[6][157] , \labels[6][156] , 
	\labels[6][155] , \labels[6][154] , \labels[6][153] , 
	\labels[6][152] , \labels[6][151] , \labels[6][150] , 
	\labels[6][149] , \labels[6][148] , \labels[6][147] , 
	\labels[6][146] , \labels[6][145] , \labels[6][144] , 
	\labels[6][143] , \labels[6][142] , \labels[6][141] , 
	\labels[6][140] , \labels[6][139] , \labels[6][138] , 
	\labels[6][137] , \labels[6][136] , \labels[6][135] , 
	\labels[6][134] , \labels[6][133] , \labels[6][132] , 
	\labels[6][131] , \labels[6][130] , \labels[6][129] , 
	\labels[6][128] , \labels[6][127] , \labels[6][126] , 
	\labels[6][125] , \labels[6][124] , \labels[6][123] , 
	\labels[6][122] , \labels[6][121] , \labels[6][120] , 
	\labels[6][119] , \labels[6][118] , \labels[6][117] , 
	\labels[6][116] , \labels[6][115] , \labels[6][114] , 
	\labels[6][113] , \labels[6][112] , \labels[6][111] , 
	\labels[6][110] , \labels[6][109] , \labels[6][108] , 
	\labels[6][107] , \labels[6][106] , \labels[6][105] , 
	\labels[6][104] , \labels[6][103] , \labels[6][102] , 
	\labels[6][101] , \labels[6][100] , \labels[6][99] , \labels[6][98] , 
	\labels[6][97] , \labels[6][96] , \labels[6][95] , \labels[6][94] , 
	\labels[6][93] , \labels[6][92] , \labels[6][91] , \labels[6][90] , 
	\labels[6][89] , \labels[6][88] , \labels[6][87] , \labels[6][86] , 
	\labels[6][85] , \labels[6][84] , \labels[6][83] , \labels[6][82] , 
	\labels[6][81] , \labels[6][80] , \labels[6][79] , \labels[6][78] , 
	\labels[6][77] , \labels[6][76] , \labels[6][75] , \labels[6][74] , 
	\labels[6][73] , \labels[6][72] , \labels[6][71] , \labels[6][70] , 
	\labels[6][69] , \labels[6][68] , \labels[6][67] , \labels[6][66] , 
	\labels[6][65] , \labels[6][64] , \labels[6][63] , \labels[6][62] , 
	\labels[6][61] , \labels[6][60] , \labels[6][59] , \labels[6][58] , 
	\labels[6][57] , \labels[6][56] , \labels[6][55] , \labels[6][54] , 
	\labels[6][53] , \labels[6][52] , \labels[6][51] , \labels[6][50] , 
	\labels[6][49] , \labels[6][48] , \labels[6][47] , \labels[6][46] , 
	\labels[6][45] , \labels[6][44] , \labels[6][43] , \labels[6][42] , 
	\labels[6][41] , \labels[6][40] , \labels[6][39] , \labels[6][38] , 
	\labels[6][37] , \labels[6][36] , \labels[6][35] , \labels[6][34] , 
	\labels[6][33] , \labels[6][32] , \labels[6][31] , \labels[6][30] , 
	\labels[6][29] , \labels[6][28] , \labels[6][27] , \labels[6][26] , 
	\labels[6][25] , \labels[6][24] , \labels[6][23] , \labels[6][22] , 
	\labels[6][21] , \labels[6][20] , \labels[6][19] , \labels[6][18] , 
	\labels[6][17] , \labels[6][16] , \labels[6][15] , \labels[6][14] , 
	\labels[6][13] , \labels[6][12] , \labels[6][11] , \labels[6][10] , 
	\labels[6][9] , \labels[6][8] , \labels[6][7] , \labels[6][6] , 
	\labels[6][5] , \labels[6][4] , \labels[6][3] , \labels[6][2] , 
	\labels[6][1] , \labels[6][0] , \labels[5][271] , \labels[5][270] , 
	\labels[5][269] , \labels[5][268] , \labels[5][267] , 
	\labels[5][266] , \labels[5][265] , \labels[5][264] , 
	\labels[5][263] , \labels[5][262] , \labels[5][261] , 
	\labels[5][260] , \labels[5][259] , \labels[5][258] , 
	\labels[5][257] , \labels[5][256] , \labels[5][255] , 
	\labels[5][254] , \labels[5][253] , \labels[5][252] , 
	\labels[5][251] , \labels[5][250] , \labels[5][249] , 
	\labels[5][248] , \labels[5][247] , \labels[5][246] , 
	\labels[5][245] , \labels[5][244] , \labels[5][243] , 
	\labels[5][242] , \labels[5][241] , \labels[5][240] , 
	\labels[5][239] , \labels[5][238] , \labels[5][237] , 
	\labels[5][236] , \labels[5][235] , \labels[5][234] , 
	\labels[5][233] , \labels[5][232] , \labels[5][231] , 
	\labels[5][230] , \labels[5][229] , \labels[5][228] , 
	\labels[5][227] , \labels[5][226] , \labels[5][225] , 
	\labels[5][224] , \labels[5][223] , \labels[5][222] , 
	\labels[5][221] , \labels[5][220] , \labels[5][219] , 
	\labels[5][218] , \labels[5][217] , \labels[5][216] , 
	\labels[5][215] , \labels[5][214] , \labels[5][213] , 
	\labels[5][212] , \labels[5][211] , \labels[5][210] , 
	\labels[5][209] , \labels[5][208] , \labels[5][207] , 
	\labels[5][206] , \labels[5][205] , \labels[5][204] , 
	\labels[5][203] , \labels[5][202] , \labels[5][201] , 
	\labels[5][200] , \labels[5][199] , \labels[5][198] , 
	\labels[5][197] , \labels[5][196] , \labels[5][195] , 
	\labels[5][194] , \labels[5][193] , \labels[5][192] , 
	\labels[5][191] , \labels[5][190] , \labels[5][189] , 
	\labels[5][188] , \labels[5][187] , \labels[5][186] , 
	\labels[5][185] , \labels[5][184] , \labels[5][183] , 
	\labels[5][182] , \labels[5][181] , \labels[5][180] , 
	\labels[5][179] , \labels[5][178] , \labels[5][177] , 
	\labels[5][176] , \labels[5][175] , \labels[5][174] , 
	\labels[5][173] , \labels[5][172] , \labels[5][171] , 
	\labels[5][170] , \labels[5][169] , \labels[5][168] , 
	\labels[5][167] , \labels[5][166] , \labels[5][165] , 
	\labels[5][164] , \labels[5][163] , \labels[5][162] , 
	\labels[5][161] , \labels[5][160] , \labels[5][159] , 
	\labels[5][158] , \labels[5][157] , \labels[5][156] , 
	\labels[5][155] , \labels[5][154] , \labels[5][153] , 
	\labels[5][152] , \labels[5][151] , \labels[5][150] , 
	\labels[5][149] , \labels[5][148] , \labels[5][147] , 
	\labels[5][146] , \labels[5][145] , \labels[5][144] , 
	\labels[5][143] , \labels[5][142] , \labels[5][141] , 
	\labels[5][140] , \labels[5][139] , \labels[5][138] , 
	\labels[5][137] , \labels[5][136] , \labels[5][135] , 
	\labels[5][134] , \labels[5][133] , \labels[5][132] , 
	\labels[5][131] , \labels[5][130] , \labels[5][129] , 
	\labels[5][128] , \labels[5][127] , \labels[5][126] , 
	\labels[5][125] , \labels[5][124] , \labels[5][123] , 
	\labels[5][122] , \labels[5][121] , \labels[5][120] , 
	\labels[5][119] , \labels[5][118] , \labels[5][117] , 
	\labels[5][116] , \labels[5][115] , \labels[5][114] , 
	\labels[5][113] , \labels[5][112] , \labels[5][111] , 
	\labels[5][110] , \labels[5][109] , \labels[5][108] , 
	\labels[5][107] , \labels[5][106] , \labels[5][105] , 
	\labels[5][104] , \labels[5][103] , \labels[5][102] , 
	\labels[5][101] , \labels[5][100] , \labels[5][99] , \labels[5][98] , 
	\labels[5][97] , \labels[5][96] , \labels[5][95] , \labels[5][94] , 
	\labels[5][93] , \labels[5][92] , \labels[5][91] , \labels[5][90] , 
	\labels[5][89] , \labels[5][88] , \labels[5][87] , \labels[5][86] , 
	\labels[5][85] , \labels[5][84] , \labels[5][83] , \labels[5][82] , 
	\labels[5][81] , \labels[5][80] , \labels[5][79] , \labels[5][78] , 
	\labels[5][77] , \labels[5][76] , \labels[5][75] , \labels[5][74] , 
	\labels[5][73] , \labels[5][72] , \labels[5][71] , \labels[5][70] , 
	\labels[5][69] , \labels[5][68] , \labels[5][67] , \labels[5][66] , 
	\labels[5][65] , \labels[5][64] , \labels[5][63] , \labels[5][62] , 
	\labels[5][61] , \labels[5][60] , \labels[5][59] , \labels[5][58] , 
	\labels[5][57] , \labels[5][56] , \labels[5][55] , \labels[5][54] , 
	\labels[5][53] , \labels[5][52] , \labels[5][51] , \labels[5][50] , 
	\labels[5][49] , \labels[5][48] , \labels[5][47] , \labels[5][46] , 
	\labels[5][45] , \labels[5][44] , \labels[5][43] , \labels[5][42] , 
	\labels[5][41] , \labels[5][40] , \labels[5][39] , \labels[5][38] , 
	\labels[5][37] , \labels[5][36] , \labels[5][35] , \labels[5][34] , 
	\labels[5][33] , \labels[5][32] , \labels[5][31] , \labels[5][30] , 
	\labels[5][29] , \labels[5][28] , \labels[5][27] , \labels[5][26] , 
	\labels[5][25] , \labels[5][24] , \labels[5][23] , \labels[5][22] , 
	\labels[5][21] , \labels[5][20] , \labels[5][19] , \labels[5][18] , 
	\labels[5][17] , \labels[5][16] , \labels[5][15] , \labels[5][14] , 
	\labels[5][13] , \labels[5][12] , \labels[5][11] , \labels[5][10] , 
	\labels[5][9] , \labels[5][8] , \labels[5][7] , \labels[5][6] , 
	\labels[5][5] , \labels[5][4] , \labels[5][3] , \labels[5][2] , 
	\labels[5][1] , \labels[5][0] , \labels[4][271] , \labels[4][270] , 
	\labels[4][269] , \labels[4][268] , \labels[4][267] , 
	\labels[4][266] , \labels[4][265] , \labels[4][264] , 
	\labels[4][263] , \labels[4][262] , \labels[4][261] , 
	\labels[4][260] , \labels[4][259] , \labels[4][258] , 
	\labels[4][257] , \labels[4][256] , \labels[4][255] , 
	\labels[4][254] , \labels[4][253] , \labels[4][252] , 
	\labels[4][251] , \labels[4][250] , \labels[4][249] , 
	\labels[4][248] , \labels[4][247] , \labels[4][246] , 
	\labels[4][245] , \labels[4][244] , \labels[4][243] , 
	\labels[4][242] , \labels[4][241] , \labels[4][240] , 
	\labels[4][239] , \labels[4][238] , \labels[4][237] , 
	\labels[4][236] , \labels[4][235] , \labels[4][234] , 
	\labels[4][233] , \labels[4][232] , \labels[4][231] , 
	\labels[4][230] , \labels[4][229] , \labels[4][228] , 
	\labels[4][227] , \labels[4][226] , \labels[4][225] , 
	\labels[4][224] , \labels[4][223] , \labels[4][222] , 
	\labels[4][221] , \labels[4][220] , \labels[4][219] , 
	\labels[4][218] , \labels[4][217] , \labels[4][216] , 
	\labels[4][215] , \labels[4][214] , \labels[4][213] , 
	\labels[4][212] , \labels[4][211] , \labels[4][210] , 
	\labels[4][209] , \labels[4][208] , \labels[4][207] , 
	\labels[4][206] , \labels[4][205] , \labels[4][204] , 
	\labels[4][203] , \labels[4][202] , \labels[4][201] , 
	\labels[4][200] , \labels[4][199] , \labels[4][198] , 
	\labels[4][197] , \labels[4][196] , \labels[4][195] , 
	\labels[4][194] , \labels[4][193] , \labels[4][192] , 
	\labels[4][191] , \labels[4][190] , \labels[4][189] , 
	\labels[4][188] , \labels[4][187] , \labels[4][186] , 
	\labels[4][185] , \labels[4][184] , \labels[4][183] , 
	\labels[4][182] , \labels[4][181] , \labels[4][180] , 
	\labels[4][179] , \labels[4][178] , \labels[4][177] , 
	\labels[4][176] , \labels[4][175] , \labels[4][174] , 
	\labels[4][173] , \labels[4][172] , \labels[4][171] , 
	\labels[4][170] , \labels[4][169] , \labels[4][168] , 
	\labels[4][167] , \labels[4][166] , \labels[4][165] , 
	\labels[4][164] , \labels[4][163] , \labels[4][162] , 
	\labels[4][161] , \labels[4][160] , \labels[4][159] , 
	\labels[4][158] , \labels[4][157] , \labels[4][156] , 
	\labels[4][155] , \labels[4][154] , \labels[4][153] , 
	\labels[4][152] , \labels[4][151] , \labels[4][150] , 
	\labels[4][149] , \labels[4][148] , \labels[4][147] , 
	\labels[4][146] , \labels[4][145] , \labels[4][144] , 
	\labels[4][143] , \labels[4][142] , \labels[4][141] , 
	\labels[4][140] , \labels[4][139] , \labels[4][138] , 
	\labels[4][137] , \labels[4][136] , \labels[4][135] , 
	\labels[4][134] , \labels[4][133] , \labels[4][132] , 
	\labels[4][131] , \labels[4][130] , \labels[4][129] , 
	\labels[4][128] , \labels[4][127] , \labels[4][126] , 
	\labels[4][125] , \labels[4][124] , \labels[4][123] , 
	\labels[4][122] , \labels[4][121] , \labels[4][120] , 
	\labels[4][119] , \labels[4][118] , \labels[4][117] , 
	\labels[4][116] , \labels[4][115] , \labels[4][114] , 
	\labels[4][113] , \labels[4][112] , \labels[4][111] , 
	\labels[4][110] , \labels[4][109] , \labels[4][108] , 
	\labels[4][107] , \labels[4][106] , \labels[4][105] , 
	\labels[4][104] , \labels[4][103] , \labels[4][102] , 
	\labels[4][101] , \labels[4][100] , \labels[4][99] , \labels[4][98] , 
	\labels[4][97] , \labels[4][96] , \labels[4][95] , \labels[4][94] , 
	\labels[4][93] , \labels[4][92] , \labels[4][91] , \labels[4][90] , 
	\labels[4][89] , \labels[4][88] , \labels[4][87] , \labels[4][86] , 
	\labels[4][85] , \labels[4][84] , \labels[4][83] , \labels[4][82] , 
	\labels[4][81] , \labels[4][80] , \labels[4][79] , \labels[4][78] , 
	\labels[4][77] , \labels[4][76] , \labels[4][75] , \labels[4][74] , 
	\labels[4][73] , \labels[4][72] , \labels[4][71] , \labels[4][70] , 
	\labels[4][69] , \labels[4][68] , \labels[4][67] , \labels[4][66] , 
	\labels[4][65] , \labels[4][64] , \labels[4][63] , \labels[4][62] , 
	\labels[4][61] , \labels[4][60] , \labels[4][59] , \labels[4][58] , 
	\labels[4][57] , \labels[4][56] , \labels[4][55] , \labels[4][54] , 
	\labels[4][53] , \labels[4][52] , \labels[4][51] , \labels[4][50] , 
	\labels[4][49] , \labels[4][48] , \labels[4][47] , \labels[4][46] , 
	\labels[4][45] , \labels[4][44] , \labels[4][43] , \labels[4][42] , 
	\labels[4][41] , \labels[4][40] , \labels[4][39] , \labels[4][38] , 
	\labels[4][37] , \labels[4][36] , \labels[4][35] , \labels[4][34] , 
	\labels[4][33] , \labels[4][32] , \labels[4][31] , \labels[4][30] , 
	\labels[4][29] , \labels[4][28] , \labels[4][27] , \labels[4][26] , 
	\labels[4][25] , \labels[4][24] , \labels[4][23] , \labels[4][22] , 
	\labels[4][21] , \labels[4][20] , \labels[4][19] , \labels[4][18] , 
	\labels[4][17] , \labels[4][16] , \labels[4][15] , \labels[4][14] , 
	\labels[4][13] , \labels[4][12] , \labels[4][11] , \labels[4][10] , 
	\labels[4][9] , \labels[4][8] , \labels[4][7] , \labels[4][6] , 
	\labels[4][5] , \labels[4][4] , \labels[4][3] , \labels[4][2] , 
	\labels[4][1] , \labels[4][0] , \labels[3][271] , \labels[3][270] , 
	\labels[3][269] , \labels[3][268] , \labels[3][267] , 
	\labels[3][266] , \labels[3][265] , \labels[3][264] , 
	\labels[3][263] , \labels[3][262] , \labels[3][261] , 
	\labels[3][260] , \labels[3][259] , \labels[3][258] , 
	\labels[3][257] , \labels[3][256] , \labels[3][255] , 
	\labels[3][254] , \labels[3][253] , \labels[3][252] , 
	\labels[3][251] , \labels[3][250] , \labels[3][249] , 
	\labels[3][248] , \labels[3][247] , \labels[3][246] , 
	\labels[3][245] , \labels[3][244] , \labels[3][243] , 
	\labels[3][242] , \labels[3][241] , \labels[3][240] , 
	\labels[3][239] , \labels[3][238] , \labels[3][237] , 
	\labels[3][236] , \labels[3][235] , \labels[3][234] , 
	\labels[3][233] , \labels[3][232] , \labels[3][231] , 
	\labels[3][230] , \labels[3][229] , \labels[3][228] , 
	\labels[3][227] , \labels[3][226] , \labels[3][225] , 
	\labels[3][224] , \labels[3][223] , \labels[3][222] , 
	\labels[3][221] , \labels[3][220] , \labels[3][219] , 
	\labels[3][218] , \labels[3][217] , \labels[3][216] , 
	\labels[3][215] , \labels[3][214] , \labels[3][213] , 
	\labels[3][212] , \labels[3][211] , \labels[3][210] , 
	\labels[3][209] , \labels[3][208] , \labels[3][207] , 
	\labels[3][206] , \labels[3][205] , \labels[3][204] , 
	\labels[3][203] , \labels[3][202] , \labels[3][201] , 
	\labels[3][200] , \labels[3][199] , \labels[3][198] , 
	\labels[3][197] , \labels[3][196] , \labels[3][195] , 
	\labels[3][194] , \labels[3][193] , \labels[3][192] , 
	\labels[3][191] , \labels[3][190] , \labels[3][189] , 
	\labels[3][188] , \labels[3][187] , \labels[3][186] , 
	\labels[3][185] , \labels[3][184] , \labels[3][183] , 
	\labels[3][182] , \labels[3][181] , \labels[3][180] , 
	\labels[3][179] , \labels[3][178] , \labels[3][177] , 
	\labels[3][176] , \labels[3][175] , \labels[3][174] , 
	\labels[3][173] , \labels[3][172] , \labels[3][171] , 
	\labels[3][170] , \labels[3][169] , \labels[3][168] , 
	\labels[3][167] , \labels[3][166] , \labels[3][165] , 
	\labels[3][164] , \labels[3][163] , \labels[3][162] , 
	\labels[3][161] , \labels[3][160] , \labels[3][159] , 
	\labels[3][158] , \labels[3][157] , \labels[3][156] , 
	\labels[3][155] , \labels[3][154] , \labels[3][153] , 
	\labels[3][152] , \labels[3][151] , \labels[3][150] , 
	\labels[3][149] , \labels[3][148] , \labels[3][147] , 
	\labels[3][146] , \labels[3][145] , \labels[3][144] , 
	\labels[3][143] , \labels[3][142] , \labels[3][141] , 
	\labels[3][140] , \labels[3][139] , \labels[3][138] , 
	\labels[3][137] , \labels[3][136] , \labels[3][135] , 
	\labels[3][134] , \labels[3][133] , \labels[3][132] , 
	\labels[3][131] , \labels[3][130] , \labels[3][129] , 
	\labels[3][128] , \labels[3][127] , \labels[3][126] , 
	\labels[3][125] , \labels[3][124] , \labels[3][123] , 
	\labels[3][122] , \labels[3][121] , \labels[3][120] , 
	\labels[3][119] , \labels[3][118] , \labels[3][117] , 
	\labels[3][116] , \labels[3][115] , \labels[3][114] , 
	\labels[3][113] , \labels[3][112] , \labels[3][111] , 
	\labels[3][110] , \labels[3][109] , \labels[3][108] , 
	\labels[3][107] , \labels[3][106] , \labels[3][105] , 
	\labels[3][104] , \labels[3][103] , \labels[3][102] , 
	\labels[3][101] , \labels[3][100] , \labels[3][99] , \labels[3][98] , 
	\labels[3][97] , \labels[3][96] , \labels[3][95] , \labels[3][94] , 
	\labels[3][93] , \labels[3][92] , \labels[3][91] , \labels[3][90] , 
	\labels[3][89] , \labels[3][88] , \labels[3][87] , \labels[3][86] , 
	\labels[3][85] , \labels[3][84] , \labels[3][83] , \labels[3][82] , 
	\labels[3][81] , \labels[3][80] , \labels[3][79] , \labels[3][78] , 
	\labels[3][77] , \labels[3][76] , \labels[3][75] , \labels[3][74] , 
	\labels[3][73] , \labels[3][72] , \labels[3][71] , \labels[3][70] , 
	\labels[3][69] , \labels[3][68] , \labels[3][67] , \labels[3][66] , 
	\labels[3][65] , \labels[3][64] , \labels[3][63] , \labels[3][62] , 
	\labels[3][61] , \labels[3][60] , \labels[3][59] , \labels[3][58] , 
	\labels[3][57] , \labels[3][56] , \labels[3][55] , \labels[3][54] , 
	\labels[3][53] , \labels[3][52] , \labels[3][51] , \labels[3][50] , 
	\labels[3][49] , \labels[3][48] , \labels[3][47] , \labels[3][46] , 
	\labels[3][45] , \labels[3][44] , \labels[3][43] , \labels[3][42] , 
	\labels[3][41] , \labels[3][40] , \labels[3][39] , \labels[3][38] , 
	\labels[3][37] , \labels[3][36] , \labels[3][35] , \labels[3][34] , 
	\labels[3][33] , \labels[3][32] , \labels[3][31] , \labels[3][30] , 
	\labels[3][29] , \labels[3][28] , \labels[3][27] , \labels[3][26] , 
	\labels[3][25] , \labels[3][24] , \labels[3][23] , \labels[3][22] , 
	\labels[3][21] , \labels[3][20] , \labels[3][19] , \labels[3][18] , 
	\labels[3][17] , \labels[3][16] , \labels[3][15] , \labels[3][14] , 
	\labels[3][13] , \labels[3][12] , \labels[3][11] , \labels[3][10] , 
	\labels[3][9] , \labels[3][8] , \labels[3][7] , \labels[3][6] , 
	\labels[3][5] , \labels[3][4] , \labels[3][3] , \labels[3][2] , 
	\labels[3][1] , \labels[3][0] , \labels[2][271] , \labels[2][270] , 
	\labels[2][269] , \labels[2][268] , \labels[2][267] , 
	\labels[2][266] , \labels[2][265] , \labels[2][264] , 
	\labels[2][263] , \labels[2][262] , \labels[2][261] , 
	\labels[2][260] , \labels[2][259] , \labels[2][258] , 
	\labels[2][257] , \labels[2][256] , \labels[2][255] , 
	\labels[2][254] , \labels[2][253] , \labels[2][252] , 
	\labels[2][251] , \labels[2][250] , \labels[2][249] , 
	\labels[2][248] , \labels[2][247] , \labels[2][246] , 
	\labels[2][245] , \labels[2][244] , \labels[2][243] , 
	\labels[2][242] , \labels[2][241] , \labels[2][240] , 
	\labels[2][239] , \labels[2][238] , \labels[2][237] , 
	\labels[2][236] , \labels[2][235] , \labels[2][234] , 
	\labels[2][233] , \labels[2][232] , \labels[2][231] , 
	\labels[2][230] , \labels[2][229] , \labels[2][228] , 
	\labels[2][227] , \labels[2][226] , \labels[2][225] , 
	\labels[2][224] , \labels[2][223] , \labels[2][222] , 
	\labels[2][221] , \labels[2][220] , \labels[2][219] , 
	\labels[2][218] , \labels[2][217] , \labels[2][216] , 
	\labels[2][215] , \labels[2][214] , \labels[2][213] , 
	\labels[2][212] , \labels[2][211] , \labels[2][210] , 
	\labels[2][209] , \labels[2][208] , \labels[2][207] , 
	\labels[2][206] , \labels[2][205] , \labels[2][204] , 
	\labels[2][203] , \labels[2][202] , \labels[2][201] , 
	\labels[2][200] , \labels[2][199] , \labels[2][198] , 
	\labels[2][197] , \labels[2][196] , \labels[2][195] , 
	\labels[2][194] , \labels[2][193] , \labels[2][192] , 
	\labels[2][191] , \labels[2][190] , \labels[2][189] , 
	\labels[2][188] , \labels[2][187] , \labels[2][186] , 
	\labels[2][185] , \labels[2][184] , \labels[2][183] , 
	\labels[2][182] , \labels[2][181] , \labels[2][180] , 
	\labels[2][179] , \labels[2][178] , \labels[2][177] , 
	\labels[2][176] , \labels[2][175] , \labels[2][174] , 
	\labels[2][173] , \labels[2][172] , \labels[2][171] , 
	\labels[2][170] , \labels[2][169] , \labels[2][168] , 
	\labels[2][167] , \labels[2][166] , \labels[2][165] , 
	\labels[2][164] , \labels[2][163] , \labels[2][162] , 
	\labels[2][161] , \labels[2][160] , \labels[2][159] , 
	\labels[2][158] , \labels[2][157] , \labels[2][156] , 
	\labels[2][155] , \labels[2][154] , \labels[2][153] , 
	\labels[2][152] , \labels[2][151] , \labels[2][150] , 
	\labels[2][149] , \labels[2][148] , \labels[2][147] , 
	\labels[2][146] , \labels[2][145] , \labels[2][144] , 
	\labels[2][143] , \labels[2][142] , \labels[2][141] , 
	\labels[2][140] , \labels[2][139] , \labels[2][138] , 
	\labels[2][137] , \labels[2][136] , \labels[2][135] , 
	\labels[2][134] , \labels[2][133] , \labels[2][132] , 
	\labels[2][131] , \labels[2][130] , \labels[2][129] , 
	\labels[2][128] , \labels[2][127] , \labels[2][126] , 
	\labels[2][125] , \labels[2][124] , \labels[2][123] , 
	\labels[2][122] , \labels[2][121] , \labels[2][120] , 
	\labels[2][119] , \labels[2][118] , \labels[2][117] , 
	\labels[2][116] , \labels[2][115] , \labels[2][114] , 
	\labels[2][113] , \labels[2][112] , \labels[2][111] , 
	\labels[2][110] , \labels[2][109] , \labels[2][108] , 
	\labels[2][107] , \labels[2][106] , \labels[2][105] , 
	\labels[2][104] , \labels[2][103] , \labels[2][102] , 
	\labels[2][101] , \labels[2][100] , \labels[2][99] , \labels[2][98] , 
	\labels[2][97] , \labels[2][96] , \labels[2][95] , \labels[2][94] , 
	\labels[2][93] , \labels[2][92] , \labels[2][91] , \labels[2][90] , 
	\labels[2][89] , \labels[2][88] , \labels[2][87] , \labels[2][86] , 
	\labels[2][85] , \labels[2][84] , \labels[2][83] , \labels[2][82] , 
	\labels[2][81] , \labels[2][80] , \labels[2][79] , \labels[2][78] , 
	\labels[2][77] , \labels[2][76] , \labels[2][75] , \labels[2][74] , 
	\labels[2][73] , \labels[2][72] , \labels[2][71] , \labels[2][70] , 
	\labels[2][69] , \labels[2][68] , \labels[2][67] , \labels[2][66] , 
	\labels[2][65] , \labels[2][64] , \labels[2][63] , \labels[2][62] , 
	\labels[2][61] , \labels[2][60] , \labels[2][59] , \labels[2][58] , 
	\labels[2][57] , \labels[2][56] , \labels[2][55] , \labels[2][54] , 
	\labels[2][53] , \labels[2][52] , \labels[2][51] , \labels[2][50] , 
	\labels[2][49] , \labels[2][48] , \labels[2][47] , \labels[2][46] , 
	\labels[2][45] , \labels[2][44] , \labels[2][43] , \labels[2][42] , 
	\labels[2][41] , \labels[2][40] , \labels[2][39] , \labels[2][38] , 
	\labels[2][37] , \labels[2][36] , \labels[2][35] , \labels[2][34] , 
	\labels[2][33] , \labels[2][32] , \labels[2][31] , \labels[2][30] , 
	\labels[2][29] , \labels[2][28] , \labels[2][27] , \labels[2][26] , 
	\labels[2][25] , \labels[2][24] , \labels[2][23] , \labels[2][22] , 
	\labels[2][21] , \labels[2][20] , \labels[2][19] , \labels[2][18] , 
	\labels[2][17] , \labels[2][16] , \labels[2][15] , \labels[2][14] , 
	\labels[2][13] , \labels[2][12] , \labels[2][11] , \labels[2][10] , 
	\labels[2][9] , \labels[2][8] , \labels[2][7] , \labels[2][6] , 
	\labels[2][5] , \labels[2][4] , \labels[2][3] , \labels[2][2] , 
	\labels[2][1] , \labels[2][0] , \labels[1][271] , \labels[1][270] , 
	\labels[1][269] , \labels[1][268] , \labels[1][267] , 
	\labels[1][266] , \labels[1][265] , \labels[1][264] , 
	\labels[1][263] , \labels[1][262] , \labels[1][261] , 
	\labels[1][260] , \labels[1][259] , \labels[1][258] , 
	\labels[1][257] , \labels[1][256] , \labels[1][255] , 
	\labels[1][254] , \labels[1][253] , \labels[1][252] , 
	\labels[1][251] , \labels[1][250] , \labels[1][249] , 
	\labels[1][248] , \labels[1][247] , \labels[1][246] , 
	\labels[1][245] , \labels[1][244] , \labels[1][243] , 
	\labels[1][242] , \labels[1][241] , \labels[1][240] , 
	\labels[1][239] , \labels[1][238] , \labels[1][237] , 
	\labels[1][236] , \labels[1][235] , \labels[1][234] , 
	\labels[1][233] , \labels[1][232] , \labels[1][231] , 
	\labels[1][230] , \labels[1][229] , \labels[1][228] , 
	\labels[1][227] , \labels[1][226] , \labels[1][225] , 
	\labels[1][224] , \labels[1][223] , \labels[1][222] , 
	\labels[1][221] , \labels[1][220] , \labels[1][219] , 
	\labels[1][218] , \labels[1][217] , \labels[1][216] , 
	\labels[1][215] , \labels[1][214] , \labels[1][213] , 
	\labels[1][212] , \labels[1][211] , \labels[1][210] , 
	\labels[1][209] , \labels[1][208] , \labels[1][207] , 
	\labels[1][206] , \labels[1][205] , \labels[1][204] , 
	\labels[1][203] , \labels[1][202] , \labels[1][201] , 
	\labels[1][200] , \labels[1][199] , \labels[1][198] , 
	\labels[1][197] , \labels[1][196] , \labels[1][195] , 
	\labels[1][194] , \labels[1][193] , \labels[1][192] , 
	\labels[1][191] , \labels[1][190] , \labels[1][189] , 
	\labels[1][188] , \labels[1][187] , \labels[1][186] , 
	\labels[1][185] , \labels[1][184] , \labels[1][183] , 
	\labels[1][182] , \labels[1][181] , \labels[1][180] , 
	\labels[1][179] , \labels[1][178] , \labels[1][177] , 
	\labels[1][176] , \labels[1][175] , \labels[1][174] , 
	\labels[1][173] , \labels[1][172] , \labels[1][171] , 
	\labels[1][170] , \labels[1][169] , \labels[1][168] , 
	\labels[1][167] , \labels[1][166] , \labels[1][165] , 
	\labels[1][164] , \labels[1][163] , \labels[1][162] , 
	\labels[1][161] , \labels[1][160] , \labels[1][159] , 
	\labels[1][158] , \labels[1][157] , \labels[1][156] , 
	\labels[1][155] , \labels[1][154] , \labels[1][153] , 
	\labels[1][152] , \labels[1][151] , \labels[1][150] , 
	\labels[1][149] , \labels[1][148] , \labels[1][147] , 
	\labels[1][146] , \labels[1][145] , \labels[1][144] , 
	\labels[1][143] , \labels[1][142] , \labels[1][141] , 
	\labels[1][140] , \labels[1][139] , \labels[1][138] , 
	\labels[1][137] , \labels[1][136] , \labels[1][135] , 
	\labels[1][134] , \labels[1][133] , \labels[1][132] , 
	\labels[1][131] , \labels[1][130] , \labels[1][129] , 
	\labels[1][128] , \labels[1][127] , \labels[1][126] , 
	\labels[1][125] , \labels[1][124] , \labels[1][123] , 
	\labels[1][122] , \labels[1][121] , \labels[1][120] , 
	\labels[1][119] , \labels[1][118] , \labels[1][117] , 
	\labels[1][116] , \labels[1][115] , \labels[1][114] , 
	\labels[1][113] , \labels[1][112] , \labels[1][111] , 
	\labels[1][110] , \labels[1][109] , \labels[1][108] , 
	\labels[1][107] , \labels[1][106] , \labels[1][105] , 
	\labels[1][104] , \labels[1][103] , \labels[1][102] , 
	\labels[1][101] , \labels[1][100] , \labels[1][99] , \labels[1][98] , 
	\labels[1][97] , \labels[1][96] , \labels[1][95] , \labels[1][94] , 
	\labels[1][93] , \labels[1][92] , \labels[1][91] , \labels[1][90] , 
	\labels[1][89] , \labels[1][88] , \labels[1][87] , \labels[1][86] , 
	\labels[1][85] , \labels[1][84] , \labels[1][83] , \labels[1][82] , 
	\labels[1][81] , \labels[1][80] , \labels[1][79] , \labels[1][78] , 
	\labels[1][77] , \labels[1][76] , \labels[1][75] , \labels[1][74] , 
	\labels[1][73] , \labels[1][72] , \labels[1][71] , \labels[1][70] , 
	\labels[1][69] , \labels[1][68] , \labels[1][67] , \labels[1][66] , 
	\labels[1][65] , \labels[1][64] , \labels[1][63] , \labels[1][62] , 
	\labels[1][61] , \labels[1][60] , \labels[1][59] , \labels[1][58] , 
	\labels[1][57] , \labels[1][56] , \labels[1][55] , \labels[1][54] , 
	\labels[1][53] , \labels[1][52] , \labels[1][51] , \labels[1][50] , 
	\labels[1][49] , \labels[1][48] , \labels[1][47] , \labels[1][46] , 
	\labels[1][45] , \labels[1][44] , \labels[1][43] , \labels[1][42] , 
	\labels[1][41] , \labels[1][40] , \labels[1][39] , \labels[1][38] , 
	\labels[1][37] , \labels[1][36] , \labels[1][35] , \labels[1][34] , 
	\labels[1][33] , \labels[1][32] , \labels[1][31] , \labels[1][30] , 
	\labels[1][29] , \labels[1][28] , \labels[1][27] , \labels[1][26] , 
	\labels[1][25] , \labels[1][24] , \labels[1][23] , \labels[1][22] , 
	\labels[1][21] , \labels[1][20] , \labels[1][19] , \labels[1][18] , 
	\labels[1][17] , \labels[1][16] , \labels[1][15] , \labels[1][14] , 
	\labels[1][13] , \labels[1][12] , \labels[1][11] , \labels[1][10] , 
	\labels[1][9] , \labels[1][8] , \labels[1][7] , \labels[1][6] , 
	\labels[1][5] , \labels[1][4] , \labels[1][3] , \labels[1][2] , 
	\labels[1][1] , \labels[1][0] , \labels[0][271] , \labels[0][270] , 
	\labels[0][269] , \labels[0][268] , \labels[0][267] , 
	\labels[0][266] , \labels[0][265] , \labels[0][264] , 
	\labels[0][263] , \labels[0][262] , \labels[0][261] , 
	\labels[0][260] , \labels[0][259] , \labels[0][258] , 
	\labels[0][257] , \labels[0][256] , \labels[0][255] , 
	\labels[0][254] , \labels[0][253] , \labels[0][252] , 
	\labels[0][251] , \labels[0][250] , \labels[0][249] , 
	\labels[0][248] , \labels[0][247] , \labels[0][246] , 
	\labels[0][245] , \labels[0][244] , \labels[0][243] , 
	\labels[0][242] , \labels[0][241] , \labels[0][240] , 
	\labels[0][239] , \labels[0][238] , \labels[0][237] , 
	\labels[0][236] , \labels[0][235] , \labels[0][234] , 
	\labels[0][233] , \labels[0][232] , \labels[0][231] , 
	\labels[0][230] , \labels[0][229] , \labels[0][228] , 
	\labels[0][227] , \labels[0][226] , \labels[0][225] , 
	\labels[0][224] , \labels[0][223] , \labels[0][222] , 
	\labels[0][221] , \labels[0][220] , \labels[0][219] , 
	\labels[0][218] , \labels[0][217] , \labels[0][216] , 
	\labels[0][215] , \labels[0][214] , \labels[0][213] , 
	\labels[0][212] , \labels[0][211] , \labels[0][210] , 
	\labels[0][209] , \labels[0][208] , \labels[0][207] , 
	\labels[0][206] , \labels[0][205] , \labels[0][204] , 
	\labels[0][203] , \labels[0][202] , \labels[0][201] , 
	\labels[0][200] , \labels[0][199] , \labels[0][198] , 
	\labels[0][197] , \labels[0][196] , \labels[0][195] , 
	\labels[0][194] , \labels[0][193] , \labels[0][192] , 
	\labels[0][191] , \labels[0][190] , \labels[0][189] , 
	\labels[0][188] , \labels[0][187] , \labels[0][186] , 
	\labels[0][185] , \labels[0][184] , \labels[0][183] , 
	\labels[0][182] , \labels[0][181] , \labels[0][180] , 
	\labels[0][179] , \labels[0][178] , \labels[0][177] , 
	\labels[0][176] , \labels[0][175] , \labels[0][174] , 
	\labels[0][173] , \labels[0][172] , \labels[0][171] , 
	\labels[0][170] , \labels[0][169] , \labels[0][168] , 
	\labels[0][167] , \labels[0][166] , \labels[0][165] , 
	\labels[0][164] , \labels[0][163] , \labels[0][162] , 
	\labels[0][161] , \labels[0][160] , \labels[0][159] , 
	\labels[0][158] , \labels[0][157] , \labels[0][156] , 
	\labels[0][155] , \labels[0][154] , \labels[0][153] , 
	\labels[0][152] , \labels[0][151] , \labels[0][150] , 
	\labels[0][149] , \labels[0][148] , \labels[0][147] , 
	\labels[0][146] , \labels[0][145] , \labels[0][144] , 
	\labels[0][143] , \labels[0][142] , \labels[0][141] , 
	\labels[0][140] , \labels[0][139] , \labels[0][138] , 
	\labels[0][137] , \labels[0][136] , \labels[0][135] , 
	\labels[0][134] , \labels[0][133] , \labels[0][132] , 
	\labels[0][131] , \labels[0][130] , \labels[0][129] , 
	\labels[0][128] , \labels[0][127] , \labels[0][126] , 
	\labels[0][125] , \labels[0][124] , \labels[0][123] , 
	\labels[0][122] , \labels[0][121] , \labels[0][120] , 
	\labels[0][119] , \labels[0][118] , \labels[0][117] , 
	\labels[0][116] , \labels[0][115] , \labels[0][114] , 
	\labels[0][113] , \labels[0][112] , \labels[0][111] , 
	\labels[0][110] , \labels[0][109] , \labels[0][108] , 
	\labels[0][107] , \labels[0][106] , \labels[0][105] , 
	\labels[0][104] , \labels[0][103] , \labels[0][102] , 
	\labels[0][101] , \labels[0][100] , \labels[0][99] , \labels[0][98] , 
	\labels[0][97] , \labels[0][96] , \labels[0][95] , \labels[0][94] , 
	\labels[0][93] , \labels[0][92] , \labels[0][91] , \labels[0][90] , 
	\labels[0][89] , \labels[0][88] , \labels[0][87] , \labels[0][86] , 
	\labels[0][85] , \labels[0][84] , \labels[0][83] , \labels[0][82] , 
	\labels[0][81] , \labels[0][80] , \labels[0][79] , \labels[0][78] , 
	\labels[0][77] , \labels[0][76] , \labels[0][75] , \labels[0][74] , 
	\labels[0][73] , \labels[0][72] , \labels[0][71] , \labels[0][70] , 
	\labels[0][69] , \labels[0][68] , \labels[0][67] , \labels[0][66] , 
	\labels[0][65] , \labels[0][64] , \labels[0][63] , \labels[0][62] , 
	\labels[0][61] , \labels[0][60] , \labels[0][59] , \labels[0][58] , 
	\labels[0][57] , \labels[0][56] , \labels[0][55] , \labels[0][54] , 
	\labels[0][53] , \labels[0][52] , \labels[0][51] , \labels[0][50] , 
	\labels[0][49] , \labels[0][48] , \labels[0][47] , \labels[0][46] , 
	\labels[0][45] , \labels[0][44] , \labels[0][43] , \labels[0][42] , 
	\labels[0][41] , \labels[0][40] , \labels[0][39] , \labels[0][38] , 
	\labels[0][37] , \labels[0][36] , \labels[0][35] , \labels[0][34] , 
	\labels[0][33] , \labels[0][32] , \labels[0][31] , \labels[0][30] , 
	\labels[0][29] , \labels[0][28] , \labels[0][27] , \labels[0][26] , 
	\labels[0][25] , \labels[0][24] , \labels[0][23] , \labels[0][22] , 
	\labels[0][21] , \labels[0][20] , \labels[0][19] , \labels[0][18] , 
	\labels[0][17] , \labels[0][16] , \labels[0][15] , \labels[0][14] , 
	\labels[0][13] , \labels[0][12] , \labels[0][11] , \labels[0][10] , 
	\labels[0][9] , \labels[0][8] , \labels[0][7] , \labels[0][6] , 
	\labels[0][5] , \labels[0][4] , \labels[0][3] , \labels[0][2] , 
	\labels[0][1] , \labels[0][0] });
cr_kme_regfile u_cr_kme_regfile ( .suppress_key_tlvs( suppress_key_tlvs), 
	.kme_interrupt( kme_interrupt), .rbus_ring_o( 
	_zy_simnet_rbus_ring_o_35_w$[0:83]), .kme_cceip0_ob_out( 
	_zy_simnet_kme_cceip0_ob_out_36_w$[0:82]), .kme_cceip0_ob_in_mod( 
	_zy_simnet_kme_cceip0_ob_in_mod_37_w$), .kme_cceip1_ob_out( 
	_zy_simnet_kme_cceip1_ob_out_38_w$[0:82]), .kme_cceip1_ob_in_mod( 
	_zy_simnet_kme_cceip1_ob_in_mod_39_w$), .kme_cceip2_ob_out( 
	_zy_simnet_kme_cceip2_ob_out_40_w$[0:82]), .kme_cceip2_ob_in_mod( 
	_zy_simnet_kme_cceip2_ob_in_mod_41_w$), .kme_cceip3_ob_out( 
	_zy_simnet_kme_cceip3_ob_out_42_w$[0:82]), .kme_cceip3_ob_in_mod( 
	_zy_simnet_kme_cceip3_ob_in_mod_43_w$), .kme_cddip0_ob_out( 
	_zy_simnet_kme_cddip0_ob_out_44_w$[0:82]), .kme_cddip0_ob_in_mod( 
	_zy_simnet_kme_cddip0_ob_in_mod_45_w$), .kme_cddip1_ob_out( 
	_zy_simnet_kme_cddip1_ob_out_46_w$[0:82]), .kme_cddip1_ob_in_mod( 
	_zy_simnet_kme_cddip1_ob_in_mod_47_w$), .kme_cddip2_ob_out( 
	_zy_simnet_kme_cddip2_ob_out_48_w$[0:82]), .kme_cddip2_ob_in_mod( 
	_zy_simnet_kme_cddip2_ob_in_mod_49_w$), .kme_cddip3_ob_out( 
	_zy_simnet_kme_cddip3_ob_out_50_w$[0:82]), .kme_cddip3_ob_in_mod( 
	_zy_simnet_kme_cddip3_ob_in_mod_51_w$), .ckv_dout( ckv_dout[63:0]), 
	.ckv_mbe( ckv_mbe), .kim_dout( _zy_simnet_kim_dout_52_w$[0:37]), 
	.kim_mbe( kim_mbe), .bimc_rst_n( bimc_rst_n), 
	.cceip_encrypt_bimc_isync( cceip_encrypt_bimc_isync), 
	.cceip_encrypt_bimc_idat( cceip_encrypt_bimc_idat), 
	.cceip_validate_bimc_isync( cceip_validate_bimc_isync), 
	.cceip_validate_bimc_idat( cceip_validate_bimc_idat), 
	.cddip_decrypt_bimc_isync( cddip_decrypt_bimc_isync), 
	.cddip_decrypt_bimc_idat( cddip_decrypt_bimc_idat), 
	.axi_bimc_isync( axi_bimc_isync), .axi_bimc_idat( axi_bimc_idat), 
	.labels( { \_zy_simnet_tvar_53[7][271] , 
	\_zy_simnet_tvar_53[7][270] , \_zy_simnet_tvar_53[7][269] , 
	\_zy_simnet_tvar_53[7][268] , \_zy_simnet_tvar_53[7][267] , 
	\_zy_simnet_tvar_53[7][266] , \_zy_simnet_tvar_53[7][265] , 
	\_zy_simnet_tvar_53[7][264] , \_zy_simnet_tvar_53[7][263] , 
	\_zy_simnet_tvar_53[7][262] , \_zy_simnet_tvar_53[7][261] , 
	\_zy_simnet_tvar_53[7][260] , \_zy_simnet_tvar_53[7][259] , 
	\_zy_simnet_tvar_53[7][258] , \_zy_simnet_tvar_53[7][257] , 
	\_zy_simnet_tvar_53[7][256] , \_zy_simnet_tvar_53[7][255] , 
	\_zy_simnet_tvar_53[7][254] , \_zy_simnet_tvar_53[7][253] , 
	\_zy_simnet_tvar_53[7][252] , \_zy_simnet_tvar_53[7][251] , 
	\_zy_simnet_tvar_53[7][250] , \_zy_simnet_tvar_53[7][249] , 
	\_zy_simnet_tvar_53[7][248] , \_zy_simnet_tvar_53[7][247] , 
	\_zy_simnet_tvar_53[7][246] , \_zy_simnet_tvar_53[7][245] , 
	\_zy_simnet_tvar_53[7][244] , \_zy_simnet_tvar_53[7][243] , 
	\_zy_simnet_tvar_53[7][242] , \_zy_simnet_tvar_53[7][241] , 
	\_zy_simnet_tvar_53[7][240] , \_zy_simnet_tvar_53[7][239] , 
	\_zy_simnet_tvar_53[7][238] , \_zy_simnet_tvar_53[7][237] , 
	\_zy_simnet_tvar_53[7][236] , \_zy_simnet_tvar_53[7][235] , 
	\_zy_simnet_tvar_53[7][234] , \_zy_simnet_tvar_53[7][233] , 
	\_zy_simnet_tvar_53[7][232] , \_zy_simnet_tvar_53[7][231] , 
	\_zy_simnet_tvar_53[7][230] , \_zy_simnet_tvar_53[7][229] , 
	\_zy_simnet_tvar_53[7][228] , \_zy_simnet_tvar_53[7][227] , 
	\_zy_simnet_tvar_53[7][226] , \_zy_simnet_tvar_53[7][225] , 
	\_zy_simnet_tvar_53[7][224] , \_zy_simnet_tvar_53[7][223] , 
	\_zy_simnet_tvar_53[7][222] , \_zy_simnet_tvar_53[7][221] , 
	\_zy_simnet_tvar_53[7][220] , \_zy_simnet_tvar_53[7][219] , 
	\_zy_simnet_tvar_53[7][218] , \_zy_simnet_tvar_53[7][217] , 
	\_zy_simnet_tvar_53[7][216] , \_zy_simnet_tvar_53[7][215] , 
	\_zy_simnet_tvar_53[7][214] , \_zy_simnet_tvar_53[7][213] , 
	\_zy_simnet_tvar_53[7][212] , \_zy_simnet_tvar_53[7][211] , 
	\_zy_simnet_tvar_53[7][210] , \_zy_simnet_tvar_53[7][209] , 
	\_zy_simnet_tvar_53[7][208] , \_zy_simnet_tvar_53[7][207] , 
	\_zy_simnet_tvar_53[7][206] , \_zy_simnet_tvar_53[7][205] , 
	\_zy_simnet_tvar_53[7][204] , \_zy_simnet_tvar_53[7][203] , 
	\_zy_simnet_tvar_53[7][202] , \_zy_simnet_tvar_53[7][201] , 
	\_zy_simnet_tvar_53[7][200] , \_zy_simnet_tvar_53[7][199] , 
	\_zy_simnet_tvar_53[7][198] , \_zy_simnet_tvar_53[7][197] , 
	\_zy_simnet_tvar_53[7][196] , \_zy_simnet_tvar_53[7][195] , 
	\_zy_simnet_tvar_53[7][194] , \_zy_simnet_tvar_53[7][193] , 
	\_zy_simnet_tvar_53[7][192] , \_zy_simnet_tvar_53[7][191] , 
	\_zy_simnet_tvar_53[7][190] , \_zy_simnet_tvar_53[7][189] , 
	\_zy_simnet_tvar_53[7][188] , \_zy_simnet_tvar_53[7][187] , 
	\_zy_simnet_tvar_53[7][186] , \_zy_simnet_tvar_53[7][185] , 
	\_zy_simnet_tvar_53[7][184] , \_zy_simnet_tvar_53[7][183] , 
	\_zy_simnet_tvar_53[7][182] , \_zy_simnet_tvar_53[7][181] , 
	\_zy_simnet_tvar_53[7][180] , \_zy_simnet_tvar_53[7][179] , 
	\_zy_simnet_tvar_53[7][178] , \_zy_simnet_tvar_53[7][177] , 
	\_zy_simnet_tvar_53[7][176] , \_zy_simnet_tvar_53[7][175] , 
	\_zy_simnet_tvar_53[7][174] , \_zy_simnet_tvar_53[7][173] , 
	\_zy_simnet_tvar_53[7][172] , \_zy_simnet_tvar_53[7][171] , 
	\_zy_simnet_tvar_53[7][170] , \_zy_simnet_tvar_53[7][169] , 
	\_zy_simnet_tvar_53[7][168] , \_zy_simnet_tvar_53[7][167] , 
	\_zy_simnet_tvar_53[7][166] , \_zy_simnet_tvar_53[7][165] , 
	\_zy_simnet_tvar_53[7][164] , \_zy_simnet_tvar_53[7][163] , 
	\_zy_simnet_tvar_53[7][162] , \_zy_simnet_tvar_53[7][161] , 
	\_zy_simnet_tvar_53[7][160] , \_zy_simnet_tvar_53[7][159] , 
	\_zy_simnet_tvar_53[7][158] , \_zy_simnet_tvar_53[7][157] , 
	\_zy_simnet_tvar_53[7][156] , \_zy_simnet_tvar_53[7][155] , 
	\_zy_simnet_tvar_53[7][154] , \_zy_simnet_tvar_53[7][153] , 
	\_zy_simnet_tvar_53[7][152] , \_zy_simnet_tvar_53[7][151] , 
	\_zy_simnet_tvar_53[7][150] , \_zy_simnet_tvar_53[7][149] , 
	\_zy_simnet_tvar_53[7][148] , \_zy_simnet_tvar_53[7][147] , 
	\_zy_simnet_tvar_53[7][146] , \_zy_simnet_tvar_53[7][145] , 
	\_zy_simnet_tvar_53[7][144] , \_zy_simnet_tvar_53[7][143] , 
	\_zy_simnet_tvar_53[7][142] , \_zy_simnet_tvar_53[7][141] , 
	\_zy_simnet_tvar_53[7][140] , \_zy_simnet_tvar_53[7][139] , 
	\_zy_simnet_tvar_53[7][138] , \_zy_simnet_tvar_53[7][137] , 
	\_zy_simnet_tvar_53[7][136] , \_zy_simnet_tvar_53[7][135] , 
	\_zy_simnet_tvar_53[7][134] , \_zy_simnet_tvar_53[7][133] , 
	\_zy_simnet_tvar_53[7][132] , \_zy_simnet_tvar_53[7][131] , 
	\_zy_simnet_tvar_53[7][130] , \_zy_simnet_tvar_53[7][129] , 
	\_zy_simnet_tvar_53[7][128] , \_zy_simnet_tvar_53[7][127] , 
	\_zy_simnet_tvar_53[7][126] , \_zy_simnet_tvar_53[7][125] , 
	\_zy_simnet_tvar_53[7][124] , \_zy_simnet_tvar_53[7][123] , 
	\_zy_simnet_tvar_53[7][122] , \_zy_simnet_tvar_53[7][121] , 
	\_zy_simnet_tvar_53[7][120] , \_zy_simnet_tvar_53[7][119] , 
	\_zy_simnet_tvar_53[7][118] , \_zy_simnet_tvar_53[7][117] , 
	\_zy_simnet_tvar_53[7][116] , \_zy_simnet_tvar_53[7][115] , 
	\_zy_simnet_tvar_53[7][114] , \_zy_simnet_tvar_53[7][113] , 
	\_zy_simnet_tvar_53[7][112] , \_zy_simnet_tvar_53[7][111] , 
	\_zy_simnet_tvar_53[7][110] , \_zy_simnet_tvar_53[7][109] , 
	\_zy_simnet_tvar_53[7][108] , \_zy_simnet_tvar_53[7][107] , 
	\_zy_simnet_tvar_53[7][106] , \_zy_simnet_tvar_53[7][105] , 
	\_zy_simnet_tvar_53[7][104] , \_zy_simnet_tvar_53[7][103] , 
	\_zy_simnet_tvar_53[7][102] , \_zy_simnet_tvar_53[7][101] , 
	\_zy_simnet_tvar_53[7][100] , \_zy_simnet_tvar_53[7][99] , 
	\_zy_simnet_tvar_53[7][98] , \_zy_simnet_tvar_53[7][97] , 
	\_zy_simnet_tvar_53[7][96] , \_zy_simnet_tvar_53[7][95] , 
	\_zy_simnet_tvar_53[7][94] , \_zy_simnet_tvar_53[7][93] , 
	\_zy_simnet_tvar_53[7][92] , \_zy_simnet_tvar_53[7][91] , 
	\_zy_simnet_tvar_53[7][90] , \_zy_simnet_tvar_53[7][89] , 
	\_zy_simnet_tvar_53[7][88] , \_zy_simnet_tvar_53[7][87] , 
	\_zy_simnet_tvar_53[7][86] , \_zy_simnet_tvar_53[7][85] , 
	\_zy_simnet_tvar_53[7][84] , \_zy_simnet_tvar_53[7][83] , 
	\_zy_simnet_tvar_53[7][82] , \_zy_simnet_tvar_53[7][81] , 
	\_zy_simnet_tvar_53[7][80] , \_zy_simnet_tvar_53[7][79] , 
	\_zy_simnet_tvar_53[7][78] , \_zy_simnet_tvar_53[7][77] , 
	\_zy_simnet_tvar_53[7][76] , \_zy_simnet_tvar_53[7][75] , 
	\_zy_simnet_tvar_53[7][74] , \_zy_simnet_tvar_53[7][73] , 
	\_zy_simnet_tvar_53[7][72] , \_zy_simnet_tvar_53[7][71] , 
	\_zy_simnet_tvar_53[7][70] , \_zy_simnet_tvar_53[7][69] , 
	\_zy_simnet_tvar_53[7][68] , \_zy_simnet_tvar_53[7][67] , 
	\_zy_simnet_tvar_53[7][66] , \_zy_simnet_tvar_53[7][65] , 
	\_zy_simnet_tvar_53[7][64] , \_zy_simnet_tvar_53[7][63] , 
	\_zy_simnet_tvar_53[7][62] , \_zy_simnet_tvar_53[7][61] , 
	\_zy_simnet_tvar_53[7][60] , \_zy_simnet_tvar_53[7][59] , 
	\_zy_simnet_tvar_53[7][58] , \_zy_simnet_tvar_53[7][57] , 
	\_zy_simnet_tvar_53[7][56] , \_zy_simnet_tvar_53[7][55] , 
	\_zy_simnet_tvar_53[7][54] , \_zy_simnet_tvar_53[7][53] , 
	\_zy_simnet_tvar_53[7][52] , \_zy_simnet_tvar_53[7][51] , 
	\_zy_simnet_tvar_53[7][50] , \_zy_simnet_tvar_53[7][49] , 
	\_zy_simnet_tvar_53[7][48] , \_zy_simnet_tvar_53[7][47] , 
	\_zy_simnet_tvar_53[7][46] , \_zy_simnet_tvar_53[7][45] , 
	\_zy_simnet_tvar_53[7][44] , \_zy_simnet_tvar_53[7][43] , 
	\_zy_simnet_tvar_53[7][42] , \_zy_simnet_tvar_53[7][41] , 
	\_zy_simnet_tvar_53[7][40] , \_zy_simnet_tvar_53[7][39] , 
	\_zy_simnet_tvar_53[7][38] , \_zy_simnet_tvar_53[7][37] , 
	\_zy_simnet_tvar_53[7][36] , \_zy_simnet_tvar_53[7][35] , 
	\_zy_simnet_tvar_53[7][34] , \_zy_simnet_tvar_53[7][33] , 
	\_zy_simnet_tvar_53[7][32] , \_zy_simnet_tvar_53[7][31] , 
	\_zy_simnet_tvar_53[7][30] , \_zy_simnet_tvar_53[7][29] , 
	\_zy_simnet_tvar_53[7][28] , \_zy_simnet_tvar_53[7][27] , 
	\_zy_simnet_tvar_53[7][26] , \_zy_simnet_tvar_53[7][25] , 
	\_zy_simnet_tvar_53[7][24] , \_zy_simnet_tvar_53[7][23] , 
	\_zy_simnet_tvar_53[7][22] , \_zy_simnet_tvar_53[7][21] , 
	\_zy_simnet_tvar_53[7][20] , \_zy_simnet_tvar_53[7][19] , 
	\_zy_simnet_tvar_53[7][18] , \_zy_simnet_tvar_53[7][17] , 
	\_zy_simnet_tvar_53[7][16] , \_zy_simnet_tvar_53[7][15] , 
	\_zy_simnet_tvar_53[7][14] , \_zy_simnet_tvar_53[7][13] , 
	\_zy_simnet_tvar_53[7][12] , \_zy_simnet_tvar_53[7][11] , 
	\_zy_simnet_tvar_53[7][10] , \_zy_simnet_tvar_53[7][9] , 
	\_zy_simnet_tvar_53[7][8] , \_zy_simnet_tvar_53[7][7] , 
	\_zy_simnet_tvar_53[7][6] , \_zy_simnet_tvar_53[7][5] , 
	\_zy_simnet_tvar_53[7][4] , \_zy_simnet_tvar_53[7][3] , 
	\_zy_simnet_tvar_53[7][2] , \_zy_simnet_tvar_53[7][1] , 
	\_zy_simnet_tvar_53[7][0] , \_zy_simnet_tvar_53[6][271] , 
	\_zy_simnet_tvar_53[6][270] , \_zy_simnet_tvar_53[6][269] , 
	\_zy_simnet_tvar_53[6][268] , \_zy_simnet_tvar_53[6][267] , 
	\_zy_simnet_tvar_53[6][266] , \_zy_simnet_tvar_53[6][265] , 
	\_zy_simnet_tvar_53[6][264] , \_zy_simnet_tvar_53[6][263] , 
	\_zy_simnet_tvar_53[6][262] , \_zy_simnet_tvar_53[6][261] , 
	\_zy_simnet_tvar_53[6][260] , \_zy_simnet_tvar_53[6][259] , 
	\_zy_simnet_tvar_53[6][258] , \_zy_simnet_tvar_53[6][257] , 
	\_zy_simnet_tvar_53[6][256] , \_zy_simnet_tvar_53[6][255] , 
	\_zy_simnet_tvar_53[6][254] , \_zy_simnet_tvar_53[6][253] , 
	\_zy_simnet_tvar_53[6][252] , \_zy_simnet_tvar_53[6][251] , 
	\_zy_simnet_tvar_53[6][250] , \_zy_simnet_tvar_53[6][249] , 
	\_zy_simnet_tvar_53[6][248] , \_zy_simnet_tvar_53[6][247] , 
	\_zy_simnet_tvar_53[6][246] , \_zy_simnet_tvar_53[6][245] , 
	\_zy_simnet_tvar_53[6][244] , \_zy_simnet_tvar_53[6][243] , 
	\_zy_simnet_tvar_53[6][242] , \_zy_simnet_tvar_53[6][241] , 
	\_zy_simnet_tvar_53[6][240] , \_zy_simnet_tvar_53[6][239] , 
	\_zy_simnet_tvar_53[6][238] , \_zy_simnet_tvar_53[6][237] , 
	\_zy_simnet_tvar_53[6][236] , \_zy_simnet_tvar_53[6][235] , 
	\_zy_simnet_tvar_53[6][234] , \_zy_simnet_tvar_53[6][233] , 
	\_zy_simnet_tvar_53[6][232] , \_zy_simnet_tvar_53[6][231] , 
	\_zy_simnet_tvar_53[6][230] , \_zy_simnet_tvar_53[6][229] , 
	\_zy_simnet_tvar_53[6][228] , \_zy_simnet_tvar_53[6][227] , 
	\_zy_simnet_tvar_53[6][226] , \_zy_simnet_tvar_53[6][225] , 
	\_zy_simnet_tvar_53[6][224] , \_zy_simnet_tvar_53[6][223] , 
	\_zy_simnet_tvar_53[6][222] , \_zy_simnet_tvar_53[6][221] , 
	\_zy_simnet_tvar_53[6][220] , \_zy_simnet_tvar_53[6][219] , 
	\_zy_simnet_tvar_53[6][218] , \_zy_simnet_tvar_53[6][217] , 
	\_zy_simnet_tvar_53[6][216] , \_zy_simnet_tvar_53[6][215] , 
	\_zy_simnet_tvar_53[6][214] , \_zy_simnet_tvar_53[6][213] , 
	\_zy_simnet_tvar_53[6][212] , \_zy_simnet_tvar_53[6][211] , 
	\_zy_simnet_tvar_53[6][210] , \_zy_simnet_tvar_53[6][209] , 
	\_zy_simnet_tvar_53[6][208] , \_zy_simnet_tvar_53[6][207] , 
	\_zy_simnet_tvar_53[6][206] , \_zy_simnet_tvar_53[6][205] , 
	\_zy_simnet_tvar_53[6][204] , \_zy_simnet_tvar_53[6][203] , 
	\_zy_simnet_tvar_53[6][202] , \_zy_simnet_tvar_53[6][201] , 
	\_zy_simnet_tvar_53[6][200] , \_zy_simnet_tvar_53[6][199] , 
	\_zy_simnet_tvar_53[6][198] , \_zy_simnet_tvar_53[6][197] , 
	\_zy_simnet_tvar_53[6][196] , \_zy_simnet_tvar_53[6][195] , 
	\_zy_simnet_tvar_53[6][194] , \_zy_simnet_tvar_53[6][193] , 
	\_zy_simnet_tvar_53[6][192] , \_zy_simnet_tvar_53[6][191] , 
	\_zy_simnet_tvar_53[6][190] , \_zy_simnet_tvar_53[6][189] , 
	\_zy_simnet_tvar_53[6][188] , \_zy_simnet_tvar_53[6][187] , 
	\_zy_simnet_tvar_53[6][186] , \_zy_simnet_tvar_53[6][185] , 
	\_zy_simnet_tvar_53[6][184] , \_zy_simnet_tvar_53[6][183] , 
	\_zy_simnet_tvar_53[6][182] , \_zy_simnet_tvar_53[6][181] , 
	\_zy_simnet_tvar_53[6][180] , \_zy_simnet_tvar_53[6][179] , 
	\_zy_simnet_tvar_53[6][178] , \_zy_simnet_tvar_53[6][177] , 
	\_zy_simnet_tvar_53[6][176] , \_zy_simnet_tvar_53[6][175] , 
	\_zy_simnet_tvar_53[6][174] , \_zy_simnet_tvar_53[6][173] , 
	\_zy_simnet_tvar_53[6][172] , \_zy_simnet_tvar_53[6][171] , 
	\_zy_simnet_tvar_53[6][170] , \_zy_simnet_tvar_53[6][169] , 
	\_zy_simnet_tvar_53[6][168] , \_zy_simnet_tvar_53[6][167] , 
	\_zy_simnet_tvar_53[6][166] , \_zy_simnet_tvar_53[6][165] , 
	\_zy_simnet_tvar_53[6][164] , \_zy_simnet_tvar_53[6][163] , 
	\_zy_simnet_tvar_53[6][162] , \_zy_simnet_tvar_53[6][161] , 
	\_zy_simnet_tvar_53[6][160] , \_zy_simnet_tvar_53[6][159] , 
	\_zy_simnet_tvar_53[6][158] , \_zy_simnet_tvar_53[6][157] , 
	\_zy_simnet_tvar_53[6][156] , \_zy_simnet_tvar_53[6][155] , 
	\_zy_simnet_tvar_53[6][154] , \_zy_simnet_tvar_53[6][153] , 
	\_zy_simnet_tvar_53[6][152] , \_zy_simnet_tvar_53[6][151] , 
	\_zy_simnet_tvar_53[6][150] , \_zy_simnet_tvar_53[6][149] , 
	\_zy_simnet_tvar_53[6][148] , \_zy_simnet_tvar_53[6][147] , 
	\_zy_simnet_tvar_53[6][146] , \_zy_simnet_tvar_53[6][145] , 
	\_zy_simnet_tvar_53[6][144] , \_zy_simnet_tvar_53[6][143] , 
	\_zy_simnet_tvar_53[6][142] , \_zy_simnet_tvar_53[6][141] , 
	\_zy_simnet_tvar_53[6][140] , \_zy_simnet_tvar_53[6][139] , 
	\_zy_simnet_tvar_53[6][138] , \_zy_simnet_tvar_53[6][137] , 
	\_zy_simnet_tvar_53[6][136] , \_zy_simnet_tvar_53[6][135] , 
	\_zy_simnet_tvar_53[6][134] , \_zy_simnet_tvar_53[6][133] , 
	\_zy_simnet_tvar_53[6][132] , \_zy_simnet_tvar_53[6][131] , 
	\_zy_simnet_tvar_53[6][130] , \_zy_simnet_tvar_53[6][129] , 
	\_zy_simnet_tvar_53[6][128] , \_zy_simnet_tvar_53[6][127] , 
	\_zy_simnet_tvar_53[6][126] , \_zy_simnet_tvar_53[6][125] , 
	\_zy_simnet_tvar_53[6][124] , \_zy_simnet_tvar_53[6][123] , 
	\_zy_simnet_tvar_53[6][122] , \_zy_simnet_tvar_53[6][121] , 
	\_zy_simnet_tvar_53[6][120] , \_zy_simnet_tvar_53[6][119] , 
	\_zy_simnet_tvar_53[6][118] , \_zy_simnet_tvar_53[6][117] , 
	\_zy_simnet_tvar_53[6][116] , \_zy_simnet_tvar_53[6][115] , 
	\_zy_simnet_tvar_53[6][114] , \_zy_simnet_tvar_53[6][113] , 
	\_zy_simnet_tvar_53[6][112] , \_zy_simnet_tvar_53[6][111] , 
	\_zy_simnet_tvar_53[6][110] , \_zy_simnet_tvar_53[6][109] , 
	\_zy_simnet_tvar_53[6][108] , \_zy_simnet_tvar_53[6][107] , 
	\_zy_simnet_tvar_53[6][106] , \_zy_simnet_tvar_53[6][105] , 
	\_zy_simnet_tvar_53[6][104] , \_zy_simnet_tvar_53[6][103] , 
	\_zy_simnet_tvar_53[6][102] , \_zy_simnet_tvar_53[6][101] , 
	\_zy_simnet_tvar_53[6][100] , \_zy_simnet_tvar_53[6][99] , 
	\_zy_simnet_tvar_53[6][98] , \_zy_simnet_tvar_53[6][97] , 
	\_zy_simnet_tvar_53[6][96] , \_zy_simnet_tvar_53[6][95] , 
	\_zy_simnet_tvar_53[6][94] , \_zy_simnet_tvar_53[6][93] , 
	\_zy_simnet_tvar_53[6][92] , \_zy_simnet_tvar_53[6][91] , 
	\_zy_simnet_tvar_53[6][90] , \_zy_simnet_tvar_53[6][89] , 
	\_zy_simnet_tvar_53[6][88] , \_zy_simnet_tvar_53[6][87] , 
	\_zy_simnet_tvar_53[6][86] , \_zy_simnet_tvar_53[6][85] , 
	\_zy_simnet_tvar_53[6][84] , \_zy_simnet_tvar_53[6][83] , 
	\_zy_simnet_tvar_53[6][82] , \_zy_simnet_tvar_53[6][81] , 
	\_zy_simnet_tvar_53[6][80] , \_zy_simnet_tvar_53[6][79] , 
	\_zy_simnet_tvar_53[6][78] , \_zy_simnet_tvar_53[6][77] , 
	\_zy_simnet_tvar_53[6][76] , \_zy_simnet_tvar_53[6][75] , 
	\_zy_simnet_tvar_53[6][74] , \_zy_simnet_tvar_53[6][73] , 
	\_zy_simnet_tvar_53[6][72] , \_zy_simnet_tvar_53[6][71] , 
	\_zy_simnet_tvar_53[6][70] , \_zy_simnet_tvar_53[6][69] , 
	\_zy_simnet_tvar_53[6][68] , \_zy_simnet_tvar_53[6][67] , 
	\_zy_simnet_tvar_53[6][66] , \_zy_simnet_tvar_53[6][65] , 
	\_zy_simnet_tvar_53[6][64] , \_zy_simnet_tvar_53[6][63] , 
	\_zy_simnet_tvar_53[6][62] , \_zy_simnet_tvar_53[6][61] , 
	\_zy_simnet_tvar_53[6][60] , \_zy_simnet_tvar_53[6][59] , 
	\_zy_simnet_tvar_53[6][58] , \_zy_simnet_tvar_53[6][57] , 
	\_zy_simnet_tvar_53[6][56] , \_zy_simnet_tvar_53[6][55] , 
	\_zy_simnet_tvar_53[6][54] , \_zy_simnet_tvar_53[6][53] , 
	\_zy_simnet_tvar_53[6][52] , \_zy_simnet_tvar_53[6][51] , 
	\_zy_simnet_tvar_53[6][50] , \_zy_simnet_tvar_53[6][49] , 
	\_zy_simnet_tvar_53[6][48] , \_zy_simnet_tvar_53[6][47] , 
	\_zy_simnet_tvar_53[6][46] , \_zy_simnet_tvar_53[6][45] , 
	\_zy_simnet_tvar_53[6][44] , \_zy_simnet_tvar_53[6][43] , 
	\_zy_simnet_tvar_53[6][42] , \_zy_simnet_tvar_53[6][41] , 
	\_zy_simnet_tvar_53[6][40] , \_zy_simnet_tvar_53[6][39] , 
	\_zy_simnet_tvar_53[6][38] , \_zy_simnet_tvar_53[6][37] , 
	\_zy_simnet_tvar_53[6][36] , \_zy_simnet_tvar_53[6][35] , 
	\_zy_simnet_tvar_53[6][34] , \_zy_simnet_tvar_53[6][33] , 
	\_zy_simnet_tvar_53[6][32] , \_zy_simnet_tvar_53[6][31] , 
	\_zy_simnet_tvar_53[6][30] , \_zy_simnet_tvar_53[6][29] , 
	\_zy_simnet_tvar_53[6][28] , \_zy_simnet_tvar_53[6][27] , 
	\_zy_simnet_tvar_53[6][26] , \_zy_simnet_tvar_53[6][25] , 
	\_zy_simnet_tvar_53[6][24] , \_zy_simnet_tvar_53[6][23] , 
	\_zy_simnet_tvar_53[6][22] , \_zy_simnet_tvar_53[6][21] , 
	\_zy_simnet_tvar_53[6][20] , \_zy_simnet_tvar_53[6][19] , 
	\_zy_simnet_tvar_53[6][18] , \_zy_simnet_tvar_53[6][17] , 
	\_zy_simnet_tvar_53[6][16] , \_zy_simnet_tvar_53[6][15] , 
	\_zy_simnet_tvar_53[6][14] , \_zy_simnet_tvar_53[6][13] , 
	\_zy_simnet_tvar_53[6][12] , \_zy_simnet_tvar_53[6][11] , 
	\_zy_simnet_tvar_53[6][10] , \_zy_simnet_tvar_53[6][9] , 
	\_zy_simnet_tvar_53[6][8] , \_zy_simnet_tvar_53[6][7] , 
	\_zy_simnet_tvar_53[6][6] , \_zy_simnet_tvar_53[6][5] , 
	\_zy_simnet_tvar_53[6][4] , \_zy_simnet_tvar_53[6][3] , 
	\_zy_simnet_tvar_53[6][2] , \_zy_simnet_tvar_53[6][1] , 
	\_zy_simnet_tvar_53[6][0] , \_zy_simnet_tvar_53[5][271] , 
	\_zy_simnet_tvar_53[5][270] , \_zy_simnet_tvar_53[5][269] , 
	\_zy_simnet_tvar_53[5][268] , \_zy_simnet_tvar_53[5][267] , 
	\_zy_simnet_tvar_53[5][266] , \_zy_simnet_tvar_53[5][265] , 
	\_zy_simnet_tvar_53[5][264] , \_zy_simnet_tvar_53[5][263] , 
	\_zy_simnet_tvar_53[5][262] , \_zy_simnet_tvar_53[5][261] , 
	\_zy_simnet_tvar_53[5][260] , \_zy_simnet_tvar_53[5][259] , 
	\_zy_simnet_tvar_53[5][258] , \_zy_simnet_tvar_53[5][257] , 
	\_zy_simnet_tvar_53[5][256] , \_zy_simnet_tvar_53[5][255] , 
	\_zy_simnet_tvar_53[5][254] , \_zy_simnet_tvar_53[5][253] , 
	\_zy_simnet_tvar_53[5][252] , \_zy_simnet_tvar_53[5][251] , 
	\_zy_simnet_tvar_53[5][250] , \_zy_simnet_tvar_53[5][249] , 
	\_zy_simnet_tvar_53[5][248] , \_zy_simnet_tvar_53[5][247] , 
	\_zy_simnet_tvar_53[5][246] , \_zy_simnet_tvar_53[5][245] , 
	\_zy_simnet_tvar_53[5][244] , \_zy_simnet_tvar_53[5][243] , 
	\_zy_simnet_tvar_53[5][242] , \_zy_simnet_tvar_53[5][241] , 
	\_zy_simnet_tvar_53[5][240] , \_zy_simnet_tvar_53[5][239] , 
	\_zy_simnet_tvar_53[5][238] , \_zy_simnet_tvar_53[5][237] , 
	\_zy_simnet_tvar_53[5][236] , \_zy_simnet_tvar_53[5][235] , 
	\_zy_simnet_tvar_53[5][234] , \_zy_simnet_tvar_53[5][233] , 
	\_zy_simnet_tvar_53[5][232] , \_zy_simnet_tvar_53[5][231] , 
	\_zy_simnet_tvar_53[5][230] , \_zy_simnet_tvar_53[5][229] , 
	\_zy_simnet_tvar_53[5][228] , \_zy_simnet_tvar_53[5][227] , 
	\_zy_simnet_tvar_53[5][226] , \_zy_simnet_tvar_53[5][225] , 
	\_zy_simnet_tvar_53[5][224] , \_zy_simnet_tvar_53[5][223] , 
	\_zy_simnet_tvar_53[5][222] , \_zy_simnet_tvar_53[5][221] , 
	\_zy_simnet_tvar_53[5][220] , \_zy_simnet_tvar_53[5][219] , 
	\_zy_simnet_tvar_53[5][218] , \_zy_simnet_tvar_53[5][217] , 
	\_zy_simnet_tvar_53[5][216] , \_zy_simnet_tvar_53[5][215] , 
	\_zy_simnet_tvar_53[5][214] , \_zy_simnet_tvar_53[5][213] , 
	\_zy_simnet_tvar_53[5][212] , \_zy_simnet_tvar_53[5][211] , 
	\_zy_simnet_tvar_53[5][210] , \_zy_simnet_tvar_53[5][209] , 
	\_zy_simnet_tvar_53[5][208] , \_zy_simnet_tvar_53[5][207] , 
	\_zy_simnet_tvar_53[5][206] , \_zy_simnet_tvar_53[5][205] , 
	\_zy_simnet_tvar_53[5][204] , \_zy_simnet_tvar_53[5][203] , 
	\_zy_simnet_tvar_53[5][202] , \_zy_simnet_tvar_53[5][201] , 
	\_zy_simnet_tvar_53[5][200] , \_zy_simnet_tvar_53[5][199] , 
	\_zy_simnet_tvar_53[5][198] , \_zy_simnet_tvar_53[5][197] , 
	\_zy_simnet_tvar_53[5][196] , \_zy_simnet_tvar_53[5][195] , 
	\_zy_simnet_tvar_53[5][194] , \_zy_simnet_tvar_53[5][193] , 
	\_zy_simnet_tvar_53[5][192] , \_zy_simnet_tvar_53[5][191] , 
	\_zy_simnet_tvar_53[5][190] , \_zy_simnet_tvar_53[5][189] , 
	\_zy_simnet_tvar_53[5][188] , \_zy_simnet_tvar_53[5][187] , 
	\_zy_simnet_tvar_53[5][186] , \_zy_simnet_tvar_53[5][185] , 
	\_zy_simnet_tvar_53[5][184] , \_zy_simnet_tvar_53[5][183] , 
	\_zy_simnet_tvar_53[5][182] , \_zy_simnet_tvar_53[5][181] , 
	\_zy_simnet_tvar_53[5][180] , \_zy_simnet_tvar_53[5][179] , 
	\_zy_simnet_tvar_53[5][178] , \_zy_simnet_tvar_53[5][177] , 
	\_zy_simnet_tvar_53[5][176] , \_zy_simnet_tvar_53[5][175] , 
	\_zy_simnet_tvar_53[5][174] , \_zy_simnet_tvar_53[5][173] , 
	\_zy_simnet_tvar_53[5][172] , \_zy_simnet_tvar_53[5][171] , 
	\_zy_simnet_tvar_53[5][170] , \_zy_simnet_tvar_53[5][169] , 
	\_zy_simnet_tvar_53[5][168] , \_zy_simnet_tvar_53[5][167] , 
	\_zy_simnet_tvar_53[5][166] , \_zy_simnet_tvar_53[5][165] , 
	\_zy_simnet_tvar_53[5][164] , \_zy_simnet_tvar_53[5][163] , 
	\_zy_simnet_tvar_53[5][162] , \_zy_simnet_tvar_53[5][161] , 
	\_zy_simnet_tvar_53[5][160] , \_zy_simnet_tvar_53[5][159] , 
	\_zy_simnet_tvar_53[5][158] , \_zy_simnet_tvar_53[5][157] , 
	\_zy_simnet_tvar_53[5][156] , \_zy_simnet_tvar_53[5][155] , 
	\_zy_simnet_tvar_53[5][154] , \_zy_simnet_tvar_53[5][153] , 
	\_zy_simnet_tvar_53[5][152] , \_zy_simnet_tvar_53[5][151] , 
	\_zy_simnet_tvar_53[5][150] , \_zy_simnet_tvar_53[5][149] , 
	\_zy_simnet_tvar_53[5][148] , \_zy_simnet_tvar_53[5][147] , 
	\_zy_simnet_tvar_53[5][146] , \_zy_simnet_tvar_53[5][145] , 
	\_zy_simnet_tvar_53[5][144] , \_zy_simnet_tvar_53[5][143] , 
	\_zy_simnet_tvar_53[5][142] , \_zy_simnet_tvar_53[5][141] , 
	\_zy_simnet_tvar_53[5][140] , \_zy_simnet_tvar_53[5][139] , 
	\_zy_simnet_tvar_53[5][138] , \_zy_simnet_tvar_53[5][137] , 
	\_zy_simnet_tvar_53[5][136] , \_zy_simnet_tvar_53[5][135] , 
	\_zy_simnet_tvar_53[5][134] , \_zy_simnet_tvar_53[5][133] , 
	\_zy_simnet_tvar_53[5][132] , \_zy_simnet_tvar_53[5][131] , 
	\_zy_simnet_tvar_53[5][130] , \_zy_simnet_tvar_53[5][129] , 
	\_zy_simnet_tvar_53[5][128] , \_zy_simnet_tvar_53[5][127] , 
	\_zy_simnet_tvar_53[5][126] , \_zy_simnet_tvar_53[5][125] , 
	\_zy_simnet_tvar_53[5][124] , \_zy_simnet_tvar_53[5][123] , 
	\_zy_simnet_tvar_53[5][122] , \_zy_simnet_tvar_53[5][121] , 
	\_zy_simnet_tvar_53[5][120] , \_zy_simnet_tvar_53[5][119] , 
	\_zy_simnet_tvar_53[5][118] , \_zy_simnet_tvar_53[5][117] , 
	\_zy_simnet_tvar_53[5][116] , \_zy_simnet_tvar_53[5][115] , 
	\_zy_simnet_tvar_53[5][114] , \_zy_simnet_tvar_53[5][113] , 
	\_zy_simnet_tvar_53[5][112] , \_zy_simnet_tvar_53[5][111] , 
	\_zy_simnet_tvar_53[5][110] , \_zy_simnet_tvar_53[5][109] , 
	\_zy_simnet_tvar_53[5][108] , \_zy_simnet_tvar_53[5][107] , 
	\_zy_simnet_tvar_53[5][106] , \_zy_simnet_tvar_53[5][105] , 
	\_zy_simnet_tvar_53[5][104] , \_zy_simnet_tvar_53[5][103] , 
	\_zy_simnet_tvar_53[5][102] , \_zy_simnet_tvar_53[5][101] , 
	\_zy_simnet_tvar_53[5][100] , \_zy_simnet_tvar_53[5][99] , 
	\_zy_simnet_tvar_53[5][98] , \_zy_simnet_tvar_53[5][97] , 
	\_zy_simnet_tvar_53[5][96] , \_zy_simnet_tvar_53[5][95] , 
	\_zy_simnet_tvar_53[5][94] , \_zy_simnet_tvar_53[5][93] , 
	\_zy_simnet_tvar_53[5][92] , \_zy_simnet_tvar_53[5][91] , 
	\_zy_simnet_tvar_53[5][90] , \_zy_simnet_tvar_53[5][89] , 
	\_zy_simnet_tvar_53[5][88] , \_zy_simnet_tvar_53[5][87] , 
	\_zy_simnet_tvar_53[5][86] , \_zy_simnet_tvar_53[5][85] , 
	\_zy_simnet_tvar_53[5][84] , \_zy_simnet_tvar_53[5][83] , 
	\_zy_simnet_tvar_53[5][82] , \_zy_simnet_tvar_53[5][81] , 
	\_zy_simnet_tvar_53[5][80] , \_zy_simnet_tvar_53[5][79] , 
	\_zy_simnet_tvar_53[5][78] , \_zy_simnet_tvar_53[5][77] , 
	\_zy_simnet_tvar_53[5][76] , \_zy_simnet_tvar_53[5][75] , 
	\_zy_simnet_tvar_53[5][74] , \_zy_simnet_tvar_53[5][73] , 
	\_zy_simnet_tvar_53[5][72] , \_zy_simnet_tvar_53[5][71] , 
	\_zy_simnet_tvar_53[5][70] , \_zy_simnet_tvar_53[5][69] , 
	\_zy_simnet_tvar_53[5][68] , \_zy_simnet_tvar_53[5][67] , 
	\_zy_simnet_tvar_53[5][66] , \_zy_simnet_tvar_53[5][65] , 
	\_zy_simnet_tvar_53[5][64] , \_zy_simnet_tvar_53[5][63] , 
	\_zy_simnet_tvar_53[5][62] , \_zy_simnet_tvar_53[5][61] , 
	\_zy_simnet_tvar_53[5][60] , \_zy_simnet_tvar_53[5][59] , 
	\_zy_simnet_tvar_53[5][58] , \_zy_simnet_tvar_53[5][57] , 
	\_zy_simnet_tvar_53[5][56] , \_zy_simnet_tvar_53[5][55] , 
	\_zy_simnet_tvar_53[5][54] , \_zy_simnet_tvar_53[5][53] , 
	\_zy_simnet_tvar_53[5][52] , \_zy_simnet_tvar_53[5][51] , 
	\_zy_simnet_tvar_53[5][50] , \_zy_simnet_tvar_53[5][49] , 
	\_zy_simnet_tvar_53[5][48] , \_zy_simnet_tvar_53[5][47] , 
	\_zy_simnet_tvar_53[5][46] , \_zy_simnet_tvar_53[5][45] , 
	\_zy_simnet_tvar_53[5][44] , \_zy_simnet_tvar_53[5][43] , 
	\_zy_simnet_tvar_53[5][42] , \_zy_simnet_tvar_53[5][41] , 
	\_zy_simnet_tvar_53[5][40] , \_zy_simnet_tvar_53[5][39] , 
	\_zy_simnet_tvar_53[5][38] , \_zy_simnet_tvar_53[5][37] , 
	\_zy_simnet_tvar_53[5][36] , \_zy_simnet_tvar_53[5][35] , 
	\_zy_simnet_tvar_53[5][34] , \_zy_simnet_tvar_53[5][33] , 
	\_zy_simnet_tvar_53[5][32] , \_zy_simnet_tvar_53[5][31] , 
	\_zy_simnet_tvar_53[5][30] , \_zy_simnet_tvar_53[5][29] , 
	\_zy_simnet_tvar_53[5][28] , \_zy_simnet_tvar_53[5][27] , 
	\_zy_simnet_tvar_53[5][26] , \_zy_simnet_tvar_53[5][25] , 
	\_zy_simnet_tvar_53[5][24] , \_zy_simnet_tvar_53[5][23] , 
	\_zy_simnet_tvar_53[5][22] , \_zy_simnet_tvar_53[5][21] , 
	\_zy_simnet_tvar_53[5][20] , \_zy_simnet_tvar_53[5][19] , 
	\_zy_simnet_tvar_53[5][18] , \_zy_simnet_tvar_53[5][17] , 
	\_zy_simnet_tvar_53[5][16] , \_zy_simnet_tvar_53[5][15] , 
	\_zy_simnet_tvar_53[5][14] , \_zy_simnet_tvar_53[5][13] , 
	\_zy_simnet_tvar_53[5][12] , \_zy_simnet_tvar_53[5][11] , 
	\_zy_simnet_tvar_53[5][10] , \_zy_simnet_tvar_53[5][9] , 
	\_zy_simnet_tvar_53[5][8] , \_zy_simnet_tvar_53[5][7] , 
	\_zy_simnet_tvar_53[5][6] , \_zy_simnet_tvar_53[5][5] , 
	\_zy_simnet_tvar_53[5][4] , \_zy_simnet_tvar_53[5][3] , 
	\_zy_simnet_tvar_53[5][2] , \_zy_simnet_tvar_53[5][1] , 
	\_zy_simnet_tvar_53[5][0] , \_zy_simnet_tvar_53[4][271] , 
	\_zy_simnet_tvar_53[4][270] , \_zy_simnet_tvar_53[4][269] , 
	\_zy_simnet_tvar_53[4][268] , \_zy_simnet_tvar_53[4][267] , 
	\_zy_simnet_tvar_53[4][266] , \_zy_simnet_tvar_53[4][265] , 
	\_zy_simnet_tvar_53[4][264] , \_zy_simnet_tvar_53[4][263] , 
	\_zy_simnet_tvar_53[4][262] , \_zy_simnet_tvar_53[4][261] , 
	\_zy_simnet_tvar_53[4][260] , \_zy_simnet_tvar_53[4][259] , 
	\_zy_simnet_tvar_53[4][258] , \_zy_simnet_tvar_53[4][257] , 
	\_zy_simnet_tvar_53[4][256] , \_zy_simnet_tvar_53[4][255] , 
	\_zy_simnet_tvar_53[4][254] , \_zy_simnet_tvar_53[4][253] , 
	\_zy_simnet_tvar_53[4][252] , \_zy_simnet_tvar_53[4][251] , 
	\_zy_simnet_tvar_53[4][250] , \_zy_simnet_tvar_53[4][249] , 
	\_zy_simnet_tvar_53[4][248] , \_zy_simnet_tvar_53[4][247] , 
	\_zy_simnet_tvar_53[4][246] , \_zy_simnet_tvar_53[4][245] , 
	\_zy_simnet_tvar_53[4][244] , \_zy_simnet_tvar_53[4][243] , 
	\_zy_simnet_tvar_53[4][242] , \_zy_simnet_tvar_53[4][241] , 
	\_zy_simnet_tvar_53[4][240] , \_zy_simnet_tvar_53[4][239] , 
	\_zy_simnet_tvar_53[4][238] , \_zy_simnet_tvar_53[4][237] , 
	\_zy_simnet_tvar_53[4][236] , \_zy_simnet_tvar_53[4][235] , 
	\_zy_simnet_tvar_53[4][234] , \_zy_simnet_tvar_53[4][233] , 
	\_zy_simnet_tvar_53[4][232] , \_zy_simnet_tvar_53[4][231] , 
	\_zy_simnet_tvar_53[4][230] , \_zy_simnet_tvar_53[4][229] , 
	\_zy_simnet_tvar_53[4][228] , \_zy_simnet_tvar_53[4][227] , 
	\_zy_simnet_tvar_53[4][226] , \_zy_simnet_tvar_53[4][225] , 
	\_zy_simnet_tvar_53[4][224] , \_zy_simnet_tvar_53[4][223] , 
	\_zy_simnet_tvar_53[4][222] , \_zy_simnet_tvar_53[4][221] , 
	\_zy_simnet_tvar_53[4][220] , \_zy_simnet_tvar_53[4][219] , 
	\_zy_simnet_tvar_53[4][218] , \_zy_simnet_tvar_53[4][217] , 
	\_zy_simnet_tvar_53[4][216] , \_zy_simnet_tvar_53[4][215] , 
	\_zy_simnet_tvar_53[4][214] , \_zy_simnet_tvar_53[4][213] , 
	\_zy_simnet_tvar_53[4][212] , \_zy_simnet_tvar_53[4][211] , 
	\_zy_simnet_tvar_53[4][210] , \_zy_simnet_tvar_53[4][209] , 
	\_zy_simnet_tvar_53[4][208] , \_zy_simnet_tvar_53[4][207] , 
	\_zy_simnet_tvar_53[4][206] , \_zy_simnet_tvar_53[4][205] , 
	\_zy_simnet_tvar_53[4][204] , \_zy_simnet_tvar_53[4][203] , 
	\_zy_simnet_tvar_53[4][202] , \_zy_simnet_tvar_53[4][201] , 
	\_zy_simnet_tvar_53[4][200] , \_zy_simnet_tvar_53[4][199] , 
	\_zy_simnet_tvar_53[4][198] , \_zy_simnet_tvar_53[4][197] , 
	\_zy_simnet_tvar_53[4][196] , \_zy_simnet_tvar_53[4][195] , 
	\_zy_simnet_tvar_53[4][194] , \_zy_simnet_tvar_53[4][193] , 
	\_zy_simnet_tvar_53[4][192] , \_zy_simnet_tvar_53[4][191] , 
	\_zy_simnet_tvar_53[4][190] , \_zy_simnet_tvar_53[4][189] , 
	\_zy_simnet_tvar_53[4][188] , \_zy_simnet_tvar_53[4][187] , 
	\_zy_simnet_tvar_53[4][186] , \_zy_simnet_tvar_53[4][185] , 
	\_zy_simnet_tvar_53[4][184] , \_zy_simnet_tvar_53[4][183] , 
	\_zy_simnet_tvar_53[4][182] , \_zy_simnet_tvar_53[4][181] , 
	\_zy_simnet_tvar_53[4][180] , \_zy_simnet_tvar_53[4][179] , 
	\_zy_simnet_tvar_53[4][178] , \_zy_simnet_tvar_53[4][177] , 
	\_zy_simnet_tvar_53[4][176] , \_zy_simnet_tvar_53[4][175] , 
	\_zy_simnet_tvar_53[4][174] , \_zy_simnet_tvar_53[4][173] , 
	\_zy_simnet_tvar_53[4][172] , \_zy_simnet_tvar_53[4][171] , 
	\_zy_simnet_tvar_53[4][170] , \_zy_simnet_tvar_53[4][169] , 
	\_zy_simnet_tvar_53[4][168] , \_zy_simnet_tvar_53[4][167] , 
	\_zy_simnet_tvar_53[4][166] , \_zy_simnet_tvar_53[4][165] , 
	\_zy_simnet_tvar_53[4][164] , \_zy_simnet_tvar_53[4][163] , 
	\_zy_simnet_tvar_53[4][162] , \_zy_simnet_tvar_53[4][161] , 
	\_zy_simnet_tvar_53[4][160] , \_zy_simnet_tvar_53[4][159] , 
	\_zy_simnet_tvar_53[4][158] , \_zy_simnet_tvar_53[4][157] , 
	\_zy_simnet_tvar_53[4][156] , \_zy_simnet_tvar_53[4][155] , 
	\_zy_simnet_tvar_53[4][154] , \_zy_simnet_tvar_53[4][153] , 
	\_zy_simnet_tvar_53[4][152] , \_zy_simnet_tvar_53[4][151] , 
	\_zy_simnet_tvar_53[4][150] , \_zy_simnet_tvar_53[4][149] , 
	\_zy_simnet_tvar_53[4][148] , \_zy_simnet_tvar_53[4][147] , 
	\_zy_simnet_tvar_53[4][146] , \_zy_simnet_tvar_53[4][145] , 
	\_zy_simnet_tvar_53[4][144] , \_zy_simnet_tvar_53[4][143] , 
	\_zy_simnet_tvar_53[4][142] , \_zy_simnet_tvar_53[4][141] , 
	\_zy_simnet_tvar_53[4][140] , \_zy_simnet_tvar_53[4][139] , 
	\_zy_simnet_tvar_53[4][138] , \_zy_simnet_tvar_53[4][137] , 
	\_zy_simnet_tvar_53[4][136] , \_zy_simnet_tvar_53[4][135] , 
	\_zy_simnet_tvar_53[4][134] , \_zy_simnet_tvar_53[4][133] , 
	\_zy_simnet_tvar_53[4][132] , \_zy_simnet_tvar_53[4][131] , 
	\_zy_simnet_tvar_53[4][130] , \_zy_simnet_tvar_53[4][129] , 
	\_zy_simnet_tvar_53[4][128] , \_zy_simnet_tvar_53[4][127] , 
	\_zy_simnet_tvar_53[4][126] , \_zy_simnet_tvar_53[4][125] , 
	\_zy_simnet_tvar_53[4][124] , \_zy_simnet_tvar_53[4][123] , 
	\_zy_simnet_tvar_53[4][122] , \_zy_simnet_tvar_53[4][121] , 
	\_zy_simnet_tvar_53[4][120] , \_zy_simnet_tvar_53[4][119] , 
	\_zy_simnet_tvar_53[4][118] , \_zy_simnet_tvar_53[4][117] , 
	\_zy_simnet_tvar_53[4][116] , \_zy_simnet_tvar_53[4][115] , 
	\_zy_simnet_tvar_53[4][114] , \_zy_simnet_tvar_53[4][113] , 
	\_zy_simnet_tvar_53[4][112] , \_zy_simnet_tvar_53[4][111] , 
	\_zy_simnet_tvar_53[4][110] , \_zy_simnet_tvar_53[4][109] , 
	\_zy_simnet_tvar_53[4][108] , \_zy_simnet_tvar_53[4][107] , 
	\_zy_simnet_tvar_53[4][106] , \_zy_simnet_tvar_53[4][105] , 
	\_zy_simnet_tvar_53[4][104] , \_zy_simnet_tvar_53[4][103] , 
	\_zy_simnet_tvar_53[4][102] , \_zy_simnet_tvar_53[4][101] , 
	\_zy_simnet_tvar_53[4][100] , \_zy_simnet_tvar_53[4][99] , 
	\_zy_simnet_tvar_53[4][98] , \_zy_simnet_tvar_53[4][97] , 
	\_zy_simnet_tvar_53[4][96] , \_zy_simnet_tvar_53[4][95] , 
	\_zy_simnet_tvar_53[4][94] , \_zy_simnet_tvar_53[4][93] , 
	\_zy_simnet_tvar_53[4][92] , \_zy_simnet_tvar_53[4][91] , 
	\_zy_simnet_tvar_53[4][90] , \_zy_simnet_tvar_53[4][89] , 
	\_zy_simnet_tvar_53[4][88] , \_zy_simnet_tvar_53[4][87] , 
	\_zy_simnet_tvar_53[4][86] , \_zy_simnet_tvar_53[4][85] , 
	\_zy_simnet_tvar_53[4][84] , \_zy_simnet_tvar_53[4][83] , 
	\_zy_simnet_tvar_53[4][82] , \_zy_simnet_tvar_53[4][81] , 
	\_zy_simnet_tvar_53[4][80] , \_zy_simnet_tvar_53[4][79] , 
	\_zy_simnet_tvar_53[4][78] , \_zy_simnet_tvar_53[4][77] , 
	\_zy_simnet_tvar_53[4][76] , \_zy_simnet_tvar_53[4][75] , 
	\_zy_simnet_tvar_53[4][74] , \_zy_simnet_tvar_53[4][73] , 
	\_zy_simnet_tvar_53[4][72] , \_zy_simnet_tvar_53[4][71] , 
	\_zy_simnet_tvar_53[4][70] , \_zy_simnet_tvar_53[4][69] , 
	\_zy_simnet_tvar_53[4][68] , \_zy_simnet_tvar_53[4][67] , 
	\_zy_simnet_tvar_53[4][66] , \_zy_simnet_tvar_53[4][65] , 
	\_zy_simnet_tvar_53[4][64] , \_zy_simnet_tvar_53[4][63] , 
	\_zy_simnet_tvar_53[4][62] , \_zy_simnet_tvar_53[4][61] , 
	\_zy_simnet_tvar_53[4][60] , \_zy_simnet_tvar_53[4][59] , 
	\_zy_simnet_tvar_53[4][58] , \_zy_simnet_tvar_53[4][57] , 
	\_zy_simnet_tvar_53[4][56] , \_zy_simnet_tvar_53[4][55] , 
	\_zy_simnet_tvar_53[4][54] , \_zy_simnet_tvar_53[4][53] , 
	\_zy_simnet_tvar_53[4][52] , \_zy_simnet_tvar_53[4][51] , 
	\_zy_simnet_tvar_53[4][50] , \_zy_simnet_tvar_53[4][49] , 
	\_zy_simnet_tvar_53[4][48] , \_zy_simnet_tvar_53[4][47] , 
	\_zy_simnet_tvar_53[4][46] , \_zy_simnet_tvar_53[4][45] , 
	\_zy_simnet_tvar_53[4][44] , \_zy_simnet_tvar_53[4][43] , 
	\_zy_simnet_tvar_53[4][42] , \_zy_simnet_tvar_53[4][41] , 
	\_zy_simnet_tvar_53[4][40] , \_zy_simnet_tvar_53[4][39] , 
	\_zy_simnet_tvar_53[4][38] , \_zy_simnet_tvar_53[4][37] , 
	\_zy_simnet_tvar_53[4][36] , \_zy_simnet_tvar_53[4][35] , 
	\_zy_simnet_tvar_53[4][34] , \_zy_simnet_tvar_53[4][33] , 
	\_zy_simnet_tvar_53[4][32] , \_zy_simnet_tvar_53[4][31] , 
	\_zy_simnet_tvar_53[4][30] , \_zy_simnet_tvar_53[4][29] , 
	\_zy_simnet_tvar_53[4][28] , \_zy_simnet_tvar_53[4][27] , 
	\_zy_simnet_tvar_53[4][26] , \_zy_simnet_tvar_53[4][25] , 
	\_zy_simnet_tvar_53[4][24] , \_zy_simnet_tvar_53[4][23] , 
	\_zy_simnet_tvar_53[4][22] , \_zy_simnet_tvar_53[4][21] , 
	\_zy_simnet_tvar_53[4][20] , \_zy_simnet_tvar_53[4][19] , 
	\_zy_simnet_tvar_53[4][18] , \_zy_simnet_tvar_53[4][17] , 
	\_zy_simnet_tvar_53[4][16] , \_zy_simnet_tvar_53[4][15] , 
	\_zy_simnet_tvar_53[4][14] , \_zy_simnet_tvar_53[4][13] , 
	\_zy_simnet_tvar_53[4][12] , \_zy_simnet_tvar_53[4][11] , 
	\_zy_simnet_tvar_53[4][10] , \_zy_simnet_tvar_53[4][9] , 
	\_zy_simnet_tvar_53[4][8] , \_zy_simnet_tvar_53[4][7] , 
	\_zy_simnet_tvar_53[4][6] , \_zy_simnet_tvar_53[4][5] , 
	\_zy_simnet_tvar_53[4][4] , \_zy_simnet_tvar_53[4][3] , 
	\_zy_simnet_tvar_53[4][2] , \_zy_simnet_tvar_53[4][1] , 
	\_zy_simnet_tvar_53[4][0] , \_zy_simnet_tvar_53[3][271] , 
	\_zy_simnet_tvar_53[3][270] , \_zy_simnet_tvar_53[3][269] , 
	\_zy_simnet_tvar_53[3][268] , \_zy_simnet_tvar_53[3][267] , 
	\_zy_simnet_tvar_53[3][266] , \_zy_simnet_tvar_53[3][265] , 
	\_zy_simnet_tvar_53[3][264] , \_zy_simnet_tvar_53[3][263] , 
	\_zy_simnet_tvar_53[3][262] , \_zy_simnet_tvar_53[3][261] , 
	\_zy_simnet_tvar_53[3][260] , \_zy_simnet_tvar_53[3][259] , 
	\_zy_simnet_tvar_53[3][258] , \_zy_simnet_tvar_53[3][257] , 
	\_zy_simnet_tvar_53[3][256] , \_zy_simnet_tvar_53[3][255] , 
	\_zy_simnet_tvar_53[3][254] , \_zy_simnet_tvar_53[3][253] , 
	\_zy_simnet_tvar_53[3][252] , \_zy_simnet_tvar_53[3][251] , 
	\_zy_simnet_tvar_53[3][250] , \_zy_simnet_tvar_53[3][249] , 
	\_zy_simnet_tvar_53[3][248] , \_zy_simnet_tvar_53[3][247] , 
	\_zy_simnet_tvar_53[3][246] , \_zy_simnet_tvar_53[3][245] , 
	\_zy_simnet_tvar_53[3][244] , \_zy_simnet_tvar_53[3][243] , 
	\_zy_simnet_tvar_53[3][242] , \_zy_simnet_tvar_53[3][241] , 
	\_zy_simnet_tvar_53[3][240] , \_zy_simnet_tvar_53[3][239] , 
	\_zy_simnet_tvar_53[3][238] , \_zy_simnet_tvar_53[3][237] , 
	\_zy_simnet_tvar_53[3][236] , \_zy_simnet_tvar_53[3][235] , 
	\_zy_simnet_tvar_53[3][234] , \_zy_simnet_tvar_53[3][233] , 
	\_zy_simnet_tvar_53[3][232] , \_zy_simnet_tvar_53[3][231] , 
	\_zy_simnet_tvar_53[3][230] , \_zy_simnet_tvar_53[3][229] , 
	\_zy_simnet_tvar_53[3][228] , \_zy_simnet_tvar_53[3][227] , 
	\_zy_simnet_tvar_53[3][226] , \_zy_simnet_tvar_53[3][225] , 
	\_zy_simnet_tvar_53[3][224] , \_zy_simnet_tvar_53[3][223] , 
	\_zy_simnet_tvar_53[3][222] , \_zy_simnet_tvar_53[3][221] , 
	\_zy_simnet_tvar_53[3][220] , \_zy_simnet_tvar_53[3][219] , 
	\_zy_simnet_tvar_53[3][218] , \_zy_simnet_tvar_53[3][217] , 
	\_zy_simnet_tvar_53[3][216] , \_zy_simnet_tvar_53[3][215] , 
	\_zy_simnet_tvar_53[3][214] , \_zy_simnet_tvar_53[3][213] , 
	\_zy_simnet_tvar_53[3][212] , \_zy_simnet_tvar_53[3][211] , 
	\_zy_simnet_tvar_53[3][210] , \_zy_simnet_tvar_53[3][209] , 
	\_zy_simnet_tvar_53[3][208] , \_zy_simnet_tvar_53[3][207] , 
	\_zy_simnet_tvar_53[3][206] , \_zy_simnet_tvar_53[3][205] , 
	\_zy_simnet_tvar_53[3][204] , \_zy_simnet_tvar_53[3][203] , 
	\_zy_simnet_tvar_53[3][202] , \_zy_simnet_tvar_53[3][201] , 
	\_zy_simnet_tvar_53[3][200] , \_zy_simnet_tvar_53[3][199] , 
	\_zy_simnet_tvar_53[3][198] , \_zy_simnet_tvar_53[3][197] , 
	\_zy_simnet_tvar_53[3][196] , \_zy_simnet_tvar_53[3][195] , 
	\_zy_simnet_tvar_53[3][194] , \_zy_simnet_tvar_53[3][193] , 
	\_zy_simnet_tvar_53[3][192] , \_zy_simnet_tvar_53[3][191] , 
	\_zy_simnet_tvar_53[3][190] , \_zy_simnet_tvar_53[3][189] , 
	\_zy_simnet_tvar_53[3][188] , \_zy_simnet_tvar_53[3][187] , 
	\_zy_simnet_tvar_53[3][186] , \_zy_simnet_tvar_53[3][185] , 
	\_zy_simnet_tvar_53[3][184] , \_zy_simnet_tvar_53[3][183] , 
	\_zy_simnet_tvar_53[3][182] , \_zy_simnet_tvar_53[3][181] , 
	\_zy_simnet_tvar_53[3][180] , \_zy_simnet_tvar_53[3][179] , 
	\_zy_simnet_tvar_53[3][178] , \_zy_simnet_tvar_53[3][177] , 
	\_zy_simnet_tvar_53[3][176] , \_zy_simnet_tvar_53[3][175] , 
	\_zy_simnet_tvar_53[3][174] , \_zy_simnet_tvar_53[3][173] , 
	\_zy_simnet_tvar_53[3][172] , \_zy_simnet_tvar_53[3][171] , 
	\_zy_simnet_tvar_53[3][170] , \_zy_simnet_tvar_53[3][169] , 
	\_zy_simnet_tvar_53[3][168] , \_zy_simnet_tvar_53[3][167] , 
	\_zy_simnet_tvar_53[3][166] , \_zy_simnet_tvar_53[3][165] , 
	\_zy_simnet_tvar_53[3][164] , \_zy_simnet_tvar_53[3][163] , 
	\_zy_simnet_tvar_53[3][162] , \_zy_simnet_tvar_53[3][161] , 
	\_zy_simnet_tvar_53[3][160] , \_zy_simnet_tvar_53[3][159] , 
	\_zy_simnet_tvar_53[3][158] , \_zy_simnet_tvar_53[3][157] , 
	\_zy_simnet_tvar_53[3][156] , \_zy_simnet_tvar_53[3][155] , 
	\_zy_simnet_tvar_53[3][154] , \_zy_simnet_tvar_53[3][153] , 
	\_zy_simnet_tvar_53[3][152] , \_zy_simnet_tvar_53[3][151] , 
	\_zy_simnet_tvar_53[3][150] , \_zy_simnet_tvar_53[3][149] , 
	\_zy_simnet_tvar_53[3][148] , \_zy_simnet_tvar_53[3][147] , 
	\_zy_simnet_tvar_53[3][146] , \_zy_simnet_tvar_53[3][145] , 
	\_zy_simnet_tvar_53[3][144] , \_zy_simnet_tvar_53[3][143] , 
	\_zy_simnet_tvar_53[3][142] , \_zy_simnet_tvar_53[3][141] , 
	\_zy_simnet_tvar_53[3][140] , \_zy_simnet_tvar_53[3][139] , 
	\_zy_simnet_tvar_53[3][138] , \_zy_simnet_tvar_53[3][137] , 
	\_zy_simnet_tvar_53[3][136] , \_zy_simnet_tvar_53[3][135] , 
	\_zy_simnet_tvar_53[3][134] , \_zy_simnet_tvar_53[3][133] , 
	\_zy_simnet_tvar_53[3][132] , \_zy_simnet_tvar_53[3][131] , 
	\_zy_simnet_tvar_53[3][130] , \_zy_simnet_tvar_53[3][129] , 
	\_zy_simnet_tvar_53[3][128] , \_zy_simnet_tvar_53[3][127] , 
	\_zy_simnet_tvar_53[3][126] , \_zy_simnet_tvar_53[3][125] , 
	\_zy_simnet_tvar_53[3][124] , \_zy_simnet_tvar_53[3][123] , 
	\_zy_simnet_tvar_53[3][122] , \_zy_simnet_tvar_53[3][121] , 
	\_zy_simnet_tvar_53[3][120] , \_zy_simnet_tvar_53[3][119] , 
	\_zy_simnet_tvar_53[3][118] , \_zy_simnet_tvar_53[3][117] , 
	\_zy_simnet_tvar_53[3][116] , \_zy_simnet_tvar_53[3][115] , 
	\_zy_simnet_tvar_53[3][114] , \_zy_simnet_tvar_53[3][113] , 
	\_zy_simnet_tvar_53[3][112] , \_zy_simnet_tvar_53[3][111] , 
	\_zy_simnet_tvar_53[3][110] , \_zy_simnet_tvar_53[3][109] , 
	\_zy_simnet_tvar_53[3][108] , \_zy_simnet_tvar_53[3][107] , 
	\_zy_simnet_tvar_53[3][106] , \_zy_simnet_tvar_53[3][105] , 
	\_zy_simnet_tvar_53[3][104] , \_zy_simnet_tvar_53[3][103] , 
	\_zy_simnet_tvar_53[3][102] , \_zy_simnet_tvar_53[3][101] , 
	\_zy_simnet_tvar_53[3][100] , \_zy_simnet_tvar_53[3][99] , 
	\_zy_simnet_tvar_53[3][98] , \_zy_simnet_tvar_53[3][97] , 
	\_zy_simnet_tvar_53[3][96] , \_zy_simnet_tvar_53[3][95] , 
	\_zy_simnet_tvar_53[3][94] , \_zy_simnet_tvar_53[3][93] , 
	\_zy_simnet_tvar_53[3][92] , \_zy_simnet_tvar_53[3][91] , 
	\_zy_simnet_tvar_53[3][90] , \_zy_simnet_tvar_53[3][89] , 
	\_zy_simnet_tvar_53[3][88] , \_zy_simnet_tvar_53[3][87] , 
	\_zy_simnet_tvar_53[3][86] , \_zy_simnet_tvar_53[3][85] , 
	\_zy_simnet_tvar_53[3][84] , \_zy_simnet_tvar_53[3][83] , 
	\_zy_simnet_tvar_53[3][82] , \_zy_simnet_tvar_53[3][81] , 
	\_zy_simnet_tvar_53[3][80] , \_zy_simnet_tvar_53[3][79] , 
	\_zy_simnet_tvar_53[3][78] , \_zy_simnet_tvar_53[3][77] , 
	\_zy_simnet_tvar_53[3][76] , \_zy_simnet_tvar_53[3][75] , 
	\_zy_simnet_tvar_53[3][74] , \_zy_simnet_tvar_53[3][73] , 
	\_zy_simnet_tvar_53[3][72] , \_zy_simnet_tvar_53[3][71] , 
	\_zy_simnet_tvar_53[3][70] , \_zy_simnet_tvar_53[3][69] , 
	\_zy_simnet_tvar_53[3][68] , \_zy_simnet_tvar_53[3][67] , 
	\_zy_simnet_tvar_53[3][66] , \_zy_simnet_tvar_53[3][65] , 
	\_zy_simnet_tvar_53[3][64] , \_zy_simnet_tvar_53[3][63] , 
	\_zy_simnet_tvar_53[3][62] , \_zy_simnet_tvar_53[3][61] , 
	\_zy_simnet_tvar_53[3][60] , \_zy_simnet_tvar_53[3][59] , 
	\_zy_simnet_tvar_53[3][58] , \_zy_simnet_tvar_53[3][57] , 
	\_zy_simnet_tvar_53[3][56] , \_zy_simnet_tvar_53[3][55] , 
	\_zy_simnet_tvar_53[3][54] , \_zy_simnet_tvar_53[3][53] , 
	\_zy_simnet_tvar_53[3][52] , \_zy_simnet_tvar_53[3][51] , 
	\_zy_simnet_tvar_53[3][50] , \_zy_simnet_tvar_53[3][49] , 
	\_zy_simnet_tvar_53[3][48] , \_zy_simnet_tvar_53[3][47] , 
	\_zy_simnet_tvar_53[3][46] , \_zy_simnet_tvar_53[3][45] , 
	\_zy_simnet_tvar_53[3][44] , \_zy_simnet_tvar_53[3][43] , 
	\_zy_simnet_tvar_53[3][42] , \_zy_simnet_tvar_53[3][41] , 
	\_zy_simnet_tvar_53[3][40] , \_zy_simnet_tvar_53[3][39] , 
	\_zy_simnet_tvar_53[3][38] , \_zy_simnet_tvar_53[3][37] , 
	\_zy_simnet_tvar_53[3][36] , \_zy_simnet_tvar_53[3][35] , 
	\_zy_simnet_tvar_53[3][34] , \_zy_simnet_tvar_53[3][33] , 
	\_zy_simnet_tvar_53[3][32] , \_zy_simnet_tvar_53[3][31] , 
	\_zy_simnet_tvar_53[3][30] , \_zy_simnet_tvar_53[3][29] , 
	\_zy_simnet_tvar_53[3][28] , \_zy_simnet_tvar_53[3][27] , 
	\_zy_simnet_tvar_53[3][26] , \_zy_simnet_tvar_53[3][25] , 
	\_zy_simnet_tvar_53[3][24] , \_zy_simnet_tvar_53[3][23] , 
	\_zy_simnet_tvar_53[3][22] , \_zy_simnet_tvar_53[3][21] , 
	\_zy_simnet_tvar_53[3][20] , \_zy_simnet_tvar_53[3][19] , 
	\_zy_simnet_tvar_53[3][18] , \_zy_simnet_tvar_53[3][17] , 
	\_zy_simnet_tvar_53[3][16] , \_zy_simnet_tvar_53[3][15] , 
	\_zy_simnet_tvar_53[3][14] , \_zy_simnet_tvar_53[3][13] , 
	\_zy_simnet_tvar_53[3][12] , \_zy_simnet_tvar_53[3][11] , 
	\_zy_simnet_tvar_53[3][10] , \_zy_simnet_tvar_53[3][9] , 
	\_zy_simnet_tvar_53[3][8] , \_zy_simnet_tvar_53[3][7] , 
	\_zy_simnet_tvar_53[3][6] , \_zy_simnet_tvar_53[3][5] , 
	\_zy_simnet_tvar_53[3][4] , \_zy_simnet_tvar_53[3][3] , 
	\_zy_simnet_tvar_53[3][2] , \_zy_simnet_tvar_53[3][1] , 
	\_zy_simnet_tvar_53[3][0] , \_zy_simnet_tvar_53[2][271] , 
	\_zy_simnet_tvar_53[2][270] , \_zy_simnet_tvar_53[2][269] , 
	\_zy_simnet_tvar_53[2][268] , \_zy_simnet_tvar_53[2][267] , 
	\_zy_simnet_tvar_53[2][266] , \_zy_simnet_tvar_53[2][265] , 
	\_zy_simnet_tvar_53[2][264] , \_zy_simnet_tvar_53[2][263] , 
	\_zy_simnet_tvar_53[2][262] , \_zy_simnet_tvar_53[2][261] , 
	\_zy_simnet_tvar_53[2][260] , \_zy_simnet_tvar_53[2][259] , 
	\_zy_simnet_tvar_53[2][258] , \_zy_simnet_tvar_53[2][257] , 
	\_zy_simnet_tvar_53[2][256] , \_zy_simnet_tvar_53[2][255] , 
	\_zy_simnet_tvar_53[2][254] , \_zy_simnet_tvar_53[2][253] , 
	\_zy_simnet_tvar_53[2][252] , \_zy_simnet_tvar_53[2][251] , 
	\_zy_simnet_tvar_53[2][250] , \_zy_simnet_tvar_53[2][249] , 
	\_zy_simnet_tvar_53[2][248] , \_zy_simnet_tvar_53[2][247] , 
	\_zy_simnet_tvar_53[2][246] , \_zy_simnet_tvar_53[2][245] , 
	\_zy_simnet_tvar_53[2][244] , \_zy_simnet_tvar_53[2][243] , 
	\_zy_simnet_tvar_53[2][242] , \_zy_simnet_tvar_53[2][241] , 
	\_zy_simnet_tvar_53[2][240] , \_zy_simnet_tvar_53[2][239] , 
	\_zy_simnet_tvar_53[2][238] , \_zy_simnet_tvar_53[2][237] , 
	\_zy_simnet_tvar_53[2][236] , \_zy_simnet_tvar_53[2][235] , 
	\_zy_simnet_tvar_53[2][234] , \_zy_simnet_tvar_53[2][233] , 
	\_zy_simnet_tvar_53[2][232] , \_zy_simnet_tvar_53[2][231] , 
	\_zy_simnet_tvar_53[2][230] , \_zy_simnet_tvar_53[2][229] , 
	\_zy_simnet_tvar_53[2][228] , \_zy_simnet_tvar_53[2][227] , 
	\_zy_simnet_tvar_53[2][226] , \_zy_simnet_tvar_53[2][225] , 
	\_zy_simnet_tvar_53[2][224] , \_zy_simnet_tvar_53[2][223] , 
	\_zy_simnet_tvar_53[2][222] , \_zy_simnet_tvar_53[2][221] , 
	\_zy_simnet_tvar_53[2][220] , \_zy_simnet_tvar_53[2][219] , 
	\_zy_simnet_tvar_53[2][218] , \_zy_simnet_tvar_53[2][217] , 
	\_zy_simnet_tvar_53[2][216] , \_zy_simnet_tvar_53[2][215] , 
	\_zy_simnet_tvar_53[2][214] , \_zy_simnet_tvar_53[2][213] , 
	\_zy_simnet_tvar_53[2][212] , \_zy_simnet_tvar_53[2][211] , 
	\_zy_simnet_tvar_53[2][210] , \_zy_simnet_tvar_53[2][209] , 
	\_zy_simnet_tvar_53[2][208] , \_zy_simnet_tvar_53[2][207] , 
	\_zy_simnet_tvar_53[2][206] , \_zy_simnet_tvar_53[2][205] , 
	\_zy_simnet_tvar_53[2][204] , \_zy_simnet_tvar_53[2][203] , 
	\_zy_simnet_tvar_53[2][202] , \_zy_simnet_tvar_53[2][201] , 
	\_zy_simnet_tvar_53[2][200] , \_zy_simnet_tvar_53[2][199] , 
	\_zy_simnet_tvar_53[2][198] , \_zy_simnet_tvar_53[2][197] , 
	\_zy_simnet_tvar_53[2][196] , \_zy_simnet_tvar_53[2][195] , 
	\_zy_simnet_tvar_53[2][194] , \_zy_simnet_tvar_53[2][193] , 
	\_zy_simnet_tvar_53[2][192] , \_zy_simnet_tvar_53[2][191] , 
	\_zy_simnet_tvar_53[2][190] , \_zy_simnet_tvar_53[2][189] , 
	\_zy_simnet_tvar_53[2][188] , \_zy_simnet_tvar_53[2][187] , 
	\_zy_simnet_tvar_53[2][186] , \_zy_simnet_tvar_53[2][185] , 
	\_zy_simnet_tvar_53[2][184] , \_zy_simnet_tvar_53[2][183] , 
	\_zy_simnet_tvar_53[2][182] , \_zy_simnet_tvar_53[2][181] , 
	\_zy_simnet_tvar_53[2][180] , \_zy_simnet_tvar_53[2][179] , 
	\_zy_simnet_tvar_53[2][178] , \_zy_simnet_tvar_53[2][177] , 
	\_zy_simnet_tvar_53[2][176] , \_zy_simnet_tvar_53[2][175] , 
	\_zy_simnet_tvar_53[2][174] , \_zy_simnet_tvar_53[2][173] , 
	\_zy_simnet_tvar_53[2][172] , \_zy_simnet_tvar_53[2][171] , 
	\_zy_simnet_tvar_53[2][170] , \_zy_simnet_tvar_53[2][169] , 
	\_zy_simnet_tvar_53[2][168] , \_zy_simnet_tvar_53[2][167] , 
	\_zy_simnet_tvar_53[2][166] , \_zy_simnet_tvar_53[2][165] , 
	\_zy_simnet_tvar_53[2][164] , \_zy_simnet_tvar_53[2][163] , 
	\_zy_simnet_tvar_53[2][162] , \_zy_simnet_tvar_53[2][161] , 
	\_zy_simnet_tvar_53[2][160] , \_zy_simnet_tvar_53[2][159] , 
	\_zy_simnet_tvar_53[2][158] , \_zy_simnet_tvar_53[2][157] , 
	\_zy_simnet_tvar_53[2][156] , \_zy_simnet_tvar_53[2][155] , 
	\_zy_simnet_tvar_53[2][154] , \_zy_simnet_tvar_53[2][153] , 
	\_zy_simnet_tvar_53[2][152] , \_zy_simnet_tvar_53[2][151] , 
	\_zy_simnet_tvar_53[2][150] , \_zy_simnet_tvar_53[2][149] , 
	\_zy_simnet_tvar_53[2][148] , \_zy_simnet_tvar_53[2][147] , 
	\_zy_simnet_tvar_53[2][146] , \_zy_simnet_tvar_53[2][145] , 
	\_zy_simnet_tvar_53[2][144] , \_zy_simnet_tvar_53[2][143] , 
	\_zy_simnet_tvar_53[2][142] , \_zy_simnet_tvar_53[2][141] , 
	\_zy_simnet_tvar_53[2][140] , \_zy_simnet_tvar_53[2][139] , 
	\_zy_simnet_tvar_53[2][138] , \_zy_simnet_tvar_53[2][137] , 
	\_zy_simnet_tvar_53[2][136] , \_zy_simnet_tvar_53[2][135] , 
	\_zy_simnet_tvar_53[2][134] , \_zy_simnet_tvar_53[2][133] , 
	\_zy_simnet_tvar_53[2][132] , \_zy_simnet_tvar_53[2][131] , 
	\_zy_simnet_tvar_53[2][130] , \_zy_simnet_tvar_53[2][129] , 
	\_zy_simnet_tvar_53[2][128] , \_zy_simnet_tvar_53[2][127] , 
	\_zy_simnet_tvar_53[2][126] , \_zy_simnet_tvar_53[2][125] , 
	\_zy_simnet_tvar_53[2][124] , \_zy_simnet_tvar_53[2][123] , 
	\_zy_simnet_tvar_53[2][122] , \_zy_simnet_tvar_53[2][121] , 
	\_zy_simnet_tvar_53[2][120] , \_zy_simnet_tvar_53[2][119] , 
	\_zy_simnet_tvar_53[2][118] , \_zy_simnet_tvar_53[2][117] , 
	\_zy_simnet_tvar_53[2][116] , \_zy_simnet_tvar_53[2][115] , 
	\_zy_simnet_tvar_53[2][114] , \_zy_simnet_tvar_53[2][113] , 
	\_zy_simnet_tvar_53[2][112] , \_zy_simnet_tvar_53[2][111] , 
	\_zy_simnet_tvar_53[2][110] , \_zy_simnet_tvar_53[2][109] , 
	\_zy_simnet_tvar_53[2][108] , \_zy_simnet_tvar_53[2][107] , 
	\_zy_simnet_tvar_53[2][106] , \_zy_simnet_tvar_53[2][105] , 
	\_zy_simnet_tvar_53[2][104] , \_zy_simnet_tvar_53[2][103] , 
	\_zy_simnet_tvar_53[2][102] , \_zy_simnet_tvar_53[2][101] , 
	\_zy_simnet_tvar_53[2][100] , \_zy_simnet_tvar_53[2][99] , 
	\_zy_simnet_tvar_53[2][98] , \_zy_simnet_tvar_53[2][97] , 
	\_zy_simnet_tvar_53[2][96] , \_zy_simnet_tvar_53[2][95] , 
	\_zy_simnet_tvar_53[2][94] , \_zy_simnet_tvar_53[2][93] , 
	\_zy_simnet_tvar_53[2][92] , \_zy_simnet_tvar_53[2][91] , 
	\_zy_simnet_tvar_53[2][90] , \_zy_simnet_tvar_53[2][89] , 
	\_zy_simnet_tvar_53[2][88] , \_zy_simnet_tvar_53[2][87] , 
	\_zy_simnet_tvar_53[2][86] , \_zy_simnet_tvar_53[2][85] , 
	\_zy_simnet_tvar_53[2][84] , \_zy_simnet_tvar_53[2][83] , 
	\_zy_simnet_tvar_53[2][82] , \_zy_simnet_tvar_53[2][81] , 
	\_zy_simnet_tvar_53[2][80] , \_zy_simnet_tvar_53[2][79] , 
	\_zy_simnet_tvar_53[2][78] , \_zy_simnet_tvar_53[2][77] , 
	\_zy_simnet_tvar_53[2][76] , \_zy_simnet_tvar_53[2][75] , 
	\_zy_simnet_tvar_53[2][74] , \_zy_simnet_tvar_53[2][73] , 
	\_zy_simnet_tvar_53[2][72] , \_zy_simnet_tvar_53[2][71] , 
	\_zy_simnet_tvar_53[2][70] , \_zy_simnet_tvar_53[2][69] , 
	\_zy_simnet_tvar_53[2][68] , \_zy_simnet_tvar_53[2][67] , 
	\_zy_simnet_tvar_53[2][66] , \_zy_simnet_tvar_53[2][65] , 
	\_zy_simnet_tvar_53[2][64] , \_zy_simnet_tvar_53[2][63] , 
	\_zy_simnet_tvar_53[2][62] , \_zy_simnet_tvar_53[2][61] , 
	\_zy_simnet_tvar_53[2][60] , \_zy_simnet_tvar_53[2][59] , 
	\_zy_simnet_tvar_53[2][58] , \_zy_simnet_tvar_53[2][57] , 
	\_zy_simnet_tvar_53[2][56] , \_zy_simnet_tvar_53[2][55] , 
	\_zy_simnet_tvar_53[2][54] , \_zy_simnet_tvar_53[2][53] , 
	\_zy_simnet_tvar_53[2][52] , \_zy_simnet_tvar_53[2][51] , 
	\_zy_simnet_tvar_53[2][50] , \_zy_simnet_tvar_53[2][49] , 
	\_zy_simnet_tvar_53[2][48] , \_zy_simnet_tvar_53[2][47] , 
	\_zy_simnet_tvar_53[2][46] , \_zy_simnet_tvar_53[2][45] , 
	\_zy_simnet_tvar_53[2][44] , \_zy_simnet_tvar_53[2][43] , 
	\_zy_simnet_tvar_53[2][42] , \_zy_simnet_tvar_53[2][41] , 
	\_zy_simnet_tvar_53[2][40] , \_zy_simnet_tvar_53[2][39] , 
	\_zy_simnet_tvar_53[2][38] , \_zy_simnet_tvar_53[2][37] , 
	\_zy_simnet_tvar_53[2][36] , \_zy_simnet_tvar_53[2][35] , 
	\_zy_simnet_tvar_53[2][34] , \_zy_simnet_tvar_53[2][33] , 
	\_zy_simnet_tvar_53[2][32] , \_zy_simnet_tvar_53[2][31] , 
	\_zy_simnet_tvar_53[2][30] , \_zy_simnet_tvar_53[2][29] , 
	\_zy_simnet_tvar_53[2][28] , \_zy_simnet_tvar_53[2][27] , 
	\_zy_simnet_tvar_53[2][26] , \_zy_simnet_tvar_53[2][25] , 
	\_zy_simnet_tvar_53[2][24] , \_zy_simnet_tvar_53[2][23] , 
	\_zy_simnet_tvar_53[2][22] , \_zy_simnet_tvar_53[2][21] , 
	\_zy_simnet_tvar_53[2][20] , \_zy_simnet_tvar_53[2][19] , 
	\_zy_simnet_tvar_53[2][18] , \_zy_simnet_tvar_53[2][17] , 
	\_zy_simnet_tvar_53[2][16] , \_zy_simnet_tvar_53[2][15] , 
	\_zy_simnet_tvar_53[2][14] , \_zy_simnet_tvar_53[2][13] , 
	\_zy_simnet_tvar_53[2][12] , \_zy_simnet_tvar_53[2][11] , 
	\_zy_simnet_tvar_53[2][10] , \_zy_simnet_tvar_53[2][9] , 
	\_zy_simnet_tvar_53[2][8] , \_zy_simnet_tvar_53[2][7] , 
	\_zy_simnet_tvar_53[2][6] , \_zy_simnet_tvar_53[2][5] , 
	\_zy_simnet_tvar_53[2][4] , \_zy_simnet_tvar_53[2][3] , 
	\_zy_simnet_tvar_53[2][2] , \_zy_simnet_tvar_53[2][1] , 
	\_zy_simnet_tvar_53[2][0] , \_zy_simnet_tvar_53[1][271] , 
	\_zy_simnet_tvar_53[1][270] , \_zy_simnet_tvar_53[1][269] , 
	\_zy_simnet_tvar_53[1][268] , \_zy_simnet_tvar_53[1][267] , 
	\_zy_simnet_tvar_53[1][266] , \_zy_simnet_tvar_53[1][265] , 
	\_zy_simnet_tvar_53[1][264] , \_zy_simnet_tvar_53[1][263] , 
	\_zy_simnet_tvar_53[1][262] , \_zy_simnet_tvar_53[1][261] , 
	\_zy_simnet_tvar_53[1][260] , \_zy_simnet_tvar_53[1][259] , 
	\_zy_simnet_tvar_53[1][258] , \_zy_simnet_tvar_53[1][257] , 
	\_zy_simnet_tvar_53[1][256] , \_zy_simnet_tvar_53[1][255] , 
	\_zy_simnet_tvar_53[1][254] , \_zy_simnet_tvar_53[1][253] , 
	\_zy_simnet_tvar_53[1][252] , \_zy_simnet_tvar_53[1][251] , 
	\_zy_simnet_tvar_53[1][250] , \_zy_simnet_tvar_53[1][249] , 
	\_zy_simnet_tvar_53[1][248] , \_zy_simnet_tvar_53[1][247] , 
	\_zy_simnet_tvar_53[1][246] , \_zy_simnet_tvar_53[1][245] , 
	\_zy_simnet_tvar_53[1][244] , \_zy_simnet_tvar_53[1][243] , 
	\_zy_simnet_tvar_53[1][242] , \_zy_simnet_tvar_53[1][241] , 
	\_zy_simnet_tvar_53[1][240] , \_zy_simnet_tvar_53[1][239] , 
	\_zy_simnet_tvar_53[1][238] , \_zy_simnet_tvar_53[1][237] , 
	\_zy_simnet_tvar_53[1][236] , \_zy_simnet_tvar_53[1][235] , 
	\_zy_simnet_tvar_53[1][234] , \_zy_simnet_tvar_53[1][233] , 
	\_zy_simnet_tvar_53[1][232] , \_zy_simnet_tvar_53[1][231] , 
	\_zy_simnet_tvar_53[1][230] , \_zy_simnet_tvar_53[1][229] , 
	\_zy_simnet_tvar_53[1][228] , \_zy_simnet_tvar_53[1][227] , 
	\_zy_simnet_tvar_53[1][226] , \_zy_simnet_tvar_53[1][225] , 
	\_zy_simnet_tvar_53[1][224] , \_zy_simnet_tvar_53[1][223] , 
	\_zy_simnet_tvar_53[1][222] , \_zy_simnet_tvar_53[1][221] , 
	\_zy_simnet_tvar_53[1][220] , \_zy_simnet_tvar_53[1][219] , 
	\_zy_simnet_tvar_53[1][218] , \_zy_simnet_tvar_53[1][217] , 
	\_zy_simnet_tvar_53[1][216] , \_zy_simnet_tvar_53[1][215] , 
	\_zy_simnet_tvar_53[1][214] , \_zy_simnet_tvar_53[1][213] , 
	\_zy_simnet_tvar_53[1][212] , \_zy_simnet_tvar_53[1][211] , 
	\_zy_simnet_tvar_53[1][210] , \_zy_simnet_tvar_53[1][209] , 
	\_zy_simnet_tvar_53[1][208] , \_zy_simnet_tvar_53[1][207] , 
	\_zy_simnet_tvar_53[1][206] , \_zy_simnet_tvar_53[1][205] , 
	\_zy_simnet_tvar_53[1][204] , \_zy_simnet_tvar_53[1][203] , 
	\_zy_simnet_tvar_53[1][202] , \_zy_simnet_tvar_53[1][201] , 
	\_zy_simnet_tvar_53[1][200] , \_zy_simnet_tvar_53[1][199] , 
	\_zy_simnet_tvar_53[1][198] , \_zy_simnet_tvar_53[1][197] , 
	\_zy_simnet_tvar_53[1][196] , \_zy_simnet_tvar_53[1][195] , 
	\_zy_simnet_tvar_53[1][194] , \_zy_simnet_tvar_53[1][193] , 
	\_zy_simnet_tvar_53[1][192] , \_zy_simnet_tvar_53[1][191] , 
	\_zy_simnet_tvar_53[1][190] , \_zy_simnet_tvar_53[1][189] , 
	\_zy_simnet_tvar_53[1][188] , \_zy_simnet_tvar_53[1][187] , 
	\_zy_simnet_tvar_53[1][186] , \_zy_simnet_tvar_53[1][185] , 
	\_zy_simnet_tvar_53[1][184] , \_zy_simnet_tvar_53[1][183] , 
	\_zy_simnet_tvar_53[1][182] , \_zy_simnet_tvar_53[1][181] , 
	\_zy_simnet_tvar_53[1][180] , \_zy_simnet_tvar_53[1][179] , 
	\_zy_simnet_tvar_53[1][178] , \_zy_simnet_tvar_53[1][177] , 
	\_zy_simnet_tvar_53[1][176] , \_zy_simnet_tvar_53[1][175] , 
	\_zy_simnet_tvar_53[1][174] , \_zy_simnet_tvar_53[1][173] , 
	\_zy_simnet_tvar_53[1][172] , \_zy_simnet_tvar_53[1][171] , 
	\_zy_simnet_tvar_53[1][170] , \_zy_simnet_tvar_53[1][169] , 
	\_zy_simnet_tvar_53[1][168] , \_zy_simnet_tvar_53[1][167] , 
	\_zy_simnet_tvar_53[1][166] , \_zy_simnet_tvar_53[1][165] , 
	\_zy_simnet_tvar_53[1][164] , \_zy_simnet_tvar_53[1][163] , 
	\_zy_simnet_tvar_53[1][162] , \_zy_simnet_tvar_53[1][161] , 
	\_zy_simnet_tvar_53[1][160] , \_zy_simnet_tvar_53[1][159] , 
	\_zy_simnet_tvar_53[1][158] , \_zy_simnet_tvar_53[1][157] , 
	\_zy_simnet_tvar_53[1][156] , \_zy_simnet_tvar_53[1][155] , 
	\_zy_simnet_tvar_53[1][154] , \_zy_simnet_tvar_53[1][153] , 
	\_zy_simnet_tvar_53[1][152] , \_zy_simnet_tvar_53[1][151] , 
	\_zy_simnet_tvar_53[1][150] , \_zy_simnet_tvar_53[1][149] , 
	\_zy_simnet_tvar_53[1][148] , \_zy_simnet_tvar_53[1][147] , 
	\_zy_simnet_tvar_53[1][146] , \_zy_simnet_tvar_53[1][145] , 
	\_zy_simnet_tvar_53[1][144] , \_zy_simnet_tvar_53[1][143] , 
	\_zy_simnet_tvar_53[1][142] , \_zy_simnet_tvar_53[1][141] , 
	\_zy_simnet_tvar_53[1][140] , \_zy_simnet_tvar_53[1][139] , 
	\_zy_simnet_tvar_53[1][138] , \_zy_simnet_tvar_53[1][137] , 
	\_zy_simnet_tvar_53[1][136] , \_zy_simnet_tvar_53[1][135] , 
	\_zy_simnet_tvar_53[1][134] , \_zy_simnet_tvar_53[1][133] , 
	\_zy_simnet_tvar_53[1][132] , \_zy_simnet_tvar_53[1][131] , 
	\_zy_simnet_tvar_53[1][130] , \_zy_simnet_tvar_53[1][129] , 
	\_zy_simnet_tvar_53[1][128] , \_zy_simnet_tvar_53[1][127] , 
	\_zy_simnet_tvar_53[1][126] , \_zy_simnet_tvar_53[1][125] , 
	\_zy_simnet_tvar_53[1][124] , \_zy_simnet_tvar_53[1][123] , 
	\_zy_simnet_tvar_53[1][122] , \_zy_simnet_tvar_53[1][121] , 
	\_zy_simnet_tvar_53[1][120] , \_zy_simnet_tvar_53[1][119] , 
	\_zy_simnet_tvar_53[1][118] , \_zy_simnet_tvar_53[1][117] , 
	\_zy_simnet_tvar_53[1][116] , \_zy_simnet_tvar_53[1][115] , 
	\_zy_simnet_tvar_53[1][114] , \_zy_simnet_tvar_53[1][113] , 
	\_zy_simnet_tvar_53[1][112] , \_zy_simnet_tvar_53[1][111] , 
	\_zy_simnet_tvar_53[1][110] , \_zy_simnet_tvar_53[1][109] , 
	\_zy_simnet_tvar_53[1][108] , \_zy_simnet_tvar_53[1][107] , 
	\_zy_simnet_tvar_53[1][106] , \_zy_simnet_tvar_53[1][105] , 
	\_zy_simnet_tvar_53[1][104] , \_zy_simnet_tvar_53[1][103] , 
	\_zy_simnet_tvar_53[1][102] , \_zy_simnet_tvar_53[1][101] , 
	\_zy_simnet_tvar_53[1][100] , \_zy_simnet_tvar_53[1][99] , 
	\_zy_simnet_tvar_53[1][98] , \_zy_simnet_tvar_53[1][97] , 
	\_zy_simnet_tvar_53[1][96] , \_zy_simnet_tvar_53[1][95] , 
	\_zy_simnet_tvar_53[1][94] , \_zy_simnet_tvar_53[1][93] , 
	\_zy_simnet_tvar_53[1][92] , \_zy_simnet_tvar_53[1][91] , 
	\_zy_simnet_tvar_53[1][90] , \_zy_simnet_tvar_53[1][89] , 
	\_zy_simnet_tvar_53[1][88] , \_zy_simnet_tvar_53[1][87] , 
	\_zy_simnet_tvar_53[1][86] , \_zy_simnet_tvar_53[1][85] , 
	\_zy_simnet_tvar_53[1][84] , \_zy_simnet_tvar_53[1][83] , 
	\_zy_simnet_tvar_53[1][82] , \_zy_simnet_tvar_53[1][81] , 
	\_zy_simnet_tvar_53[1][80] , \_zy_simnet_tvar_53[1][79] , 
	\_zy_simnet_tvar_53[1][78] , \_zy_simnet_tvar_53[1][77] , 
	\_zy_simnet_tvar_53[1][76] , \_zy_simnet_tvar_53[1][75] , 
	\_zy_simnet_tvar_53[1][74] , \_zy_simnet_tvar_53[1][73] , 
	\_zy_simnet_tvar_53[1][72] , \_zy_simnet_tvar_53[1][71] , 
	\_zy_simnet_tvar_53[1][70] , \_zy_simnet_tvar_53[1][69] , 
	\_zy_simnet_tvar_53[1][68] , \_zy_simnet_tvar_53[1][67] , 
	\_zy_simnet_tvar_53[1][66] , \_zy_simnet_tvar_53[1][65] , 
	\_zy_simnet_tvar_53[1][64] , \_zy_simnet_tvar_53[1][63] , 
	\_zy_simnet_tvar_53[1][62] , \_zy_simnet_tvar_53[1][61] , 
	\_zy_simnet_tvar_53[1][60] , \_zy_simnet_tvar_53[1][59] , 
	\_zy_simnet_tvar_53[1][58] , \_zy_simnet_tvar_53[1][57] , 
	\_zy_simnet_tvar_53[1][56] , \_zy_simnet_tvar_53[1][55] , 
	\_zy_simnet_tvar_53[1][54] , \_zy_simnet_tvar_53[1][53] , 
	\_zy_simnet_tvar_53[1][52] , \_zy_simnet_tvar_53[1][51] , 
	\_zy_simnet_tvar_53[1][50] , \_zy_simnet_tvar_53[1][49] , 
	\_zy_simnet_tvar_53[1][48] , \_zy_simnet_tvar_53[1][47] , 
	\_zy_simnet_tvar_53[1][46] , \_zy_simnet_tvar_53[1][45] , 
	\_zy_simnet_tvar_53[1][44] , \_zy_simnet_tvar_53[1][43] , 
	\_zy_simnet_tvar_53[1][42] , \_zy_simnet_tvar_53[1][41] , 
	\_zy_simnet_tvar_53[1][40] , \_zy_simnet_tvar_53[1][39] , 
	\_zy_simnet_tvar_53[1][38] , \_zy_simnet_tvar_53[1][37] , 
	\_zy_simnet_tvar_53[1][36] , \_zy_simnet_tvar_53[1][35] , 
	\_zy_simnet_tvar_53[1][34] , \_zy_simnet_tvar_53[1][33] , 
	\_zy_simnet_tvar_53[1][32] , \_zy_simnet_tvar_53[1][31] , 
	\_zy_simnet_tvar_53[1][30] , \_zy_simnet_tvar_53[1][29] , 
	\_zy_simnet_tvar_53[1][28] , \_zy_simnet_tvar_53[1][27] , 
	\_zy_simnet_tvar_53[1][26] , \_zy_simnet_tvar_53[1][25] , 
	\_zy_simnet_tvar_53[1][24] , \_zy_simnet_tvar_53[1][23] , 
	\_zy_simnet_tvar_53[1][22] , \_zy_simnet_tvar_53[1][21] , 
	\_zy_simnet_tvar_53[1][20] , \_zy_simnet_tvar_53[1][19] , 
	\_zy_simnet_tvar_53[1][18] , \_zy_simnet_tvar_53[1][17] , 
	\_zy_simnet_tvar_53[1][16] , \_zy_simnet_tvar_53[1][15] , 
	\_zy_simnet_tvar_53[1][14] , \_zy_simnet_tvar_53[1][13] , 
	\_zy_simnet_tvar_53[1][12] , \_zy_simnet_tvar_53[1][11] , 
	\_zy_simnet_tvar_53[1][10] , \_zy_simnet_tvar_53[1][9] , 
	\_zy_simnet_tvar_53[1][8] , \_zy_simnet_tvar_53[1][7] , 
	\_zy_simnet_tvar_53[1][6] , \_zy_simnet_tvar_53[1][5] , 
	\_zy_simnet_tvar_53[1][4] , \_zy_simnet_tvar_53[1][3] , 
	\_zy_simnet_tvar_53[1][2] , \_zy_simnet_tvar_53[1][1] , 
	\_zy_simnet_tvar_53[1][0] , \_zy_simnet_tvar_53[0][271] , 
	\_zy_simnet_tvar_53[0][270] , \_zy_simnet_tvar_53[0][269] , 
	\_zy_simnet_tvar_53[0][268] , \_zy_simnet_tvar_53[0][267] , 
	\_zy_simnet_tvar_53[0][266] , \_zy_simnet_tvar_53[0][265] , 
	\_zy_simnet_tvar_53[0][264] , \_zy_simnet_tvar_53[0][263] , 
	\_zy_simnet_tvar_53[0][262] , \_zy_simnet_tvar_53[0][261] , 
	\_zy_simnet_tvar_53[0][260] , \_zy_simnet_tvar_53[0][259] , 
	\_zy_simnet_tvar_53[0][258] , \_zy_simnet_tvar_53[0][257] , 
	\_zy_simnet_tvar_53[0][256] , \_zy_simnet_tvar_53[0][255] , 
	\_zy_simnet_tvar_53[0][254] , \_zy_simnet_tvar_53[0][253] , 
	\_zy_simnet_tvar_53[0][252] , \_zy_simnet_tvar_53[0][251] , 
	\_zy_simnet_tvar_53[0][250] , \_zy_simnet_tvar_53[0][249] , 
	\_zy_simnet_tvar_53[0][248] , \_zy_simnet_tvar_53[0][247] , 
	\_zy_simnet_tvar_53[0][246] , \_zy_simnet_tvar_53[0][245] , 
	\_zy_simnet_tvar_53[0][244] , \_zy_simnet_tvar_53[0][243] , 
	\_zy_simnet_tvar_53[0][242] , \_zy_simnet_tvar_53[0][241] , 
	\_zy_simnet_tvar_53[0][240] , \_zy_simnet_tvar_53[0][239] , 
	\_zy_simnet_tvar_53[0][238] , \_zy_simnet_tvar_53[0][237] , 
	\_zy_simnet_tvar_53[0][236] , \_zy_simnet_tvar_53[0][235] , 
	\_zy_simnet_tvar_53[0][234] , \_zy_simnet_tvar_53[0][233] , 
	\_zy_simnet_tvar_53[0][232] , \_zy_simnet_tvar_53[0][231] , 
	\_zy_simnet_tvar_53[0][230] , \_zy_simnet_tvar_53[0][229] , 
	\_zy_simnet_tvar_53[0][228] , \_zy_simnet_tvar_53[0][227] , 
	\_zy_simnet_tvar_53[0][226] , \_zy_simnet_tvar_53[0][225] , 
	\_zy_simnet_tvar_53[0][224] , \_zy_simnet_tvar_53[0][223] , 
	\_zy_simnet_tvar_53[0][222] , \_zy_simnet_tvar_53[0][221] , 
	\_zy_simnet_tvar_53[0][220] , \_zy_simnet_tvar_53[0][219] , 
	\_zy_simnet_tvar_53[0][218] , \_zy_simnet_tvar_53[0][217] , 
	\_zy_simnet_tvar_53[0][216] , \_zy_simnet_tvar_53[0][215] , 
	\_zy_simnet_tvar_53[0][214] , \_zy_simnet_tvar_53[0][213] , 
	\_zy_simnet_tvar_53[0][212] , \_zy_simnet_tvar_53[0][211] , 
	\_zy_simnet_tvar_53[0][210] , \_zy_simnet_tvar_53[0][209] , 
	\_zy_simnet_tvar_53[0][208] , \_zy_simnet_tvar_53[0][207] , 
	\_zy_simnet_tvar_53[0][206] , \_zy_simnet_tvar_53[0][205] , 
	\_zy_simnet_tvar_53[0][204] , \_zy_simnet_tvar_53[0][203] , 
	\_zy_simnet_tvar_53[0][202] , \_zy_simnet_tvar_53[0][201] , 
	\_zy_simnet_tvar_53[0][200] , \_zy_simnet_tvar_53[0][199] , 
	\_zy_simnet_tvar_53[0][198] , \_zy_simnet_tvar_53[0][197] , 
	\_zy_simnet_tvar_53[0][196] , \_zy_simnet_tvar_53[0][195] , 
	\_zy_simnet_tvar_53[0][194] , \_zy_simnet_tvar_53[0][193] , 
	\_zy_simnet_tvar_53[0][192] , \_zy_simnet_tvar_53[0][191] , 
	\_zy_simnet_tvar_53[0][190] , \_zy_simnet_tvar_53[0][189] , 
	\_zy_simnet_tvar_53[0][188] , \_zy_simnet_tvar_53[0][187] , 
	\_zy_simnet_tvar_53[0][186] , \_zy_simnet_tvar_53[0][185] , 
	\_zy_simnet_tvar_53[0][184] , \_zy_simnet_tvar_53[0][183] , 
	\_zy_simnet_tvar_53[0][182] , \_zy_simnet_tvar_53[0][181] , 
	\_zy_simnet_tvar_53[0][180] , \_zy_simnet_tvar_53[0][179] , 
	\_zy_simnet_tvar_53[0][178] , \_zy_simnet_tvar_53[0][177] , 
	\_zy_simnet_tvar_53[0][176] , \_zy_simnet_tvar_53[0][175] , 
	\_zy_simnet_tvar_53[0][174] , \_zy_simnet_tvar_53[0][173] , 
	\_zy_simnet_tvar_53[0][172] , \_zy_simnet_tvar_53[0][171] , 
	\_zy_simnet_tvar_53[0][170] , \_zy_simnet_tvar_53[0][169] , 
	\_zy_simnet_tvar_53[0][168] , \_zy_simnet_tvar_53[0][167] , 
	\_zy_simnet_tvar_53[0][166] , \_zy_simnet_tvar_53[0][165] , 
	\_zy_simnet_tvar_53[0][164] , \_zy_simnet_tvar_53[0][163] , 
	\_zy_simnet_tvar_53[0][162] , \_zy_simnet_tvar_53[0][161] , 
	\_zy_simnet_tvar_53[0][160] , \_zy_simnet_tvar_53[0][159] , 
	\_zy_simnet_tvar_53[0][158] , \_zy_simnet_tvar_53[0][157] , 
	\_zy_simnet_tvar_53[0][156] , \_zy_simnet_tvar_53[0][155] , 
	\_zy_simnet_tvar_53[0][154] , \_zy_simnet_tvar_53[0][153] , 
	\_zy_simnet_tvar_53[0][152] , \_zy_simnet_tvar_53[0][151] , 
	\_zy_simnet_tvar_53[0][150] , \_zy_simnet_tvar_53[0][149] , 
	\_zy_simnet_tvar_53[0][148] , \_zy_simnet_tvar_53[0][147] , 
	\_zy_simnet_tvar_53[0][146] , \_zy_simnet_tvar_53[0][145] , 
	\_zy_simnet_tvar_53[0][144] , \_zy_simnet_tvar_53[0][143] , 
	\_zy_simnet_tvar_53[0][142] , \_zy_simnet_tvar_53[0][141] , 
	\_zy_simnet_tvar_53[0][140] , \_zy_simnet_tvar_53[0][139] , 
	\_zy_simnet_tvar_53[0][138] , \_zy_simnet_tvar_53[0][137] , 
	\_zy_simnet_tvar_53[0][136] , \_zy_simnet_tvar_53[0][135] , 
	\_zy_simnet_tvar_53[0][134] , \_zy_simnet_tvar_53[0][133] , 
	\_zy_simnet_tvar_53[0][132] , \_zy_simnet_tvar_53[0][131] , 
	\_zy_simnet_tvar_53[0][130] , \_zy_simnet_tvar_53[0][129] , 
	\_zy_simnet_tvar_53[0][128] , \_zy_simnet_tvar_53[0][127] , 
	\_zy_simnet_tvar_53[0][126] , \_zy_simnet_tvar_53[0][125] , 
	\_zy_simnet_tvar_53[0][124] , \_zy_simnet_tvar_53[0][123] , 
	\_zy_simnet_tvar_53[0][122] , \_zy_simnet_tvar_53[0][121] , 
	\_zy_simnet_tvar_53[0][120] , \_zy_simnet_tvar_53[0][119] , 
	\_zy_simnet_tvar_53[0][118] , \_zy_simnet_tvar_53[0][117] , 
	\_zy_simnet_tvar_53[0][116] , \_zy_simnet_tvar_53[0][115] , 
	\_zy_simnet_tvar_53[0][114] , \_zy_simnet_tvar_53[0][113] , 
	\_zy_simnet_tvar_53[0][112] , \_zy_simnet_tvar_53[0][111] , 
	\_zy_simnet_tvar_53[0][110] , \_zy_simnet_tvar_53[0][109] , 
	\_zy_simnet_tvar_53[0][108] , \_zy_simnet_tvar_53[0][107] , 
	\_zy_simnet_tvar_53[0][106] , \_zy_simnet_tvar_53[0][105] , 
	\_zy_simnet_tvar_53[0][104] , \_zy_simnet_tvar_53[0][103] , 
	\_zy_simnet_tvar_53[0][102] , \_zy_simnet_tvar_53[0][101] , 
	\_zy_simnet_tvar_53[0][100] , \_zy_simnet_tvar_53[0][99] , 
	\_zy_simnet_tvar_53[0][98] , \_zy_simnet_tvar_53[0][97] , 
	\_zy_simnet_tvar_53[0][96] , \_zy_simnet_tvar_53[0][95] , 
	\_zy_simnet_tvar_53[0][94] , \_zy_simnet_tvar_53[0][93] , 
	\_zy_simnet_tvar_53[0][92] , \_zy_simnet_tvar_53[0][91] , 
	\_zy_simnet_tvar_53[0][90] , \_zy_simnet_tvar_53[0][89] , 
	\_zy_simnet_tvar_53[0][88] , \_zy_simnet_tvar_53[0][87] , 
	\_zy_simnet_tvar_53[0][86] , \_zy_simnet_tvar_53[0][85] , 
	\_zy_simnet_tvar_53[0][84] , \_zy_simnet_tvar_53[0][83] , 
	\_zy_simnet_tvar_53[0][82] , \_zy_simnet_tvar_53[0][81] , 
	\_zy_simnet_tvar_53[0][80] , \_zy_simnet_tvar_53[0][79] , 
	\_zy_simnet_tvar_53[0][78] , \_zy_simnet_tvar_53[0][77] , 
	\_zy_simnet_tvar_53[0][76] , \_zy_simnet_tvar_53[0][75] , 
	\_zy_simnet_tvar_53[0][74] , \_zy_simnet_tvar_53[0][73] , 
	\_zy_simnet_tvar_53[0][72] , \_zy_simnet_tvar_53[0][71] , 
	\_zy_simnet_tvar_53[0][70] , \_zy_simnet_tvar_53[0][69] , 
	\_zy_simnet_tvar_53[0][68] , \_zy_simnet_tvar_53[0][67] , 
	\_zy_simnet_tvar_53[0][66] , \_zy_simnet_tvar_53[0][65] , 
	\_zy_simnet_tvar_53[0][64] , \_zy_simnet_tvar_53[0][63] , 
	\_zy_simnet_tvar_53[0][62] , \_zy_simnet_tvar_53[0][61] , 
	\_zy_simnet_tvar_53[0][60] , \_zy_simnet_tvar_53[0][59] , 
	\_zy_simnet_tvar_53[0][58] , \_zy_simnet_tvar_53[0][57] , 
	\_zy_simnet_tvar_53[0][56] , \_zy_simnet_tvar_53[0][55] , 
	\_zy_simnet_tvar_53[0][54] , \_zy_simnet_tvar_53[0][53] , 
	\_zy_simnet_tvar_53[0][52] , \_zy_simnet_tvar_53[0][51] , 
	\_zy_simnet_tvar_53[0][50] , \_zy_simnet_tvar_53[0][49] , 
	\_zy_simnet_tvar_53[0][48] , \_zy_simnet_tvar_53[0][47] , 
	\_zy_simnet_tvar_53[0][46] , \_zy_simnet_tvar_53[0][45] , 
	\_zy_simnet_tvar_53[0][44] , \_zy_simnet_tvar_53[0][43] , 
	\_zy_simnet_tvar_53[0][42] , \_zy_simnet_tvar_53[0][41] , 
	\_zy_simnet_tvar_53[0][40] , \_zy_simnet_tvar_53[0][39] , 
	\_zy_simnet_tvar_53[0][38] , \_zy_simnet_tvar_53[0][37] , 
	\_zy_simnet_tvar_53[0][36] , \_zy_simnet_tvar_53[0][35] , 
	\_zy_simnet_tvar_53[0][34] , \_zy_simnet_tvar_53[0][33] , 
	\_zy_simnet_tvar_53[0][32] , \_zy_simnet_tvar_53[0][31] , 
	\_zy_simnet_tvar_53[0][30] , \_zy_simnet_tvar_53[0][29] , 
	\_zy_simnet_tvar_53[0][28] , \_zy_simnet_tvar_53[0][27] , 
	\_zy_simnet_tvar_53[0][26] , \_zy_simnet_tvar_53[0][25] , 
	\_zy_simnet_tvar_53[0][24] , \_zy_simnet_tvar_53[0][23] , 
	\_zy_simnet_tvar_53[0][22] , \_zy_simnet_tvar_53[0][21] , 
	\_zy_simnet_tvar_53[0][20] , \_zy_simnet_tvar_53[0][19] , 
	\_zy_simnet_tvar_53[0][18] , \_zy_simnet_tvar_53[0][17] , 
	\_zy_simnet_tvar_53[0][16] , \_zy_simnet_tvar_53[0][15] , 
	\_zy_simnet_tvar_53[0][14] , \_zy_simnet_tvar_53[0][13] , 
	\_zy_simnet_tvar_53[0][12] , \_zy_simnet_tvar_53[0][11] , 
	\_zy_simnet_tvar_53[0][10] , \_zy_simnet_tvar_53[0][9] , 
	\_zy_simnet_tvar_53[0][8] , \_zy_simnet_tvar_53[0][7] , 
	\_zy_simnet_tvar_53[0][6] , \_zy_simnet_tvar_53[0][5] , 
	\_zy_simnet_tvar_53[0][4] , \_zy_simnet_tvar_53[0][3] , 
	\_zy_simnet_tvar_53[0][2] , \_zy_simnet_tvar_53[0][1] , 
	\_zy_simnet_tvar_53[0][0] }), .seed0_valid( seed0_valid), 
	.seed0_internal_state_key( seed0_internal_state_key[255:0]), 
	.seed0_internal_state_value( seed0_internal_state_value[127:0]), 
	.seed0_reseed_interval( seed0_reseed_interval[47:0]), 
	.seed1_valid( seed1_valid), .seed1_internal_state_key( 
	seed1_internal_state_key[255:0]), .seed1_internal_state_value( 
	seed1_internal_state_value[127:0]), .seed1_reseed_interval( 
	seed1_reseed_interval[47:0]), .tready_override( 
	_zy_simnet_tready_override_54_w$[0:8]), 
	.cceip_encrypt_kop_fifo_override( 
	_zy_simnet_cceip_encrypt_kop_fifo_override_55_w$[0:6]), 
	.cceip_validate_kop_fifo_override( 
	_zy_simnet_cceip_validate_kop_fifo_override_56_w$[0:6]), 
	.cddip_decrypt_kop_fifo_override( 
	_zy_simnet_cddip_decrypt_kop_fifo_override_57_w$[0:6]), .manual_txc( 
	manual_txc), .always_validate_kim_ref( always_validate_kim_ref), 
	.kdf_test_mode_en( kdf_test_mode_en), .kdf_test_key_size( 
	kdf_test_key_size[31:0]), .sa_global_ctrl( 
	_zy_simnet_sa_global_ctrl_58_w$[0:31]), .sa_ctrl( { \sa_ctrl[31][31] , 
	\sa_ctrl[31][30] , \sa_ctrl[31][29] , \sa_ctrl[31][28] , 
	\sa_ctrl[31][27] , \sa_ctrl[31][26] , \sa_ctrl[31][25] , 
	\sa_ctrl[31][24] , \sa_ctrl[31][23] , \sa_ctrl[31][22] , 
	\sa_ctrl[31][21] , \sa_ctrl[31][20] , \sa_ctrl[31][19] , 
	\sa_ctrl[31][18] , \sa_ctrl[31][17] , \sa_ctrl[31][16] , 
	\sa_ctrl[31][15] , \sa_ctrl[31][14] , \sa_ctrl[31][13] , 
	\sa_ctrl[31][12] , \sa_ctrl[31][11] , \sa_ctrl[31][10] , 
	\sa_ctrl[31][9] , \sa_ctrl[31][8] , \sa_ctrl[31][7] , 
	\sa_ctrl[31][6] , \sa_ctrl[31][5] , \sa_ctrl[31][4] , 
	\sa_ctrl[31][3] , \sa_ctrl[31][2] , \sa_ctrl[31][1] , 
	\sa_ctrl[31][0] , \sa_ctrl[30][31] , \sa_ctrl[30][30] , 
	\sa_ctrl[30][29] , \sa_ctrl[30][28] , \sa_ctrl[30][27] , 
	\sa_ctrl[30][26] , \sa_ctrl[30][25] , \sa_ctrl[30][24] , 
	\sa_ctrl[30][23] , \sa_ctrl[30][22] , \sa_ctrl[30][21] , 
	\sa_ctrl[30][20] , \sa_ctrl[30][19] , \sa_ctrl[30][18] , 
	\sa_ctrl[30][17] , \sa_ctrl[30][16] , \sa_ctrl[30][15] , 
	\sa_ctrl[30][14] , \sa_ctrl[30][13] , \sa_ctrl[30][12] , 
	\sa_ctrl[30][11] , \sa_ctrl[30][10] , \sa_ctrl[30][9] , 
	\sa_ctrl[30][8] , \sa_ctrl[30][7] , \sa_ctrl[30][6] , 
	\sa_ctrl[30][5] , \sa_ctrl[30][4] , \sa_ctrl[30][3] , 
	\sa_ctrl[30][2] , \sa_ctrl[30][1] , \sa_ctrl[30][0] , 
	\sa_ctrl[29][31] , \sa_ctrl[29][30] , \sa_ctrl[29][29] , 
	\sa_ctrl[29][28] , \sa_ctrl[29][27] , \sa_ctrl[29][26] , 
	\sa_ctrl[29][25] , \sa_ctrl[29][24] , \sa_ctrl[29][23] , 
	\sa_ctrl[29][22] , \sa_ctrl[29][21] , \sa_ctrl[29][20] , 
	\sa_ctrl[29][19] , \sa_ctrl[29][18] , \sa_ctrl[29][17] , 
	\sa_ctrl[29][16] , \sa_ctrl[29][15] , \sa_ctrl[29][14] , 
	\sa_ctrl[29][13] , \sa_ctrl[29][12] , \sa_ctrl[29][11] , 
	\sa_ctrl[29][10] , \sa_ctrl[29][9] , \sa_ctrl[29][8] , 
	\sa_ctrl[29][7] , \sa_ctrl[29][6] , \sa_ctrl[29][5] , 
	\sa_ctrl[29][4] , \sa_ctrl[29][3] , \sa_ctrl[29][2] , 
	\sa_ctrl[29][1] , \sa_ctrl[29][0] , \sa_ctrl[28][31] , 
	\sa_ctrl[28][30] , \sa_ctrl[28][29] , \sa_ctrl[28][28] , 
	\sa_ctrl[28][27] , \sa_ctrl[28][26] , \sa_ctrl[28][25] , 
	\sa_ctrl[28][24] , \sa_ctrl[28][23] , \sa_ctrl[28][22] , 
	\sa_ctrl[28][21] , \sa_ctrl[28][20] , \sa_ctrl[28][19] , 
	\sa_ctrl[28][18] , \sa_ctrl[28][17] , \sa_ctrl[28][16] , 
	\sa_ctrl[28][15] , \sa_ctrl[28][14] , \sa_ctrl[28][13] , 
	\sa_ctrl[28][12] , \sa_ctrl[28][11] , \sa_ctrl[28][10] , 
	\sa_ctrl[28][9] , \sa_ctrl[28][8] , \sa_ctrl[28][7] , 
	\sa_ctrl[28][6] , \sa_ctrl[28][5] , \sa_ctrl[28][4] , 
	\sa_ctrl[28][3] , \sa_ctrl[28][2] , \sa_ctrl[28][1] , 
	\sa_ctrl[28][0] , \sa_ctrl[27][31] , \sa_ctrl[27][30] , 
	\sa_ctrl[27][29] , \sa_ctrl[27][28] , \sa_ctrl[27][27] , 
	\sa_ctrl[27][26] , \sa_ctrl[27][25] , \sa_ctrl[27][24] , 
	\sa_ctrl[27][23] , \sa_ctrl[27][22] , \sa_ctrl[27][21] , 
	\sa_ctrl[27][20] , \sa_ctrl[27][19] , \sa_ctrl[27][18] , 
	\sa_ctrl[27][17] , \sa_ctrl[27][16] , \sa_ctrl[27][15] , 
	\sa_ctrl[27][14] , \sa_ctrl[27][13] , \sa_ctrl[27][12] , 
	\sa_ctrl[27][11] , \sa_ctrl[27][10] , \sa_ctrl[27][9] , 
	\sa_ctrl[27][8] , \sa_ctrl[27][7] , \sa_ctrl[27][6] , 
	\sa_ctrl[27][5] , \sa_ctrl[27][4] , \sa_ctrl[27][3] , 
	\sa_ctrl[27][2] , \sa_ctrl[27][1] , \sa_ctrl[27][0] , 
	\sa_ctrl[26][31] , \sa_ctrl[26][30] , \sa_ctrl[26][29] , 
	\sa_ctrl[26][28] , \sa_ctrl[26][27] , \sa_ctrl[26][26] , 
	\sa_ctrl[26][25] , \sa_ctrl[26][24] , \sa_ctrl[26][23] , 
	\sa_ctrl[26][22] , \sa_ctrl[26][21] , \sa_ctrl[26][20] , 
	\sa_ctrl[26][19] , \sa_ctrl[26][18] , \sa_ctrl[26][17] , 
	\sa_ctrl[26][16] , \sa_ctrl[26][15] , \sa_ctrl[26][14] , 
	\sa_ctrl[26][13] , \sa_ctrl[26][12] , \sa_ctrl[26][11] , 
	\sa_ctrl[26][10] , \sa_ctrl[26][9] , \sa_ctrl[26][8] , 
	\sa_ctrl[26][7] , \sa_ctrl[26][6] , \sa_ctrl[26][5] , 
	\sa_ctrl[26][4] , \sa_ctrl[26][3] , \sa_ctrl[26][2] , 
	\sa_ctrl[26][1] , \sa_ctrl[26][0] , \sa_ctrl[25][31] , 
	\sa_ctrl[25][30] , \sa_ctrl[25][29] , \sa_ctrl[25][28] , 
	\sa_ctrl[25][27] , \sa_ctrl[25][26] , \sa_ctrl[25][25] , 
	\sa_ctrl[25][24] , \sa_ctrl[25][23] , \sa_ctrl[25][22] , 
	\sa_ctrl[25][21] , \sa_ctrl[25][20] , \sa_ctrl[25][19] , 
	\sa_ctrl[25][18] , \sa_ctrl[25][17] , \sa_ctrl[25][16] , 
	\sa_ctrl[25][15] , \sa_ctrl[25][14] , \sa_ctrl[25][13] , 
	\sa_ctrl[25][12] , \sa_ctrl[25][11] , \sa_ctrl[25][10] , 
	\sa_ctrl[25][9] , \sa_ctrl[25][8] , \sa_ctrl[25][7] , 
	\sa_ctrl[25][6] , \sa_ctrl[25][5] , \sa_ctrl[25][4] , 
	\sa_ctrl[25][3] , \sa_ctrl[25][2] , \sa_ctrl[25][1] , 
	\sa_ctrl[25][0] , \sa_ctrl[24][31] , \sa_ctrl[24][30] , 
	\sa_ctrl[24][29] , \sa_ctrl[24][28] , \sa_ctrl[24][27] , 
	\sa_ctrl[24][26] , \sa_ctrl[24][25] , \sa_ctrl[24][24] , 
	\sa_ctrl[24][23] , \sa_ctrl[24][22] , \sa_ctrl[24][21] , 
	\sa_ctrl[24][20] , \sa_ctrl[24][19] , \sa_ctrl[24][18] , 
	\sa_ctrl[24][17] , \sa_ctrl[24][16] , \sa_ctrl[24][15] , 
	\sa_ctrl[24][14] , \sa_ctrl[24][13] , \sa_ctrl[24][12] , 
	\sa_ctrl[24][11] , \sa_ctrl[24][10] , \sa_ctrl[24][9] , 
	\sa_ctrl[24][8] , \sa_ctrl[24][7] , \sa_ctrl[24][6] , 
	\sa_ctrl[24][5] , \sa_ctrl[24][4] , \sa_ctrl[24][3] , 
	\sa_ctrl[24][2] , \sa_ctrl[24][1] , \sa_ctrl[24][0] , 
	\sa_ctrl[23][31] , \sa_ctrl[23][30] , \sa_ctrl[23][29] , 
	\sa_ctrl[23][28] , \sa_ctrl[23][27] , \sa_ctrl[23][26] , 
	\sa_ctrl[23][25] , \sa_ctrl[23][24] , \sa_ctrl[23][23] , 
	\sa_ctrl[23][22] , \sa_ctrl[23][21] , \sa_ctrl[23][20] , 
	\sa_ctrl[23][19] , \sa_ctrl[23][18] , \sa_ctrl[23][17] , 
	\sa_ctrl[23][16] , \sa_ctrl[23][15] , \sa_ctrl[23][14] , 
	\sa_ctrl[23][13] , \sa_ctrl[23][12] , \sa_ctrl[23][11] , 
	\sa_ctrl[23][10] , \sa_ctrl[23][9] , \sa_ctrl[23][8] , 
	\sa_ctrl[23][7] , \sa_ctrl[23][6] , \sa_ctrl[23][5] , 
	\sa_ctrl[23][4] , \sa_ctrl[23][3] , \sa_ctrl[23][2] , 
	\sa_ctrl[23][1] , \sa_ctrl[23][0] , \sa_ctrl[22][31] , 
	\sa_ctrl[22][30] , \sa_ctrl[22][29] , \sa_ctrl[22][28] , 
	\sa_ctrl[22][27] , \sa_ctrl[22][26] , \sa_ctrl[22][25] , 
	\sa_ctrl[22][24] , \sa_ctrl[22][23] , \sa_ctrl[22][22] , 
	\sa_ctrl[22][21] , \sa_ctrl[22][20] , \sa_ctrl[22][19] , 
	\sa_ctrl[22][18] , \sa_ctrl[22][17] , \sa_ctrl[22][16] , 
	\sa_ctrl[22][15] , \sa_ctrl[22][14] , \sa_ctrl[22][13] , 
	\sa_ctrl[22][12] , \sa_ctrl[22][11] , \sa_ctrl[22][10] , 
	\sa_ctrl[22][9] , \sa_ctrl[22][8] , \sa_ctrl[22][7] , 
	\sa_ctrl[22][6] , \sa_ctrl[22][5] , \sa_ctrl[22][4] , 
	\sa_ctrl[22][3] , \sa_ctrl[22][2] , \sa_ctrl[22][1] , 
	\sa_ctrl[22][0] , \sa_ctrl[21][31] , \sa_ctrl[21][30] , 
	\sa_ctrl[21][29] , \sa_ctrl[21][28] , \sa_ctrl[21][27] , 
	\sa_ctrl[21][26] , \sa_ctrl[21][25] , \sa_ctrl[21][24] , 
	\sa_ctrl[21][23] , \sa_ctrl[21][22] , \sa_ctrl[21][21] , 
	\sa_ctrl[21][20] , \sa_ctrl[21][19] , \sa_ctrl[21][18] , 
	\sa_ctrl[21][17] , \sa_ctrl[21][16] , \sa_ctrl[21][15] , 
	\sa_ctrl[21][14] , \sa_ctrl[21][13] , \sa_ctrl[21][12] , 
	\sa_ctrl[21][11] , \sa_ctrl[21][10] , \sa_ctrl[21][9] , 
	\sa_ctrl[21][8] , \sa_ctrl[21][7] , \sa_ctrl[21][6] , 
	\sa_ctrl[21][5] , \sa_ctrl[21][4] , \sa_ctrl[21][3] , 
	\sa_ctrl[21][2] , \sa_ctrl[21][1] , \sa_ctrl[21][0] , 
	\sa_ctrl[20][31] , \sa_ctrl[20][30] , \sa_ctrl[20][29] , 
	\sa_ctrl[20][28] , \sa_ctrl[20][27] , \sa_ctrl[20][26] , 
	\sa_ctrl[20][25] , \sa_ctrl[20][24] , \sa_ctrl[20][23] , 
	\sa_ctrl[20][22] , \sa_ctrl[20][21] , \sa_ctrl[20][20] , 
	\sa_ctrl[20][19] , \sa_ctrl[20][18] , \sa_ctrl[20][17] , 
	\sa_ctrl[20][16] , \sa_ctrl[20][15] , \sa_ctrl[20][14] , 
	\sa_ctrl[20][13] , \sa_ctrl[20][12] , \sa_ctrl[20][11] , 
	\sa_ctrl[20][10] , \sa_ctrl[20][9] , \sa_ctrl[20][8] , 
	\sa_ctrl[20][7] , \sa_ctrl[20][6] , \sa_ctrl[20][5] , 
	\sa_ctrl[20][4] , \sa_ctrl[20][3] , \sa_ctrl[20][2] , 
	\sa_ctrl[20][1] , \sa_ctrl[20][0] , \sa_ctrl[19][31] , 
	\sa_ctrl[19][30] , \sa_ctrl[19][29] , \sa_ctrl[19][28] , 
	\sa_ctrl[19][27] , \sa_ctrl[19][26] , \sa_ctrl[19][25] , 
	\sa_ctrl[19][24] , \sa_ctrl[19][23] , \sa_ctrl[19][22] , 
	\sa_ctrl[19][21] , \sa_ctrl[19][20] , \sa_ctrl[19][19] , 
	\sa_ctrl[19][18] , \sa_ctrl[19][17] , \sa_ctrl[19][16] , 
	\sa_ctrl[19][15] , \sa_ctrl[19][14] , \sa_ctrl[19][13] , 
	\sa_ctrl[19][12] , \sa_ctrl[19][11] , \sa_ctrl[19][10] , 
	\sa_ctrl[19][9] , \sa_ctrl[19][8] , \sa_ctrl[19][7] , 
	\sa_ctrl[19][6] , \sa_ctrl[19][5] , \sa_ctrl[19][4] , 
	\sa_ctrl[19][3] , \sa_ctrl[19][2] , \sa_ctrl[19][1] , 
	\sa_ctrl[19][0] , \sa_ctrl[18][31] , \sa_ctrl[18][30] , 
	\sa_ctrl[18][29] , \sa_ctrl[18][28] , \sa_ctrl[18][27] , 
	\sa_ctrl[18][26] , \sa_ctrl[18][25] , \sa_ctrl[18][24] , 
	\sa_ctrl[18][23] , \sa_ctrl[18][22] , \sa_ctrl[18][21] , 
	\sa_ctrl[18][20] , \sa_ctrl[18][19] , \sa_ctrl[18][18] , 
	\sa_ctrl[18][17] , \sa_ctrl[18][16] , \sa_ctrl[18][15] , 
	\sa_ctrl[18][14] , \sa_ctrl[18][13] , \sa_ctrl[18][12] , 
	\sa_ctrl[18][11] , \sa_ctrl[18][10] , \sa_ctrl[18][9] , 
	\sa_ctrl[18][8] , \sa_ctrl[18][7] , \sa_ctrl[18][6] , 
	\sa_ctrl[18][5] , \sa_ctrl[18][4] , \sa_ctrl[18][3] , 
	\sa_ctrl[18][2] , \sa_ctrl[18][1] , \sa_ctrl[18][0] , 
	\sa_ctrl[17][31] , \sa_ctrl[17][30] , \sa_ctrl[17][29] , 
	\sa_ctrl[17][28] , \sa_ctrl[17][27] , \sa_ctrl[17][26] , 
	\sa_ctrl[17][25] , \sa_ctrl[17][24] , \sa_ctrl[17][23] , 
	\sa_ctrl[17][22] , \sa_ctrl[17][21] , \sa_ctrl[17][20] , 
	\sa_ctrl[17][19] , \sa_ctrl[17][18] , \sa_ctrl[17][17] , 
	\sa_ctrl[17][16] , \sa_ctrl[17][15] , \sa_ctrl[17][14] , 
	\sa_ctrl[17][13] , \sa_ctrl[17][12] , \sa_ctrl[17][11] , 
	\sa_ctrl[17][10] , \sa_ctrl[17][9] , \sa_ctrl[17][8] , 
	\sa_ctrl[17][7] , \sa_ctrl[17][6] , \sa_ctrl[17][5] , 
	\sa_ctrl[17][4] , \sa_ctrl[17][3] , \sa_ctrl[17][2] , 
	\sa_ctrl[17][1] , \sa_ctrl[17][0] , \sa_ctrl[16][31] , 
	\sa_ctrl[16][30] , \sa_ctrl[16][29] , \sa_ctrl[16][28] , 
	\sa_ctrl[16][27] , \sa_ctrl[16][26] , \sa_ctrl[16][25] , 
	\sa_ctrl[16][24] , \sa_ctrl[16][23] , \sa_ctrl[16][22] , 
	\sa_ctrl[16][21] , \sa_ctrl[16][20] , \sa_ctrl[16][19] , 
	\sa_ctrl[16][18] , \sa_ctrl[16][17] , \sa_ctrl[16][16] , 
	\sa_ctrl[16][15] , \sa_ctrl[16][14] , \sa_ctrl[16][13] , 
	\sa_ctrl[16][12] , \sa_ctrl[16][11] , \sa_ctrl[16][10] , 
	\sa_ctrl[16][9] , \sa_ctrl[16][8] , \sa_ctrl[16][7] , 
	\sa_ctrl[16][6] , \sa_ctrl[16][5] , \sa_ctrl[16][4] , 
	\sa_ctrl[16][3] , \sa_ctrl[16][2] , \sa_ctrl[16][1] , 
	\sa_ctrl[16][0] , \sa_ctrl[15][31] , \sa_ctrl[15][30] , 
	\sa_ctrl[15][29] , \sa_ctrl[15][28] , \sa_ctrl[15][27] , 
	\sa_ctrl[15][26] , \sa_ctrl[15][25] , \sa_ctrl[15][24] , 
	\sa_ctrl[15][23] , \sa_ctrl[15][22] , \sa_ctrl[15][21] , 
	\sa_ctrl[15][20] , \sa_ctrl[15][19] , \sa_ctrl[15][18] , 
	\sa_ctrl[15][17] , \sa_ctrl[15][16] , \sa_ctrl[15][15] , 
	\sa_ctrl[15][14] , \sa_ctrl[15][13] , \sa_ctrl[15][12] , 
	\sa_ctrl[15][11] , \sa_ctrl[15][10] , \sa_ctrl[15][9] , 
	\sa_ctrl[15][8] , \sa_ctrl[15][7] , \sa_ctrl[15][6] , 
	\sa_ctrl[15][5] , \sa_ctrl[15][4] , \sa_ctrl[15][3] , 
	\sa_ctrl[15][2] , \sa_ctrl[15][1] , \sa_ctrl[15][0] , 
	\sa_ctrl[14][31] , \sa_ctrl[14][30] , \sa_ctrl[14][29] , 
	\sa_ctrl[14][28] , \sa_ctrl[14][27] , \sa_ctrl[14][26] , 
	\sa_ctrl[14][25] , \sa_ctrl[14][24] , \sa_ctrl[14][23] , 
	\sa_ctrl[14][22] , \sa_ctrl[14][21] , \sa_ctrl[14][20] , 
	\sa_ctrl[14][19] , \sa_ctrl[14][18] , \sa_ctrl[14][17] , 
	\sa_ctrl[14][16] , \sa_ctrl[14][15] , \sa_ctrl[14][14] , 
	\sa_ctrl[14][13] , \sa_ctrl[14][12] , \sa_ctrl[14][11] , 
	\sa_ctrl[14][10] , \sa_ctrl[14][9] , \sa_ctrl[14][8] , 
	\sa_ctrl[14][7] , \sa_ctrl[14][6] , \sa_ctrl[14][5] , 
	\sa_ctrl[14][4] , \sa_ctrl[14][3] , \sa_ctrl[14][2] , 
	\sa_ctrl[14][1] , \sa_ctrl[14][0] , \sa_ctrl[13][31] , 
	\sa_ctrl[13][30] , \sa_ctrl[13][29] , \sa_ctrl[13][28] , 
	\sa_ctrl[13][27] , \sa_ctrl[13][26] , \sa_ctrl[13][25] , 
	\sa_ctrl[13][24] , \sa_ctrl[13][23] , \sa_ctrl[13][22] , 
	\sa_ctrl[13][21] , \sa_ctrl[13][20] , \sa_ctrl[13][19] , 
	\sa_ctrl[13][18] , \sa_ctrl[13][17] , \sa_ctrl[13][16] , 
	\sa_ctrl[13][15] , \sa_ctrl[13][14] , \sa_ctrl[13][13] , 
	\sa_ctrl[13][12] , \sa_ctrl[13][11] , \sa_ctrl[13][10] , 
	\sa_ctrl[13][9] , \sa_ctrl[13][8] , \sa_ctrl[13][7] , 
	\sa_ctrl[13][6] , \sa_ctrl[13][5] , \sa_ctrl[13][4] , 
	\sa_ctrl[13][3] , \sa_ctrl[13][2] , \sa_ctrl[13][1] , 
	\sa_ctrl[13][0] , \sa_ctrl[12][31] , \sa_ctrl[12][30] , 
	\sa_ctrl[12][29] , \sa_ctrl[12][28] , \sa_ctrl[12][27] , 
	\sa_ctrl[12][26] , \sa_ctrl[12][25] , \sa_ctrl[12][24] , 
	\sa_ctrl[12][23] , \sa_ctrl[12][22] , \sa_ctrl[12][21] , 
	\sa_ctrl[12][20] , \sa_ctrl[12][19] , \sa_ctrl[12][18] , 
	\sa_ctrl[12][17] , \sa_ctrl[12][16] , \sa_ctrl[12][15] , 
	\sa_ctrl[12][14] , \sa_ctrl[12][13] , \sa_ctrl[12][12] , 
	\sa_ctrl[12][11] , \sa_ctrl[12][10] , \sa_ctrl[12][9] , 
	\sa_ctrl[12][8] , \sa_ctrl[12][7] , \sa_ctrl[12][6] , 
	\sa_ctrl[12][5] , \sa_ctrl[12][4] , \sa_ctrl[12][3] , 
	\sa_ctrl[12][2] , \sa_ctrl[12][1] , \sa_ctrl[12][0] , 
	\sa_ctrl[11][31] , \sa_ctrl[11][30] , \sa_ctrl[11][29] , 
	\sa_ctrl[11][28] , \sa_ctrl[11][27] , \sa_ctrl[11][26] , 
	\sa_ctrl[11][25] , \sa_ctrl[11][24] , \sa_ctrl[11][23] , 
	\sa_ctrl[11][22] , \sa_ctrl[11][21] , \sa_ctrl[11][20] , 
	\sa_ctrl[11][19] , \sa_ctrl[11][18] , \sa_ctrl[11][17] , 
	\sa_ctrl[11][16] , \sa_ctrl[11][15] , \sa_ctrl[11][14] , 
	\sa_ctrl[11][13] , \sa_ctrl[11][12] , \sa_ctrl[11][11] , 
	\sa_ctrl[11][10] , \sa_ctrl[11][9] , \sa_ctrl[11][8] , 
	\sa_ctrl[11][7] , \sa_ctrl[11][6] , \sa_ctrl[11][5] , 
	\sa_ctrl[11][4] , \sa_ctrl[11][3] , \sa_ctrl[11][2] , 
	\sa_ctrl[11][1] , \sa_ctrl[11][0] , \sa_ctrl[10][31] , 
	\sa_ctrl[10][30] , \sa_ctrl[10][29] , \sa_ctrl[10][28] , 
	\sa_ctrl[10][27] , \sa_ctrl[10][26] , \sa_ctrl[10][25] , 
	\sa_ctrl[10][24] , \sa_ctrl[10][23] , \sa_ctrl[10][22] , 
	\sa_ctrl[10][21] , \sa_ctrl[10][20] , \sa_ctrl[10][19] , 
	\sa_ctrl[10][18] , \sa_ctrl[10][17] , \sa_ctrl[10][16] , 
	\sa_ctrl[10][15] , \sa_ctrl[10][14] , \sa_ctrl[10][13] , 
	\sa_ctrl[10][12] , \sa_ctrl[10][11] , \sa_ctrl[10][10] , 
	\sa_ctrl[10][9] , \sa_ctrl[10][8] , \sa_ctrl[10][7] , 
	\sa_ctrl[10][6] , \sa_ctrl[10][5] , \sa_ctrl[10][4] , 
	\sa_ctrl[10][3] , \sa_ctrl[10][2] , \sa_ctrl[10][1] , 
	\sa_ctrl[10][0] , \sa_ctrl[9][31] , \sa_ctrl[9][30] , 
	\sa_ctrl[9][29] , \sa_ctrl[9][28] , \sa_ctrl[9][27] , 
	\sa_ctrl[9][26] , \sa_ctrl[9][25] , \sa_ctrl[9][24] , 
	\sa_ctrl[9][23] , \sa_ctrl[9][22] , \sa_ctrl[9][21] , 
	\sa_ctrl[9][20] , \sa_ctrl[9][19] , \sa_ctrl[9][18] , 
	\sa_ctrl[9][17] , \sa_ctrl[9][16] , \sa_ctrl[9][15] , 
	\sa_ctrl[9][14] , \sa_ctrl[9][13] , \sa_ctrl[9][12] , 
	\sa_ctrl[9][11] , \sa_ctrl[9][10] , \sa_ctrl[9][9] , \sa_ctrl[9][8] , 
	\sa_ctrl[9][7] , \sa_ctrl[9][6] , \sa_ctrl[9][5] , \sa_ctrl[9][4] , 
	\sa_ctrl[9][3] , \sa_ctrl[9][2] , \sa_ctrl[9][1] , \sa_ctrl[9][0] , 
	\sa_ctrl[8][31] , \sa_ctrl[8][30] , \sa_ctrl[8][29] , 
	\sa_ctrl[8][28] , \sa_ctrl[8][27] , \sa_ctrl[8][26] , 
	\sa_ctrl[8][25] , \sa_ctrl[8][24] , \sa_ctrl[8][23] , 
	\sa_ctrl[8][22] , \sa_ctrl[8][21] , \sa_ctrl[8][20] , 
	\sa_ctrl[8][19] , \sa_ctrl[8][18] , \sa_ctrl[8][17] , 
	\sa_ctrl[8][16] , \sa_ctrl[8][15] , \sa_ctrl[8][14] , 
	\sa_ctrl[8][13] , \sa_ctrl[8][12] , \sa_ctrl[8][11] , 
	\sa_ctrl[8][10] , \sa_ctrl[8][9] , \sa_ctrl[8][8] , \sa_ctrl[8][7] , 
	\sa_ctrl[8][6] , \sa_ctrl[8][5] , \sa_ctrl[8][4] , \sa_ctrl[8][3] , 
	\sa_ctrl[8][2] , \sa_ctrl[8][1] , \sa_ctrl[8][0] , \sa_ctrl[7][31] , 
	\sa_ctrl[7][30] , \sa_ctrl[7][29] , \sa_ctrl[7][28] , 
	\sa_ctrl[7][27] , \sa_ctrl[7][26] , \sa_ctrl[7][25] , 
	\sa_ctrl[7][24] , \sa_ctrl[7][23] , \sa_ctrl[7][22] , 
	\sa_ctrl[7][21] , \sa_ctrl[7][20] , \sa_ctrl[7][19] , 
	\sa_ctrl[7][18] , \sa_ctrl[7][17] , \sa_ctrl[7][16] , 
	\sa_ctrl[7][15] , \sa_ctrl[7][14] , \sa_ctrl[7][13] , 
	\sa_ctrl[7][12] , \sa_ctrl[7][11] , \sa_ctrl[7][10] , 
	\sa_ctrl[7][9] , \sa_ctrl[7][8] , \sa_ctrl[7][7] , \sa_ctrl[7][6] , 
	\sa_ctrl[7][5] , \sa_ctrl[7][4] , \sa_ctrl[7][3] , \sa_ctrl[7][2] , 
	\sa_ctrl[7][1] , \sa_ctrl[7][0] , \sa_ctrl[6][31] , \sa_ctrl[6][30] , 
	\sa_ctrl[6][29] , \sa_ctrl[6][28] , \sa_ctrl[6][27] , 
	\sa_ctrl[6][26] , \sa_ctrl[6][25] , \sa_ctrl[6][24] , 
	\sa_ctrl[6][23] , \sa_ctrl[6][22] , \sa_ctrl[6][21] , 
	\sa_ctrl[6][20] , \sa_ctrl[6][19] , \sa_ctrl[6][18] , 
	\sa_ctrl[6][17] , \sa_ctrl[6][16] , \sa_ctrl[6][15] , 
	\sa_ctrl[6][14] , \sa_ctrl[6][13] , \sa_ctrl[6][12] , 
	\sa_ctrl[6][11] , \sa_ctrl[6][10] , \sa_ctrl[6][9] , \sa_ctrl[6][8] , 
	\sa_ctrl[6][7] , \sa_ctrl[6][6] , \sa_ctrl[6][5] , \sa_ctrl[6][4] , 
	\sa_ctrl[6][3] , \sa_ctrl[6][2] , \sa_ctrl[6][1] , \sa_ctrl[6][0] , 
	\sa_ctrl[5][31] , \sa_ctrl[5][30] , \sa_ctrl[5][29] , 
	\sa_ctrl[5][28] , \sa_ctrl[5][27] , \sa_ctrl[5][26] , 
	\sa_ctrl[5][25] , \sa_ctrl[5][24] , \sa_ctrl[5][23] , 
	\sa_ctrl[5][22] , \sa_ctrl[5][21] , \sa_ctrl[5][20] , 
	\sa_ctrl[5][19] , \sa_ctrl[5][18] , \sa_ctrl[5][17] , 
	\sa_ctrl[5][16] , \sa_ctrl[5][15] , \sa_ctrl[5][14] , 
	\sa_ctrl[5][13] , \sa_ctrl[5][12] , \sa_ctrl[5][11] , 
	\sa_ctrl[5][10] , \sa_ctrl[5][9] , \sa_ctrl[5][8] , \sa_ctrl[5][7] , 
	\sa_ctrl[5][6] , \sa_ctrl[5][5] , \sa_ctrl[5][4] , \sa_ctrl[5][3] , 
	\sa_ctrl[5][2] , \sa_ctrl[5][1] , \sa_ctrl[5][0] , \sa_ctrl[4][31] , 
	\sa_ctrl[4][30] , \sa_ctrl[4][29] , \sa_ctrl[4][28] , 
	\sa_ctrl[4][27] , \sa_ctrl[4][26] , \sa_ctrl[4][25] , 
	\sa_ctrl[4][24] , \sa_ctrl[4][23] , \sa_ctrl[4][22] , 
	\sa_ctrl[4][21] , \sa_ctrl[4][20] , \sa_ctrl[4][19] , 
	\sa_ctrl[4][18] , \sa_ctrl[4][17] , \sa_ctrl[4][16] , 
	\sa_ctrl[4][15] , \sa_ctrl[4][14] , \sa_ctrl[4][13] , 
	\sa_ctrl[4][12] , \sa_ctrl[4][11] , \sa_ctrl[4][10] , 
	\sa_ctrl[4][9] , \sa_ctrl[4][8] , \sa_ctrl[4][7] , \sa_ctrl[4][6] , 
	\sa_ctrl[4][5] , \sa_ctrl[4][4] , \sa_ctrl[4][3] , \sa_ctrl[4][2] , 
	\sa_ctrl[4][1] , \sa_ctrl[4][0] , \sa_ctrl[3][31] , \sa_ctrl[3][30] , 
	\sa_ctrl[3][29] , \sa_ctrl[3][28] , \sa_ctrl[3][27] , 
	\sa_ctrl[3][26] , \sa_ctrl[3][25] , \sa_ctrl[3][24] , 
	\sa_ctrl[3][23] , \sa_ctrl[3][22] , \sa_ctrl[3][21] , 
	\sa_ctrl[3][20] , \sa_ctrl[3][19] , \sa_ctrl[3][18] , 
	\sa_ctrl[3][17] , \sa_ctrl[3][16] , \sa_ctrl[3][15] , 
	\sa_ctrl[3][14] , \sa_ctrl[3][13] , \sa_ctrl[3][12] , 
	\sa_ctrl[3][11] , \sa_ctrl[3][10] , \sa_ctrl[3][9] , \sa_ctrl[3][8] , 
	\sa_ctrl[3][7] , \sa_ctrl[3][6] , \sa_ctrl[3][5] , \sa_ctrl[3][4] , 
	\sa_ctrl[3][3] , \sa_ctrl[3][2] , \sa_ctrl[3][1] , \sa_ctrl[3][0] , 
	\sa_ctrl[2][31] , \sa_ctrl[2][30] , \sa_ctrl[2][29] , 
	\sa_ctrl[2][28] , \sa_ctrl[2][27] , \sa_ctrl[2][26] , 
	\sa_ctrl[2][25] , \sa_ctrl[2][24] , \sa_ctrl[2][23] , 
	\sa_ctrl[2][22] , \sa_ctrl[2][21] , \sa_ctrl[2][20] , 
	\sa_ctrl[2][19] , \sa_ctrl[2][18] , \sa_ctrl[2][17] , 
	\sa_ctrl[2][16] , \sa_ctrl[2][15] , \sa_ctrl[2][14] , 
	\sa_ctrl[2][13] , \sa_ctrl[2][12] , \sa_ctrl[2][11] , 
	\sa_ctrl[2][10] , \sa_ctrl[2][9] , \sa_ctrl[2][8] , \sa_ctrl[2][7] , 
	\sa_ctrl[2][6] , \sa_ctrl[2][5] , \sa_ctrl[2][4] , \sa_ctrl[2][3] , 
	\sa_ctrl[2][2] , \sa_ctrl[2][1] , \sa_ctrl[2][0] , \sa_ctrl[1][31] , 
	\sa_ctrl[1][30] , \sa_ctrl[1][29] , \sa_ctrl[1][28] , 
	\sa_ctrl[1][27] , \sa_ctrl[1][26] , \sa_ctrl[1][25] , 
	\sa_ctrl[1][24] , \sa_ctrl[1][23] , \sa_ctrl[1][22] , 
	\sa_ctrl[1][21] , \sa_ctrl[1][20] , \sa_ctrl[1][19] , 
	\sa_ctrl[1][18] , \sa_ctrl[1][17] , \sa_ctrl[1][16] , 
	\sa_ctrl[1][15] , \sa_ctrl[1][14] , \sa_ctrl[1][13] , 
	\sa_ctrl[1][12] , \sa_ctrl[1][11] , \sa_ctrl[1][10] , 
	\sa_ctrl[1][9] , \sa_ctrl[1][8] , \sa_ctrl[1][7] , \sa_ctrl[1][6] , 
	\sa_ctrl[1][5] , \sa_ctrl[1][4] , \sa_ctrl[1][3] , \sa_ctrl[1][2] , 
	\sa_ctrl[1][1] , \sa_ctrl[1][0] , \sa_ctrl[0][31] , \sa_ctrl[0][30] , 
	\sa_ctrl[0][29] , \sa_ctrl[0][28] , \sa_ctrl[0][27] , 
	\sa_ctrl[0][26] , \sa_ctrl[0][25] , \sa_ctrl[0][24] , 
	\sa_ctrl[0][23] , \sa_ctrl[0][22] , \sa_ctrl[0][21] , 
	\sa_ctrl[0][20] , \sa_ctrl[0][19] , \sa_ctrl[0][18] , 
	\sa_ctrl[0][17] , \sa_ctrl[0][16] , \sa_ctrl[0][15] , 
	\sa_ctrl[0][14] , \sa_ctrl[0][13] , \sa_ctrl[0][12] , 
	\sa_ctrl[0][11] , \sa_ctrl[0][10] , \sa_ctrl[0][9] , \sa_ctrl[0][8] , 
	\sa_ctrl[0][7] , \sa_ctrl[0][6] , \sa_ctrl[0][5] , \sa_ctrl[0][4] , 
	\sa_ctrl[0][3] , \sa_ctrl[0][2] , \sa_ctrl[0][1] , \sa_ctrl[0][0] }), 
	.debug_kme_ib_tvalid( debug_kme_ib_tvalid), .debug_kme_ib_tlast( 
	debug_kme_ib_tlast), .debug_kme_ib_tid( debug_kme_ib_tid[0]), 
	.debug_kme_ib_tstrb( debug_kme_ib_tstrb[7:0]), .debug_kme_ib_tuser( 
	debug_kme_ib_tuser[7:0]), .debug_kme_ib_tdata( 
	debug_kme_ib_tdata[63:0]), .clk( clk), .rst_n( rst_sync_n), .ovstb( 
	ovstb), .lvm( lvm), .mlvm( mlvm), .rbus_ring_i( 
	_zy_simnet_rbus_ring_i_59_w$[0:83]), .cfg_start_addr( 
	_zy_simnet_cio_60[0:15]), .cfg_end_addr( _zy_simnet_cio_61[0:15]), 
	.kme_cceip0_ob_out_pre( _zy_simnet_kme_cceip0_ob_out_pre_62_w$[0:82]), 
	.kme_cceip0_ob_in( _zy_simnet_kme_cceip0_ob_in_63_w$), 
	.kme_cceip1_ob_out_pre( _zy_simnet_kme_cceip1_ob_out_pre_64_w$[0:82]), 
	.kme_cceip1_ob_in( _zy_simnet_kme_cceip1_ob_in_65_w$), 
	.kme_cceip2_ob_out_pre( _zy_simnet_kme_cceip2_ob_out_pre_66_w$[0:82]), 
	.kme_cceip2_ob_in( _zy_simnet_kme_cceip2_ob_in_67_w$), 
	.kme_cceip3_ob_out_pre( _zy_simnet_kme_cceip3_ob_out_pre_68_w$[0:82]), 
	.kme_cceip3_ob_in( _zy_simnet_kme_cceip3_ob_in_69_w$), 
	.kme_cddip0_ob_out_pre( _zy_simnet_kme_cddip0_ob_out_pre_70_w$[0:82]), 
	.kme_cddip0_ob_in( _zy_simnet_kme_cddip0_ob_in_71_w$), 
	.kme_cddip1_ob_out_pre( _zy_simnet_kme_cddip1_ob_out_pre_72_w$[0:82]), 
	.kme_cddip1_ob_in( _zy_simnet_kme_cddip1_ob_in_73_w$), 
	.kme_cddip2_ob_out_pre( _zy_simnet_kme_cddip2_ob_out_pre_74_w$[0:82]), 
	.kme_cddip2_ob_in( _zy_simnet_kme_cddip2_ob_in_75_w$), 
	.kme_cddip3_ob_out_pre( _zy_simnet_kme_cddip3_ob_out_pre_76_w$[0:82]), 
	.kme_cddip3_ob_in( _zy_simnet_kme_cddip3_ob_in_77_w$), .ckv_rd( 
	ckv_rd), .ckv_addr( ckv_addr[14:0]), .kim_rd( kim_rd), .kim_addr( 
	kim_addr[13:0]), .cceip_encrypt_bimc_osync( cceip_encrypt_bimc_osync), 
	.cceip_encrypt_bimc_odat( cceip_encrypt_bimc_odat), 
	.cceip_encrypt_mbe( cceip_encrypt_mbe), .cceip_validate_bimc_osync( 
	cceip_validate_bimc_osync), .cceip_validate_bimc_odat( 
	cceip_validate_bimc_odat), .cceip_validate_mbe( cceip_validate_mbe), 
	.cddip_decrypt_bimc_osync( cddip_decrypt_bimc_osync), 
	.cddip_decrypt_bimc_odat( cddip_decrypt_bimc_odat), 
	.cddip_decrypt_mbe( cddip_decrypt_mbe), .axi_bimc_osync( 
	axi_bimc_osync), .axi_bimc_odat( axi_bimc_odat), .axi_mbe( axi_mbe), 
	.seed0_invalidate( seed0_invalidate), .seed1_invalidate( 
	seed1_invalidate), .set_txc_bp_int( set_txc_bp_int), 
	.set_gcm_tag_fail_int( set_gcm_tag_fail_int), 
	.set_key_tlv_miscmp_int( set_key_tlv_miscmp_int), 
	.set_tlv_bip2_error_int( set_tlv_bip2_error_int), 
	.set_rsm_is_backpressuring( set_rsm_is_backpressuring[7:0]), 
	.idle_components( _zy_simnet_idle_components_78_w$[0:31]), 
	.sa_snapshot( { \sa_snapshot[31][63] , \sa_snapshot[31][62] , 
	\sa_snapshot[31][61] , \sa_snapshot[31][60] , \sa_snapshot[31][59] , 
	\sa_snapshot[31][58] , \sa_snapshot[31][57] , \sa_snapshot[31][56] , 
	\sa_snapshot[31][55] , \sa_snapshot[31][54] , \sa_snapshot[31][53] , 
	\sa_snapshot[31][52] , \sa_snapshot[31][51] , \sa_snapshot[31][50] , 
	\sa_snapshot[31][49] , \sa_snapshot[31][48] , \sa_snapshot[31][47] , 
	\sa_snapshot[31][46] , \sa_snapshot[31][45] , \sa_snapshot[31][44] , 
	\sa_snapshot[31][43] , \sa_snapshot[31][42] , \sa_snapshot[31][41] , 
	\sa_snapshot[31][40] , \sa_snapshot[31][39] , \sa_snapshot[31][38] , 
	\sa_snapshot[31][37] , \sa_snapshot[31][36] , \sa_snapshot[31][35] , 
	\sa_snapshot[31][34] , \sa_snapshot[31][33] , \sa_snapshot[31][32] , 
	\sa_snapshot[31][31] , \sa_snapshot[31][30] , \sa_snapshot[31][29] , 
	\sa_snapshot[31][28] , \sa_snapshot[31][27] , \sa_snapshot[31][26] , 
	\sa_snapshot[31][25] , \sa_snapshot[31][24] , \sa_snapshot[31][23] , 
	\sa_snapshot[31][22] , \sa_snapshot[31][21] , \sa_snapshot[31][20] , 
	\sa_snapshot[31][19] , \sa_snapshot[31][18] , \sa_snapshot[31][17] , 
	\sa_snapshot[31][16] , \sa_snapshot[31][15] , \sa_snapshot[31][14] , 
	\sa_snapshot[31][13] , \sa_snapshot[31][12] , \sa_snapshot[31][11] , 
	\sa_snapshot[31][10] , \sa_snapshot[31][9] , \sa_snapshot[31][8] , 
	\sa_snapshot[31][7] , \sa_snapshot[31][6] , \sa_snapshot[31][5] , 
	\sa_snapshot[31][4] , \sa_snapshot[31][3] , \sa_snapshot[31][2] , 
	\sa_snapshot[31][1] , \sa_snapshot[31][0] , \sa_snapshot[30][63] , 
	\sa_snapshot[30][62] , \sa_snapshot[30][61] , \sa_snapshot[30][60] , 
	\sa_snapshot[30][59] , \sa_snapshot[30][58] , \sa_snapshot[30][57] , 
	\sa_snapshot[30][56] , \sa_snapshot[30][55] , \sa_snapshot[30][54] , 
	\sa_snapshot[30][53] , \sa_snapshot[30][52] , \sa_snapshot[30][51] , 
	\sa_snapshot[30][50] , \sa_snapshot[30][49] , \sa_snapshot[30][48] , 
	\sa_snapshot[30][47] , \sa_snapshot[30][46] , \sa_snapshot[30][45] , 
	\sa_snapshot[30][44] , \sa_snapshot[30][43] , \sa_snapshot[30][42] , 
	\sa_snapshot[30][41] , \sa_snapshot[30][40] , \sa_snapshot[30][39] , 
	\sa_snapshot[30][38] , \sa_snapshot[30][37] , \sa_snapshot[30][36] , 
	\sa_snapshot[30][35] , \sa_snapshot[30][34] , \sa_snapshot[30][33] , 
	\sa_snapshot[30][32] , \sa_snapshot[30][31] , \sa_snapshot[30][30] , 
	\sa_snapshot[30][29] , \sa_snapshot[30][28] , \sa_snapshot[30][27] , 
	\sa_snapshot[30][26] , \sa_snapshot[30][25] , \sa_snapshot[30][24] , 
	\sa_snapshot[30][23] , \sa_snapshot[30][22] , \sa_snapshot[30][21] , 
	\sa_snapshot[30][20] , \sa_snapshot[30][19] , \sa_snapshot[30][18] , 
	\sa_snapshot[30][17] , \sa_snapshot[30][16] , \sa_snapshot[30][15] , 
	\sa_snapshot[30][14] , \sa_snapshot[30][13] , \sa_snapshot[30][12] , 
	\sa_snapshot[30][11] , \sa_snapshot[30][10] , \sa_snapshot[30][9] , 
	\sa_snapshot[30][8] , \sa_snapshot[30][7] , \sa_snapshot[30][6] , 
	\sa_snapshot[30][5] , \sa_snapshot[30][4] , \sa_snapshot[30][3] , 
	\sa_snapshot[30][2] , \sa_snapshot[30][1] , \sa_snapshot[30][0] , 
	\sa_snapshot[29][63] , \sa_snapshot[29][62] , \sa_snapshot[29][61] , 
	\sa_snapshot[29][60] , \sa_snapshot[29][59] , \sa_snapshot[29][58] , 
	\sa_snapshot[29][57] , \sa_snapshot[29][56] , \sa_snapshot[29][55] , 
	\sa_snapshot[29][54] , \sa_snapshot[29][53] , \sa_snapshot[29][52] , 
	\sa_snapshot[29][51] , \sa_snapshot[29][50] , \sa_snapshot[29][49] , 
	\sa_snapshot[29][48] , \sa_snapshot[29][47] , \sa_snapshot[29][46] , 
	\sa_snapshot[29][45] , \sa_snapshot[29][44] , \sa_snapshot[29][43] , 
	\sa_snapshot[29][42] , \sa_snapshot[29][41] , \sa_snapshot[29][40] , 
	\sa_snapshot[29][39] , \sa_snapshot[29][38] , \sa_snapshot[29][37] , 
	\sa_snapshot[29][36] , \sa_snapshot[29][35] , \sa_snapshot[29][34] , 
	\sa_snapshot[29][33] , \sa_snapshot[29][32] , \sa_snapshot[29][31] , 
	\sa_snapshot[29][30] , \sa_snapshot[29][29] , \sa_snapshot[29][28] , 
	\sa_snapshot[29][27] , \sa_snapshot[29][26] , \sa_snapshot[29][25] , 
	\sa_snapshot[29][24] , \sa_snapshot[29][23] , \sa_snapshot[29][22] , 
	\sa_snapshot[29][21] , \sa_snapshot[29][20] , \sa_snapshot[29][19] , 
	\sa_snapshot[29][18] , \sa_snapshot[29][17] , \sa_snapshot[29][16] , 
	\sa_snapshot[29][15] , \sa_snapshot[29][14] , \sa_snapshot[29][13] , 
	\sa_snapshot[29][12] , \sa_snapshot[29][11] , \sa_snapshot[29][10] , 
	\sa_snapshot[29][9] , \sa_snapshot[29][8] , \sa_snapshot[29][7] , 
	\sa_snapshot[29][6] , \sa_snapshot[29][5] , \sa_snapshot[29][4] , 
	\sa_snapshot[29][3] , \sa_snapshot[29][2] , \sa_snapshot[29][1] , 
	\sa_snapshot[29][0] , \sa_snapshot[28][63] , \sa_snapshot[28][62] , 
	\sa_snapshot[28][61] , \sa_snapshot[28][60] , \sa_snapshot[28][59] , 
	\sa_snapshot[28][58] , \sa_snapshot[28][57] , \sa_snapshot[28][56] , 
	\sa_snapshot[28][55] , \sa_snapshot[28][54] , \sa_snapshot[28][53] , 
	\sa_snapshot[28][52] , \sa_snapshot[28][51] , \sa_snapshot[28][50] , 
	\sa_snapshot[28][49] , \sa_snapshot[28][48] , \sa_snapshot[28][47] , 
	\sa_snapshot[28][46] , \sa_snapshot[28][45] , \sa_snapshot[28][44] , 
	\sa_snapshot[28][43] , \sa_snapshot[28][42] , \sa_snapshot[28][41] , 
	\sa_snapshot[28][40] , \sa_snapshot[28][39] , \sa_snapshot[28][38] , 
	\sa_snapshot[28][37] , \sa_snapshot[28][36] , \sa_snapshot[28][35] , 
	\sa_snapshot[28][34] , \sa_snapshot[28][33] , \sa_snapshot[28][32] , 
	\sa_snapshot[28][31] , \sa_snapshot[28][30] , \sa_snapshot[28][29] , 
	\sa_snapshot[28][28] , \sa_snapshot[28][27] , \sa_snapshot[28][26] , 
	\sa_snapshot[28][25] , \sa_snapshot[28][24] , \sa_snapshot[28][23] , 
	\sa_snapshot[28][22] , \sa_snapshot[28][21] , \sa_snapshot[28][20] , 
	\sa_snapshot[28][19] , \sa_snapshot[28][18] , \sa_snapshot[28][17] , 
	\sa_snapshot[28][16] , \sa_snapshot[28][15] , \sa_snapshot[28][14] , 
	\sa_snapshot[28][13] , \sa_snapshot[28][12] , \sa_snapshot[28][11] , 
	\sa_snapshot[28][10] , \sa_snapshot[28][9] , \sa_snapshot[28][8] , 
	\sa_snapshot[28][7] , \sa_snapshot[28][6] , \sa_snapshot[28][5] , 
	\sa_snapshot[28][4] , \sa_snapshot[28][3] , \sa_snapshot[28][2] , 
	\sa_snapshot[28][1] , \sa_snapshot[28][0] , \sa_snapshot[27][63] , 
	\sa_snapshot[27][62] , \sa_snapshot[27][61] , \sa_snapshot[27][60] , 
	\sa_snapshot[27][59] , \sa_snapshot[27][58] , \sa_snapshot[27][57] , 
	\sa_snapshot[27][56] , \sa_snapshot[27][55] , \sa_snapshot[27][54] , 
	\sa_snapshot[27][53] , \sa_snapshot[27][52] , \sa_snapshot[27][51] , 
	\sa_snapshot[27][50] , \sa_snapshot[27][49] , \sa_snapshot[27][48] , 
	\sa_snapshot[27][47] , \sa_snapshot[27][46] , \sa_snapshot[27][45] , 
	\sa_snapshot[27][44] , \sa_snapshot[27][43] , \sa_snapshot[27][42] , 
	\sa_snapshot[27][41] , \sa_snapshot[27][40] , \sa_snapshot[27][39] , 
	\sa_snapshot[27][38] , \sa_snapshot[27][37] , \sa_snapshot[27][36] , 
	\sa_snapshot[27][35] , \sa_snapshot[27][34] , \sa_snapshot[27][33] , 
	\sa_snapshot[27][32] , \sa_snapshot[27][31] , \sa_snapshot[27][30] , 
	\sa_snapshot[27][29] , \sa_snapshot[27][28] , \sa_snapshot[27][27] , 
	\sa_snapshot[27][26] , \sa_snapshot[27][25] , \sa_snapshot[27][24] , 
	\sa_snapshot[27][23] , \sa_snapshot[27][22] , \sa_snapshot[27][21] , 
	\sa_snapshot[27][20] , \sa_snapshot[27][19] , \sa_snapshot[27][18] , 
	\sa_snapshot[27][17] , \sa_snapshot[27][16] , \sa_snapshot[27][15] , 
	\sa_snapshot[27][14] , \sa_snapshot[27][13] , \sa_snapshot[27][12] , 
	\sa_snapshot[27][11] , \sa_snapshot[27][10] , \sa_snapshot[27][9] , 
	\sa_snapshot[27][8] , \sa_snapshot[27][7] , \sa_snapshot[27][6] , 
	\sa_snapshot[27][5] , \sa_snapshot[27][4] , \sa_snapshot[27][3] , 
	\sa_snapshot[27][2] , \sa_snapshot[27][1] , \sa_snapshot[27][0] , 
	\sa_snapshot[26][63] , \sa_snapshot[26][62] , \sa_snapshot[26][61] , 
	\sa_snapshot[26][60] , \sa_snapshot[26][59] , \sa_snapshot[26][58] , 
	\sa_snapshot[26][57] , \sa_snapshot[26][56] , \sa_snapshot[26][55] , 
	\sa_snapshot[26][54] , \sa_snapshot[26][53] , \sa_snapshot[26][52] , 
	\sa_snapshot[26][51] , \sa_snapshot[26][50] , \sa_snapshot[26][49] , 
	\sa_snapshot[26][48] , \sa_snapshot[26][47] , \sa_snapshot[26][46] , 
	\sa_snapshot[26][45] , \sa_snapshot[26][44] , \sa_snapshot[26][43] , 
	\sa_snapshot[26][42] , \sa_snapshot[26][41] , \sa_snapshot[26][40] , 
	\sa_snapshot[26][39] , \sa_snapshot[26][38] , \sa_snapshot[26][37] , 
	\sa_snapshot[26][36] , \sa_snapshot[26][35] , \sa_snapshot[26][34] , 
	\sa_snapshot[26][33] , \sa_snapshot[26][32] , \sa_snapshot[26][31] , 
	\sa_snapshot[26][30] , \sa_snapshot[26][29] , \sa_snapshot[26][28] , 
	\sa_snapshot[26][27] , \sa_snapshot[26][26] , \sa_snapshot[26][25] , 
	\sa_snapshot[26][24] , \sa_snapshot[26][23] , \sa_snapshot[26][22] , 
	\sa_snapshot[26][21] , \sa_snapshot[26][20] , \sa_snapshot[26][19] , 
	\sa_snapshot[26][18] , \sa_snapshot[26][17] , \sa_snapshot[26][16] , 
	\sa_snapshot[26][15] , \sa_snapshot[26][14] , \sa_snapshot[26][13] , 
	\sa_snapshot[26][12] , \sa_snapshot[26][11] , \sa_snapshot[26][10] , 
	\sa_snapshot[26][9] , \sa_snapshot[26][8] , \sa_snapshot[26][7] , 
	\sa_snapshot[26][6] , \sa_snapshot[26][5] , \sa_snapshot[26][4] , 
	\sa_snapshot[26][3] , \sa_snapshot[26][2] , \sa_snapshot[26][1] , 
	\sa_snapshot[26][0] , \sa_snapshot[25][63] , \sa_snapshot[25][62] , 
	\sa_snapshot[25][61] , \sa_snapshot[25][60] , \sa_snapshot[25][59] , 
	\sa_snapshot[25][58] , \sa_snapshot[25][57] , \sa_snapshot[25][56] , 
	\sa_snapshot[25][55] , \sa_snapshot[25][54] , \sa_snapshot[25][53] , 
	\sa_snapshot[25][52] , \sa_snapshot[25][51] , \sa_snapshot[25][50] , 
	\sa_snapshot[25][49] , \sa_snapshot[25][48] , \sa_snapshot[25][47] , 
	\sa_snapshot[25][46] , \sa_snapshot[25][45] , \sa_snapshot[25][44] , 
	\sa_snapshot[25][43] , \sa_snapshot[25][42] , \sa_snapshot[25][41] , 
	\sa_snapshot[25][40] , \sa_snapshot[25][39] , \sa_snapshot[25][38] , 
	\sa_snapshot[25][37] , \sa_snapshot[25][36] , \sa_snapshot[25][35] , 
	\sa_snapshot[25][34] , \sa_snapshot[25][33] , \sa_snapshot[25][32] , 
	\sa_snapshot[25][31] , \sa_snapshot[25][30] , \sa_snapshot[25][29] , 
	\sa_snapshot[25][28] , \sa_snapshot[25][27] , \sa_snapshot[25][26] , 
	\sa_snapshot[25][25] , \sa_snapshot[25][24] , \sa_snapshot[25][23] , 
	\sa_snapshot[25][22] , \sa_snapshot[25][21] , \sa_snapshot[25][20] , 
	\sa_snapshot[25][19] , \sa_snapshot[25][18] , \sa_snapshot[25][17] , 
	\sa_snapshot[25][16] , \sa_snapshot[25][15] , \sa_snapshot[25][14] , 
	\sa_snapshot[25][13] , \sa_snapshot[25][12] , \sa_snapshot[25][11] , 
	\sa_snapshot[25][10] , \sa_snapshot[25][9] , \sa_snapshot[25][8] , 
	\sa_snapshot[25][7] , \sa_snapshot[25][6] , \sa_snapshot[25][5] , 
	\sa_snapshot[25][4] , \sa_snapshot[25][3] , \sa_snapshot[25][2] , 
	\sa_snapshot[25][1] , \sa_snapshot[25][0] , \sa_snapshot[24][63] , 
	\sa_snapshot[24][62] , \sa_snapshot[24][61] , \sa_snapshot[24][60] , 
	\sa_snapshot[24][59] , \sa_snapshot[24][58] , \sa_snapshot[24][57] , 
	\sa_snapshot[24][56] , \sa_snapshot[24][55] , \sa_snapshot[24][54] , 
	\sa_snapshot[24][53] , \sa_snapshot[24][52] , \sa_snapshot[24][51] , 
	\sa_snapshot[24][50] , \sa_snapshot[24][49] , \sa_snapshot[24][48] , 
	\sa_snapshot[24][47] , \sa_snapshot[24][46] , \sa_snapshot[24][45] , 
	\sa_snapshot[24][44] , \sa_snapshot[24][43] , \sa_snapshot[24][42] , 
	\sa_snapshot[24][41] , \sa_snapshot[24][40] , \sa_snapshot[24][39] , 
	\sa_snapshot[24][38] , \sa_snapshot[24][37] , \sa_snapshot[24][36] , 
	\sa_snapshot[24][35] , \sa_snapshot[24][34] , \sa_snapshot[24][33] , 
	\sa_snapshot[24][32] , \sa_snapshot[24][31] , \sa_snapshot[24][30] , 
	\sa_snapshot[24][29] , \sa_snapshot[24][28] , \sa_snapshot[24][27] , 
	\sa_snapshot[24][26] , \sa_snapshot[24][25] , \sa_snapshot[24][24] , 
	\sa_snapshot[24][23] , \sa_snapshot[24][22] , \sa_snapshot[24][21] , 
	\sa_snapshot[24][20] , \sa_snapshot[24][19] , \sa_snapshot[24][18] , 
	\sa_snapshot[24][17] , \sa_snapshot[24][16] , \sa_snapshot[24][15] , 
	\sa_snapshot[24][14] , \sa_snapshot[24][13] , \sa_snapshot[24][12] , 
	\sa_snapshot[24][11] , \sa_snapshot[24][10] , \sa_snapshot[24][9] , 
	\sa_snapshot[24][8] , \sa_snapshot[24][7] , \sa_snapshot[24][6] , 
	\sa_snapshot[24][5] , \sa_snapshot[24][4] , \sa_snapshot[24][3] , 
	\sa_snapshot[24][2] , \sa_snapshot[24][1] , \sa_snapshot[24][0] , 
	\sa_snapshot[23][63] , \sa_snapshot[23][62] , \sa_snapshot[23][61] , 
	\sa_snapshot[23][60] , \sa_snapshot[23][59] , \sa_snapshot[23][58] , 
	\sa_snapshot[23][57] , \sa_snapshot[23][56] , \sa_snapshot[23][55] , 
	\sa_snapshot[23][54] , \sa_snapshot[23][53] , \sa_snapshot[23][52] , 
	\sa_snapshot[23][51] , \sa_snapshot[23][50] , \sa_snapshot[23][49] , 
	\sa_snapshot[23][48] , \sa_snapshot[23][47] , \sa_snapshot[23][46] , 
	\sa_snapshot[23][45] , \sa_snapshot[23][44] , \sa_snapshot[23][43] , 
	\sa_snapshot[23][42] , \sa_snapshot[23][41] , \sa_snapshot[23][40] , 
	\sa_snapshot[23][39] , \sa_snapshot[23][38] , \sa_snapshot[23][37] , 
	\sa_snapshot[23][36] , \sa_snapshot[23][35] , \sa_snapshot[23][34] , 
	\sa_snapshot[23][33] , \sa_snapshot[23][32] , \sa_snapshot[23][31] , 
	\sa_snapshot[23][30] , \sa_snapshot[23][29] , \sa_snapshot[23][28] , 
	\sa_snapshot[23][27] , \sa_snapshot[23][26] , \sa_snapshot[23][25] , 
	\sa_snapshot[23][24] , \sa_snapshot[23][23] , \sa_snapshot[23][22] , 
	\sa_snapshot[23][21] , \sa_snapshot[23][20] , \sa_snapshot[23][19] , 
	\sa_snapshot[23][18] , \sa_snapshot[23][17] , \sa_snapshot[23][16] , 
	\sa_snapshot[23][15] , \sa_snapshot[23][14] , \sa_snapshot[23][13] , 
	\sa_snapshot[23][12] , \sa_snapshot[23][11] , \sa_snapshot[23][10] , 
	\sa_snapshot[23][9] , \sa_snapshot[23][8] , \sa_snapshot[23][7] , 
	\sa_snapshot[23][6] , \sa_snapshot[23][5] , \sa_snapshot[23][4] , 
	\sa_snapshot[23][3] , \sa_snapshot[23][2] , \sa_snapshot[23][1] , 
	\sa_snapshot[23][0] , \sa_snapshot[22][63] , \sa_snapshot[22][62] , 
	\sa_snapshot[22][61] , \sa_snapshot[22][60] , \sa_snapshot[22][59] , 
	\sa_snapshot[22][58] , \sa_snapshot[22][57] , \sa_snapshot[22][56] , 
	\sa_snapshot[22][55] , \sa_snapshot[22][54] , \sa_snapshot[22][53] , 
	\sa_snapshot[22][52] , \sa_snapshot[22][51] , \sa_snapshot[22][50] , 
	\sa_snapshot[22][49] , \sa_snapshot[22][48] , \sa_snapshot[22][47] , 
	\sa_snapshot[22][46] , \sa_snapshot[22][45] , \sa_snapshot[22][44] , 
	\sa_snapshot[22][43] , \sa_snapshot[22][42] , \sa_snapshot[22][41] , 
	\sa_snapshot[22][40] , \sa_snapshot[22][39] , \sa_snapshot[22][38] , 
	\sa_snapshot[22][37] , \sa_snapshot[22][36] , \sa_snapshot[22][35] , 
	\sa_snapshot[22][34] , \sa_snapshot[22][33] , \sa_snapshot[22][32] , 
	\sa_snapshot[22][31] , \sa_snapshot[22][30] , \sa_snapshot[22][29] , 
	\sa_snapshot[22][28] , \sa_snapshot[22][27] , \sa_snapshot[22][26] , 
	\sa_snapshot[22][25] , \sa_snapshot[22][24] , \sa_snapshot[22][23] , 
	\sa_snapshot[22][22] , \sa_snapshot[22][21] , \sa_snapshot[22][20] , 
	\sa_snapshot[22][19] , \sa_snapshot[22][18] , \sa_snapshot[22][17] , 
	\sa_snapshot[22][16] , \sa_snapshot[22][15] , \sa_snapshot[22][14] , 
	\sa_snapshot[22][13] , \sa_snapshot[22][12] , \sa_snapshot[22][11] , 
	\sa_snapshot[22][10] , \sa_snapshot[22][9] , \sa_snapshot[22][8] , 
	\sa_snapshot[22][7] , \sa_snapshot[22][6] , \sa_snapshot[22][5] , 
	\sa_snapshot[22][4] , \sa_snapshot[22][3] , \sa_snapshot[22][2] , 
	\sa_snapshot[22][1] , \sa_snapshot[22][0] , \sa_snapshot[21][63] , 
	\sa_snapshot[21][62] , \sa_snapshot[21][61] , \sa_snapshot[21][60] , 
	\sa_snapshot[21][59] , \sa_snapshot[21][58] , \sa_snapshot[21][57] , 
	\sa_snapshot[21][56] , \sa_snapshot[21][55] , \sa_snapshot[21][54] , 
	\sa_snapshot[21][53] , \sa_snapshot[21][52] , \sa_snapshot[21][51] , 
	\sa_snapshot[21][50] , \sa_snapshot[21][49] , \sa_snapshot[21][48] , 
	\sa_snapshot[21][47] , \sa_snapshot[21][46] , \sa_snapshot[21][45] , 
	\sa_snapshot[21][44] , \sa_snapshot[21][43] , \sa_snapshot[21][42] , 
	\sa_snapshot[21][41] , \sa_snapshot[21][40] , \sa_snapshot[21][39] , 
	\sa_snapshot[21][38] , \sa_snapshot[21][37] , \sa_snapshot[21][36] , 
	\sa_snapshot[21][35] , \sa_snapshot[21][34] , \sa_snapshot[21][33] , 
	\sa_snapshot[21][32] , \sa_snapshot[21][31] , \sa_snapshot[21][30] , 
	\sa_snapshot[21][29] , \sa_snapshot[21][28] , \sa_snapshot[21][27] , 
	\sa_snapshot[21][26] , \sa_snapshot[21][25] , \sa_snapshot[21][24] , 
	\sa_snapshot[21][23] , \sa_snapshot[21][22] , \sa_snapshot[21][21] , 
	\sa_snapshot[21][20] , \sa_snapshot[21][19] , \sa_snapshot[21][18] , 
	\sa_snapshot[21][17] , \sa_snapshot[21][16] , \sa_snapshot[21][15] , 
	\sa_snapshot[21][14] , \sa_snapshot[21][13] , \sa_snapshot[21][12] , 
	\sa_snapshot[21][11] , \sa_snapshot[21][10] , \sa_snapshot[21][9] , 
	\sa_snapshot[21][8] , \sa_snapshot[21][7] , \sa_snapshot[21][6] , 
	\sa_snapshot[21][5] , \sa_snapshot[21][4] , \sa_snapshot[21][3] , 
	\sa_snapshot[21][2] , \sa_snapshot[21][1] , \sa_snapshot[21][0] , 
	\sa_snapshot[20][63] , \sa_snapshot[20][62] , \sa_snapshot[20][61] , 
	\sa_snapshot[20][60] , \sa_snapshot[20][59] , \sa_snapshot[20][58] , 
	\sa_snapshot[20][57] , \sa_snapshot[20][56] , \sa_snapshot[20][55] , 
	\sa_snapshot[20][54] , \sa_snapshot[20][53] , \sa_snapshot[20][52] , 
	\sa_snapshot[20][51] , \sa_snapshot[20][50] , \sa_snapshot[20][49] , 
	\sa_snapshot[20][48] , \sa_snapshot[20][47] , \sa_snapshot[20][46] , 
	\sa_snapshot[20][45] , \sa_snapshot[20][44] , \sa_snapshot[20][43] , 
	\sa_snapshot[20][42] , \sa_snapshot[20][41] , \sa_snapshot[20][40] , 
	\sa_snapshot[20][39] , \sa_snapshot[20][38] , \sa_snapshot[20][37] , 
	\sa_snapshot[20][36] , \sa_snapshot[20][35] , \sa_snapshot[20][34] , 
	\sa_snapshot[20][33] , \sa_snapshot[20][32] , \sa_snapshot[20][31] , 
	\sa_snapshot[20][30] , \sa_snapshot[20][29] , \sa_snapshot[20][28] , 
	\sa_snapshot[20][27] , \sa_snapshot[20][26] , \sa_snapshot[20][25] , 
	\sa_snapshot[20][24] , \sa_snapshot[20][23] , \sa_snapshot[20][22] , 
	\sa_snapshot[20][21] , \sa_snapshot[20][20] , \sa_snapshot[20][19] , 
	\sa_snapshot[20][18] , \sa_snapshot[20][17] , \sa_snapshot[20][16] , 
	\sa_snapshot[20][15] , \sa_snapshot[20][14] , \sa_snapshot[20][13] , 
	\sa_snapshot[20][12] , \sa_snapshot[20][11] , \sa_snapshot[20][10] , 
	\sa_snapshot[20][9] , \sa_snapshot[20][8] , \sa_snapshot[20][7] , 
	\sa_snapshot[20][6] , \sa_snapshot[20][5] , \sa_snapshot[20][4] , 
	\sa_snapshot[20][3] , \sa_snapshot[20][2] , \sa_snapshot[20][1] , 
	\sa_snapshot[20][0] , \sa_snapshot[19][63] , \sa_snapshot[19][62] , 
	\sa_snapshot[19][61] , \sa_snapshot[19][60] , \sa_snapshot[19][59] , 
	\sa_snapshot[19][58] , \sa_snapshot[19][57] , \sa_snapshot[19][56] , 
	\sa_snapshot[19][55] , \sa_snapshot[19][54] , \sa_snapshot[19][53] , 
	\sa_snapshot[19][52] , \sa_snapshot[19][51] , \sa_snapshot[19][50] , 
	\sa_snapshot[19][49] , \sa_snapshot[19][48] , \sa_snapshot[19][47] , 
	\sa_snapshot[19][46] , \sa_snapshot[19][45] , \sa_snapshot[19][44] , 
	\sa_snapshot[19][43] , \sa_snapshot[19][42] , \sa_snapshot[19][41] , 
	\sa_snapshot[19][40] , \sa_snapshot[19][39] , \sa_snapshot[19][38] , 
	\sa_snapshot[19][37] , \sa_snapshot[19][36] , \sa_snapshot[19][35] , 
	\sa_snapshot[19][34] , \sa_snapshot[19][33] , \sa_snapshot[19][32] , 
	\sa_snapshot[19][31] , \sa_snapshot[19][30] , \sa_snapshot[19][29] , 
	\sa_snapshot[19][28] , \sa_snapshot[19][27] , \sa_snapshot[19][26] , 
	\sa_snapshot[19][25] , \sa_snapshot[19][24] , \sa_snapshot[19][23] , 
	\sa_snapshot[19][22] , \sa_snapshot[19][21] , \sa_snapshot[19][20] , 
	\sa_snapshot[19][19] , \sa_snapshot[19][18] , \sa_snapshot[19][17] , 
	\sa_snapshot[19][16] , \sa_snapshot[19][15] , \sa_snapshot[19][14] , 
	\sa_snapshot[19][13] , \sa_snapshot[19][12] , \sa_snapshot[19][11] , 
	\sa_snapshot[19][10] , \sa_snapshot[19][9] , \sa_snapshot[19][8] , 
	\sa_snapshot[19][7] , \sa_snapshot[19][6] , \sa_snapshot[19][5] , 
	\sa_snapshot[19][4] , \sa_snapshot[19][3] , \sa_snapshot[19][2] , 
	\sa_snapshot[19][1] , \sa_snapshot[19][0] , \sa_snapshot[18][63] , 
	\sa_snapshot[18][62] , \sa_snapshot[18][61] , \sa_snapshot[18][60] , 
	\sa_snapshot[18][59] , \sa_snapshot[18][58] , \sa_snapshot[18][57] , 
	\sa_snapshot[18][56] , \sa_snapshot[18][55] , \sa_snapshot[18][54] , 
	\sa_snapshot[18][53] , \sa_snapshot[18][52] , \sa_snapshot[18][51] , 
	\sa_snapshot[18][50] , \sa_snapshot[18][49] , \sa_snapshot[18][48] , 
	\sa_snapshot[18][47] , \sa_snapshot[18][46] , \sa_snapshot[18][45] , 
	\sa_snapshot[18][44] , \sa_snapshot[18][43] , \sa_snapshot[18][42] , 
	\sa_snapshot[18][41] , \sa_snapshot[18][40] , \sa_snapshot[18][39] , 
	\sa_snapshot[18][38] , \sa_snapshot[18][37] , \sa_snapshot[18][36] , 
	\sa_snapshot[18][35] , \sa_snapshot[18][34] , \sa_snapshot[18][33] , 
	\sa_snapshot[18][32] , \sa_snapshot[18][31] , \sa_snapshot[18][30] , 
	\sa_snapshot[18][29] , \sa_snapshot[18][28] , \sa_snapshot[18][27] , 
	\sa_snapshot[18][26] , \sa_snapshot[18][25] , \sa_snapshot[18][24] , 
	\sa_snapshot[18][23] , \sa_snapshot[18][22] , \sa_snapshot[18][21] , 
	\sa_snapshot[18][20] , \sa_snapshot[18][19] , \sa_snapshot[18][18] , 
	\sa_snapshot[18][17] , \sa_snapshot[18][16] , \sa_snapshot[18][15] , 
	\sa_snapshot[18][14] , \sa_snapshot[18][13] , \sa_snapshot[18][12] , 
	\sa_snapshot[18][11] , \sa_snapshot[18][10] , \sa_snapshot[18][9] , 
	\sa_snapshot[18][8] , \sa_snapshot[18][7] , \sa_snapshot[18][6] , 
	\sa_snapshot[18][5] , \sa_snapshot[18][4] , \sa_snapshot[18][3] , 
	\sa_snapshot[18][2] , \sa_snapshot[18][1] , \sa_snapshot[18][0] , 
	\sa_snapshot[17][63] , \sa_snapshot[17][62] , \sa_snapshot[17][61] , 
	\sa_snapshot[17][60] , \sa_snapshot[17][59] , \sa_snapshot[17][58] , 
	\sa_snapshot[17][57] , \sa_snapshot[17][56] , \sa_snapshot[17][55] , 
	\sa_snapshot[17][54] , \sa_snapshot[17][53] , \sa_snapshot[17][52] , 
	\sa_snapshot[17][51] , \sa_snapshot[17][50] , \sa_snapshot[17][49] , 
	\sa_snapshot[17][48] , \sa_snapshot[17][47] , \sa_snapshot[17][46] , 
	\sa_snapshot[17][45] , \sa_snapshot[17][44] , \sa_snapshot[17][43] , 
	\sa_snapshot[17][42] , \sa_snapshot[17][41] , \sa_snapshot[17][40] , 
	\sa_snapshot[17][39] , \sa_snapshot[17][38] , \sa_snapshot[17][37] , 
	\sa_snapshot[17][36] , \sa_snapshot[17][35] , \sa_snapshot[17][34] , 
	\sa_snapshot[17][33] , \sa_snapshot[17][32] , \sa_snapshot[17][31] , 
	\sa_snapshot[17][30] , \sa_snapshot[17][29] , \sa_snapshot[17][28] , 
	\sa_snapshot[17][27] , \sa_snapshot[17][26] , \sa_snapshot[17][25] , 
	\sa_snapshot[17][24] , \sa_snapshot[17][23] , \sa_snapshot[17][22] , 
	\sa_snapshot[17][21] , \sa_snapshot[17][20] , \sa_snapshot[17][19] , 
	\sa_snapshot[17][18] , \sa_snapshot[17][17] , \sa_snapshot[17][16] , 
	\sa_snapshot[17][15] , \sa_snapshot[17][14] , \sa_snapshot[17][13] , 
	\sa_snapshot[17][12] , \sa_snapshot[17][11] , \sa_snapshot[17][10] , 
	\sa_snapshot[17][9] , \sa_snapshot[17][8] , \sa_snapshot[17][7] , 
	\sa_snapshot[17][6] , \sa_snapshot[17][5] , \sa_snapshot[17][4] , 
	\sa_snapshot[17][3] , \sa_snapshot[17][2] , \sa_snapshot[17][1] , 
	\sa_snapshot[17][0] , \sa_snapshot[16][63] , \sa_snapshot[16][62] , 
	\sa_snapshot[16][61] , \sa_snapshot[16][60] , \sa_snapshot[16][59] , 
	\sa_snapshot[16][58] , \sa_snapshot[16][57] , \sa_snapshot[16][56] , 
	\sa_snapshot[16][55] , \sa_snapshot[16][54] , \sa_snapshot[16][53] , 
	\sa_snapshot[16][52] , \sa_snapshot[16][51] , \sa_snapshot[16][50] , 
	\sa_snapshot[16][49] , \sa_snapshot[16][48] , \sa_snapshot[16][47] , 
	\sa_snapshot[16][46] , \sa_snapshot[16][45] , \sa_snapshot[16][44] , 
	\sa_snapshot[16][43] , \sa_snapshot[16][42] , \sa_snapshot[16][41] , 
	\sa_snapshot[16][40] , \sa_snapshot[16][39] , \sa_snapshot[16][38] , 
	\sa_snapshot[16][37] , \sa_snapshot[16][36] , \sa_snapshot[16][35] , 
	\sa_snapshot[16][34] , \sa_snapshot[16][33] , \sa_snapshot[16][32] , 
	\sa_snapshot[16][31] , \sa_snapshot[16][30] , \sa_snapshot[16][29] , 
	\sa_snapshot[16][28] , \sa_snapshot[16][27] , \sa_snapshot[16][26] , 
	\sa_snapshot[16][25] , \sa_snapshot[16][24] , \sa_snapshot[16][23] , 
	\sa_snapshot[16][22] , \sa_snapshot[16][21] , \sa_snapshot[16][20] , 
	\sa_snapshot[16][19] , \sa_snapshot[16][18] , \sa_snapshot[16][17] , 
	\sa_snapshot[16][16] , \sa_snapshot[16][15] , \sa_snapshot[16][14] , 
	\sa_snapshot[16][13] , \sa_snapshot[16][12] , \sa_snapshot[16][11] , 
	\sa_snapshot[16][10] , \sa_snapshot[16][9] , \sa_snapshot[16][8] , 
	\sa_snapshot[16][7] , \sa_snapshot[16][6] , \sa_snapshot[16][5] , 
	\sa_snapshot[16][4] , \sa_snapshot[16][3] , \sa_snapshot[16][2] , 
	\sa_snapshot[16][1] , \sa_snapshot[16][0] , \sa_snapshot[15][63] , 
	\sa_snapshot[15][62] , \sa_snapshot[15][61] , \sa_snapshot[15][60] , 
	\sa_snapshot[15][59] , \sa_snapshot[15][58] , \sa_snapshot[15][57] , 
	\sa_snapshot[15][56] , \sa_snapshot[15][55] , \sa_snapshot[15][54] , 
	\sa_snapshot[15][53] , \sa_snapshot[15][52] , \sa_snapshot[15][51] , 
	\sa_snapshot[15][50] , \sa_snapshot[15][49] , \sa_snapshot[15][48] , 
	\sa_snapshot[15][47] , \sa_snapshot[15][46] , \sa_snapshot[15][45] , 
	\sa_snapshot[15][44] , \sa_snapshot[15][43] , \sa_snapshot[15][42] , 
	\sa_snapshot[15][41] , \sa_snapshot[15][40] , \sa_snapshot[15][39] , 
	\sa_snapshot[15][38] , \sa_snapshot[15][37] , \sa_snapshot[15][36] , 
	\sa_snapshot[15][35] , \sa_snapshot[15][34] , \sa_snapshot[15][33] , 
	\sa_snapshot[15][32] , \sa_snapshot[15][31] , \sa_snapshot[15][30] , 
	\sa_snapshot[15][29] , \sa_snapshot[15][28] , \sa_snapshot[15][27] , 
	\sa_snapshot[15][26] , \sa_snapshot[15][25] , \sa_snapshot[15][24] , 
	\sa_snapshot[15][23] , \sa_snapshot[15][22] , \sa_snapshot[15][21] , 
	\sa_snapshot[15][20] , \sa_snapshot[15][19] , \sa_snapshot[15][18] , 
	\sa_snapshot[15][17] , \sa_snapshot[15][16] , \sa_snapshot[15][15] , 
	\sa_snapshot[15][14] , \sa_snapshot[15][13] , \sa_snapshot[15][12] , 
	\sa_snapshot[15][11] , \sa_snapshot[15][10] , \sa_snapshot[15][9] , 
	\sa_snapshot[15][8] , \sa_snapshot[15][7] , \sa_snapshot[15][6] , 
	\sa_snapshot[15][5] , \sa_snapshot[15][4] , \sa_snapshot[15][3] , 
	\sa_snapshot[15][2] , \sa_snapshot[15][1] , \sa_snapshot[15][0] , 
	\sa_snapshot[14][63] , \sa_snapshot[14][62] , \sa_snapshot[14][61] , 
	\sa_snapshot[14][60] , \sa_snapshot[14][59] , \sa_snapshot[14][58] , 
	\sa_snapshot[14][57] , \sa_snapshot[14][56] , \sa_snapshot[14][55] , 
	\sa_snapshot[14][54] , \sa_snapshot[14][53] , \sa_snapshot[14][52] , 
	\sa_snapshot[14][51] , \sa_snapshot[14][50] , \sa_snapshot[14][49] , 
	\sa_snapshot[14][48] , \sa_snapshot[14][47] , \sa_snapshot[14][46] , 
	\sa_snapshot[14][45] , \sa_snapshot[14][44] , \sa_snapshot[14][43] , 
	\sa_snapshot[14][42] , \sa_snapshot[14][41] , \sa_snapshot[14][40] , 
	\sa_snapshot[14][39] , \sa_snapshot[14][38] , \sa_snapshot[14][37] , 
	\sa_snapshot[14][36] , \sa_snapshot[14][35] , \sa_snapshot[14][34] , 
	\sa_snapshot[14][33] , \sa_snapshot[14][32] , \sa_snapshot[14][31] , 
	\sa_snapshot[14][30] , \sa_snapshot[14][29] , \sa_snapshot[14][28] , 
	\sa_snapshot[14][27] , \sa_snapshot[14][26] , \sa_snapshot[14][25] , 
	\sa_snapshot[14][24] , \sa_snapshot[14][23] , \sa_snapshot[14][22] , 
	\sa_snapshot[14][21] , \sa_snapshot[14][20] , \sa_snapshot[14][19] , 
	\sa_snapshot[14][18] , \sa_snapshot[14][17] , \sa_snapshot[14][16] , 
	\sa_snapshot[14][15] , \sa_snapshot[14][14] , \sa_snapshot[14][13] , 
	\sa_snapshot[14][12] , \sa_snapshot[14][11] , \sa_snapshot[14][10] , 
	\sa_snapshot[14][9] , \sa_snapshot[14][8] , \sa_snapshot[14][7] , 
	\sa_snapshot[14][6] , \sa_snapshot[14][5] , \sa_snapshot[14][4] , 
	\sa_snapshot[14][3] , \sa_snapshot[14][2] , \sa_snapshot[14][1] , 
	\sa_snapshot[14][0] , \sa_snapshot[13][63] , \sa_snapshot[13][62] , 
	\sa_snapshot[13][61] , \sa_snapshot[13][60] , \sa_snapshot[13][59] , 
	\sa_snapshot[13][58] , \sa_snapshot[13][57] , \sa_snapshot[13][56] , 
	\sa_snapshot[13][55] , \sa_snapshot[13][54] , \sa_snapshot[13][53] , 
	\sa_snapshot[13][52] , \sa_snapshot[13][51] , \sa_snapshot[13][50] , 
	\sa_snapshot[13][49] , \sa_snapshot[13][48] , \sa_snapshot[13][47] , 
	\sa_snapshot[13][46] , \sa_snapshot[13][45] , \sa_snapshot[13][44] , 
	\sa_snapshot[13][43] , \sa_snapshot[13][42] , \sa_snapshot[13][41] , 
	\sa_snapshot[13][40] , \sa_snapshot[13][39] , \sa_snapshot[13][38] , 
	\sa_snapshot[13][37] , \sa_snapshot[13][36] , \sa_snapshot[13][35] , 
	\sa_snapshot[13][34] , \sa_snapshot[13][33] , \sa_snapshot[13][32] , 
	\sa_snapshot[13][31] , \sa_snapshot[13][30] , \sa_snapshot[13][29] , 
	\sa_snapshot[13][28] , \sa_snapshot[13][27] , \sa_snapshot[13][26] , 
	\sa_snapshot[13][25] , \sa_snapshot[13][24] , \sa_snapshot[13][23] , 
	\sa_snapshot[13][22] , \sa_snapshot[13][21] , \sa_snapshot[13][20] , 
	\sa_snapshot[13][19] , \sa_snapshot[13][18] , \sa_snapshot[13][17] , 
	\sa_snapshot[13][16] , \sa_snapshot[13][15] , \sa_snapshot[13][14] , 
	\sa_snapshot[13][13] , \sa_snapshot[13][12] , \sa_snapshot[13][11] , 
	\sa_snapshot[13][10] , \sa_snapshot[13][9] , \sa_snapshot[13][8] , 
	\sa_snapshot[13][7] , \sa_snapshot[13][6] , \sa_snapshot[13][5] , 
	\sa_snapshot[13][4] , \sa_snapshot[13][3] , \sa_snapshot[13][2] , 
	\sa_snapshot[13][1] , \sa_snapshot[13][0] , \sa_snapshot[12][63] , 
	\sa_snapshot[12][62] , \sa_snapshot[12][61] , \sa_snapshot[12][60] , 
	\sa_snapshot[12][59] , \sa_snapshot[12][58] , \sa_snapshot[12][57] , 
	\sa_snapshot[12][56] , \sa_snapshot[12][55] , \sa_snapshot[12][54] , 
	\sa_snapshot[12][53] , \sa_snapshot[12][52] , \sa_snapshot[12][51] , 
	\sa_snapshot[12][50] , \sa_snapshot[12][49] , \sa_snapshot[12][48] , 
	\sa_snapshot[12][47] , \sa_snapshot[12][46] , \sa_snapshot[12][45] , 
	\sa_snapshot[12][44] , \sa_snapshot[12][43] , \sa_snapshot[12][42] , 
	\sa_snapshot[12][41] , \sa_snapshot[12][40] , \sa_snapshot[12][39] , 
	\sa_snapshot[12][38] , \sa_snapshot[12][37] , \sa_snapshot[12][36] , 
	\sa_snapshot[12][35] , \sa_snapshot[12][34] , \sa_snapshot[12][33] , 
	\sa_snapshot[12][32] , \sa_snapshot[12][31] , \sa_snapshot[12][30] , 
	\sa_snapshot[12][29] , \sa_snapshot[12][28] , \sa_snapshot[12][27] , 
	\sa_snapshot[12][26] , \sa_snapshot[12][25] , \sa_snapshot[12][24] , 
	\sa_snapshot[12][23] , \sa_snapshot[12][22] , \sa_snapshot[12][21] , 
	\sa_snapshot[12][20] , \sa_snapshot[12][19] , \sa_snapshot[12][18] , 
	\sa_snapshot[12][17] , \sa_snapshot[12][16] , \sa_snapshot[12][15] , 
	\sa_snapshot[12][14] , \sa_snapshot[12][13] , \sa_snapshot[12][12] , 
	\sa_snapshot[12][11] , \sa_snapshot[12][10] , \sa_snapshot[12][9] , 
	\sa_snapshot[12][8] , \sa_snapshot[12][7] , \sa_snapshot[12][6] , 
	\sa_snapshot[12][5] , \sa_snapshot[12][4] , \sa_snapshot[12][3] , 
	\sa_snapshot[12][2] , \sa_snapshot[12][1] , \sa_snapshot[12][0] , 
	\sa_snapshot[11][63] , \sa_snapshot[11][62] , \sa_snapshot[11][61] , 
	\sa_snapshot[11][60] , \sa_snapshot[11][59] , \sa_snapshot[11][58] , 
	\sa_snapshot[11][57] , \sa_snapshot[11][56] , \sa_snapshot[11][55] , 
	\sa_snapshot[11][54] , \sa_snapshot[11][53] , \sa_snapshot[11][52] , 
	\sa_snapshot[11][51] , \sa_snapshot[11][50] , \sa_snapshot[11][49] , 
	\sa_snapshot[11][48] , \sa_snapshot[11][47] , \sa_snapshot[11][46] , 
	\sa_snapshot[11][45] , \sa_snapshot[11][44] , \sa_snapshot[11][43] , 
	\sa_snapshot[11][42] , \sa_snapshot[11][41] , \sa_snapshot[11][40] , 
	\sa_snapshot[11][39] , \sa_snapshot[11][38] , \sa_snapshot[11][37] , 
	\sa_snapshot[11][36] , \sa_snapshot[11][35] , \sa_snapshot[11][34] , 
	\sa_snapshot[11][33] , \sa_snapshot[11][32] , \sa_snapshot[11][31] , 
	\sa_snapshot[11][30] , \sa_snapshot[11][29] , \sa_snapshot[11][28] , 
	\sa_snapshot[11][27] , \sa_snapshot[11][26] , \sa_snapshot[11][25] , 
	\sa_snapshot[11][24] , \sa_snapshot[11][23] , \sa_snapshot[11][22] , 
	\sa_snapshot[11][21] , \sa_snapshot[11][20] , \sa_snapshot[11][19] , 
	\sa_snapshot[11][18] , \sa_snapshot[11][17] , \sa_snapshot[11][16] , 
	\sa_snapshot[11][15] , \sa_snapshot[11][14] , \sa_snapshot[11][13] , 
	\sa_snapshot[11][12] , \sa_snapshot[11][11] , \sa_snapshot[11][10] , 
	\sa_snapshot[11][9] , \sa_snapshot[11][8] , \sa_snapshot[11][7] , 
	\sa_snapshot[11][6] , \sa_snapshot[11][5] , \sa_snapshot[11][4] , 
	\sa_snapshot[11][3] , \sa_snapshot[11][2] , \sa_snapshot[11][1] , 
	\sa_snapshot[11][0] , \sa_snapshot[10][63] , \sa_snapshot[10][62] , 
	\sa_snapshot[10][61] , \sa_snapshot[10][60] , \sa_snapshot[10][59] , 
	\sa_snapshot[10][58] , \sa_snapshot[10][57] , \sa_snapshot[10][56] , 
	\sa_snapshot[10][55] , \sa_snapshot[10][54] , \sa_snapshot[10][53] , 
	\sa_snapshot[10][52] , \sa_snapshot[10][51] , \sa_snapshot[10][50] , 
	\sa_snapshot[10][49] , \sa_snapshot[10][48] , \sa_snapshot[10][47] , 
	\sa_snapshot[10][46] , \sa_snapshot[10][45] , \sa_snapshot[10][44] , 
	\sa_snapshot[10][43] , \sa_snapshot[10][42] , \sa_snapshot[10][41] , 
	\sa_snapshot[10][40] , \sa_snapshot[10][39] , \sa_snapshot[10][38] , 
	\sa_snapshot[10][37] , \sa_snapshot[10][36] , \sa_snapshot[10][35] , 
	\sa_snapshot[10][34] , \sa_snapshot[10][33] , \sa_snapshot[10][32] , 
	\sa_snapshot[10][31] , \sa_snapshot[10][30] , \sa_snapshot[10][29] , 
	\sa_snapshot[10][28] , \sa_snapshot[10][27] , \sa_snapshot[10][26] , 
	\sa_snapshot[10][25] , \sa_snapshot[10][24] , \sa_snapshot[10][23] , 
	\sa_snapshot[10][22] , \sa_snapshot[10][21] , \sa_snapshot[10][20] , 
	\sa_snapshot[10][19] , \sa_snapshot[10][18] , \sa_snapshot[10][17] , 
	\sa_snapshot[10][16] , \sa_snapshot[10][15] , \sa_snapshot[10][14] , 
	\sa_snapshot[10][13] , \sa_snapshot[10][12] , \sa_snapshot[10][11] , 
	\sa_snapshot[10][10] , \sa_snapshot[10][9] , \sa_snapshot[10][8] , 
	\sa_snapshot[10][7] , \sa_snapshot[10][6] , \sa_snapshot[10][5] , 
	\sa_snapshot[10][4] , \sa_snapshot[10][3] , \sa_snapshot[10][2] , 
	\sa_snapshot[10][1] , \sa_snapshot[10][0] , \sa_snapshot[9][63] , 
	\sa_snapshot[9][62] , \sa_snapshot[9][61] , \sa_snapshot[9][60] , 
	\sa_snapshot[9][59] , \sa_snapshot[9][58] , \sa_snapshot[9][57] , 
	\sa_snapshot[9][56] , \sa_snapshot[9][55] , \sa_snapshot[9][54] , 
	\sa_snapshot[9][53] , \sa_snapshot[9][52] , \sa_snapshot[9][51] , 
	\sa_snapshot[9][50] , \sa_snapshot[9][49] , \sa_snapshot[9][48] , 
	\sa_snapshot[9][47] , \sa_snapshot[9][46] , \sa_snapshot[9][45] , 
	\sa_snapshot[9][44] , \sa_snapshot[9][43] , \sa_snapshot[9][42] , 
	\sa_snapshot[9][41] , \sa_snapshot[9][40] , \sa_snapshot[9][39] , 
	\sa_snapshot[9][38] , \sa_snapshot[9][37] , \sa_snapshot[9][36] , 
	\sa_snapshot[9][35] , \sa_snapshot[9][34] , \sa_snapshot[9][33] , 
	\sa_snapshot[9][32] , \sa_snapshot[9][31] , \sa_snapshot[9][30] , 
	\sa_snapshot[9][29] , \sa_snapshot[9][28] , \sa_snapshot[9][27] , 
	\sa_snapshot[9][26] , \sa_snapshot[9][25] , \sa_snapshot[9][24] , 
	\sa_snapshot[9][23] , \sa_snapshot[9][22] , \sa_snapshot[9][21] , 
	\sa_snapshot[9][20] , \sa_snapshot[9][19] , \sa_snapshot[9][18] , 
	\sa_snapshot[9][17] , \sa_snapshot[9][16] , \sa_snapshot[9][15] , 
	\sa_snapshot[9][14] , \sa_snapshot[9][13] , \sa_snapshot[9][12] , 
	\sa_snapshot[9][11] , \sa_snapshot[9][10] , \sa_snapshot[9][9] , 
	\sa_snapshot[9][8] , \sa_snapshot[9][7] , \sa_snapshot[9][6] , 
	\sa_snapshot[9][5] , \sa_snapshot[9][4] , \sa_snapshot[9][3] , 
	\sa_snapshot[9][2] , \sa_snapshot[9][1] , \sa_snapshot[9][0] , 
	\sa_snapshot[8][63] , \sa_snapshot[8][62] , \sa_snapshot[8][61] , 
	\sa_snapshot[8][60] , \sa_snapshot[8][59] , \sa_snapshot[8][58] , 
	\sa_snapshot[8][57] , \sa_snapshot[8][56] , \sa_snapshot[8][55] , 
	\sa_snapshot[8][54] , \sa_snapshot[8][53] , \sa_snapshot[8][52] , 
	\sa_snapshot[8][51] , \sa_snapshot[8][50] , \sa_snapshot[8][49] , 
	\sa_snapshot[8][48] , \sa_snapshot[8][47] , \sa_snapshot[8][46] , 
	\sa_snapshot[8][45] , \sa_snapshot[8][44] , \sa_snapshot[8][43] , 
	\sa_snapshot[8][42] , \sa_snapshot[8][41] , \sa_snapshot[8][40] , 
	\sa_snapshot[8][39] , \sa_snapshot[8][38] , \sa_snapshot[8][37] , 
	\sa_snapshot[8][36] , \sa_snapshot[8][35] , \sa_snapshot[8][34] , 
	\sa_snapshot[8][33] , \sa_snapshot[8][32] , \sa_snapshot[8][31] , 
	\sa_snapshot[8][30] , \sa_snapshot[8][29] , \sa_snapshot[8][28] , 
	\sa_snapshot[8][27] , \sa_snapshot[8][26] , \sa_snapshot[8][25] , 
	\sa_snapshot[8][24] , \sa_snapshot[8][23] , \sa_snapshot[8][22] , 
	\sa_snapshot[8][21] , \sa_snapshot[8][20] , \sa_snapshot[8][19] , 
	\sa_snapshot[8][18] , \sa_snapshot[8][17] , \sa_snapshot[8][16] , 
	\sa_snapshot[8][15] , \sa_snapshot[8][14] , \sa_snapshot[8][13] , 
	\sa_snapshot[8][12] , \sa_snapshot[8][11] , \sa_snapshot[8][10] , 
	\sa_snapshot[8][9] , \sa_snapshot[8][8] , \sa_snapshot[8][7] , 
	\sa_snapshot[8][6] , \sa_snapshot[8][5] , \sa_snapshot[8][4] , 
	\sa_snapshot[8][3] , \sa_snapshot[8][2] , \sa_snapshot[8][1] , 
	\sa_snapshot[8][0] , \sa_snapshot[7][63] , \sa_snapshot[7][62] , 
	\sa_snapshot[7][61] , \sa_snapshot[7][60] , \sa_snapshot[7][59] , 
	\sa_snapshot[7][58] , \sa_snapshot[7][57] , \sa_snapshot[7][56] , 
	\sa_snapshot[7][55] , \sa_snapshot[7][54] , \sa_snapshot[7][53] , 
	\sa_snapshot[7][52] , \sa_snapshot[7][51] , \sa_snapshot[7][50] , 
	\sa_snapshot[7][49] , \sa_snapshot[7][48] , \sa_snapshot[7][47] , 
	\sa_snapshot[7][46] , \sa_snapshot[7][45] , \sa_snapshot[7][44] , 
	\sa_snapshot[7][43] , \sa_snapshot[7][42] , \sa_snapshot[7][41] , 
	\sa_snapshot[7][40] , \sa_snapshot[7][39] , \sa_snapshot[7][38] , 
	\sa_snapshot[7][37] , \sa_snapshot[7][36] , \sa_snapshot[7][35] , 
	\sa_snapshot[7][34] , \sa_snapshot[7][33] , \sa_snapshot[7][32] , 
	\sa_snapshot[7][31] , \sa_snapshot[7][30] , \sa_snapshot[7][29] , 
	\sa_snapshot[7][28] , \sa_snapshot[7][27] , \sa_snapshot[7][26] , 
	\sa_snapshot[7][25] , \sa_snapshot[7][24] , \sa_snapshot[7][23] , 
	\sa_snapshot[7][22] , \sa_snapshot[7][21] , \sa_snapshot[7][20] , 
	\sa_snapshot[7][19] , \sa_snapshot[7][18] , \sa_snapshot[7][17] , 
	\sa_snapshot[7][16] , \sa_snapshot[7][15] , \sa_snapshot[7][14] , 
	\sa_snapshot[7][13] , \sa_snapshot[7][12] , \sa_snapshot[7][11] , 
	\sa_snapshot[7][10] , \sa_snapshot[7][9] , \sa_snapshot[7][8] , 
	\sa_snapshot[7][7] , \sa_snapshot[7][6] , \sa_snapshot[7][5] , 
	\sa_snapshot[7][4] , \sa_snapshot[7][3] , \sa_snapshot[7][2] , 
	\sa_snapshot[7][1] , \sa_snapshot[7][0] , \sa_snapshot[6][63] , 
	\sa_snapshot[6][62] , \sa_snapshot[6][61] , \sa_snapshot[6][60] , 
	\sa_snapshot[6][59] , \sa_snapshot[6][58] , \sa_snapshot[6][57] , 
	\sa_snapshot[6][56] , \sa_snapshot[6][55] , \sa_snapshot[6][54] , 
	\sa_snapshot[6][53] , \sa_snapshot[6][52] , \sa_snapshot[6][51] , 
	\sa_snapshot[6][50] , \sa_snapshot[6][49] , \sa_snapshot[6][48] , 
	\sa_snapshot[6][47] , \sa_snapshot[6][46] , \sa_snapshot[6][45] , 
	\sa_snapshot[6][44] , \sa_snapshot[6][43] , \sa_snapshot[6][42] , 
	\sa_snapshot[6][41] , \sa_snapshot[6][40] , \sa_snapshot[6][39] , 
	\sa_snapshot[6][38] , \sa_snapshot[6][37] , \sa_snapshot[6][36] , 
	\sa_snapshot[6][35] , \sa_snapshot[6][34] , \sa_snapshot[6][33] , 
	\sa_snapshot[6][32] , \sa_snapshot[6][31] , \sa_snapshot[6][30] , 
	\sa_snapshot[6][29] , \sa_snapshot[6][28] , \sa_snapshot[6][27] , 
	\sa_snapshot[6][26] , \sa_snapshot[6][25] , \sa_snapshot[6][24] , 
	\sa_snapshot[6][23] , \sa_snapshot[6][22] , \sa_snapshot[6][21] , 
	\sa_snapshot[6][20] , \sa_snapshot[6][19] , \sa_snapshot[6][18] , 
	\sa_snapshot[6][17] , \sa_snapshot[6][16] , \sa_snapshot[6][15] , 
	\sa_snapshot[6][14] , \sa_snapshot[6][13] , \sa_snapshot[6][12] , 
	\sa_snapshot[6][11] , \sa_snapshot[6][10] , \sa_snapshot[6][9] , 
	\sa_snapshot[6][8] , \sa_snapshot[6][7] , \sa_snapshot[6][6] , 
	\sa_snapshot[6][5] , \sa_snapshot[6][4] , \sa_snapshot[6][3] , 
	\sa_snapshot[6][2] , \sa_snapshot[6][1] , \sa_snapshot[6][0] , 
	\sa_snapshot[5][63] , \sa_snapshot[5][62] , \sa_snapshot[5][61] , 
	\sa_snapshot[5][60] , \sa_snapshot[5][59] , \sa_snapshot[5][58] , 
	\sa_snapshot[5][57] , \sa_snapshot[5][56] , \sa_snapshot[5][55] , 
	\sa_snapshot[5][54] , \sa_snapshot[5][53] , \sa_snapshot[5][52] , 
	\sa_snapshot[5][51] , \sa_snapshot[5][50] , \sa_snapshot[5][49] , 
	\sa_snapshot[5][48] , \sa_snapshot[5][47] , \sa_snapshot[5][46] , 
	\sa_snapshot[5][45] , \sa_snapshot[5][44] , \sa_snapshot[5][43] , 
	\sa_snapshot[5][42] , \sa_snapshot[5][41] , \sa_snapshot[5][40] , 
	\sa_snapshot[5][39] , \sa_snapshot[5][38] , \sa_snapshot[5][37] , 
	\sa_snapshot[5][36] , \sa_snapshot[5][35] , \sa_snapshot[5][34] , 
	\sa_snapshot[5][33] , \sa_snapshot[5][32] , \sa_snapshot[5][31] , 
	\sa_snapshot[5][30] , \sa_snapshot[5][29] , \sa_snapshot[5][28] , 
	\sa_snapshot[5][27] , \sa_snapshot[5][26] , \sa_snapshot[5][25] , 
	\sa_snapshot[5][24] , \sa_snapshot[5][23] , \sa_snapshot[5][22] , 
	\sa_snapshot[5][21] , \sa_snapshot[5][20] , \sa_snapshot[5][19] , 
	\sa_snapshot[5][18] , \sa_snapshot[5][17] , \sa_snapshot[5][16] , 
	\sa_snapshot[5][15] , \sa_snapshot[5][14] , \sa_snapshot[5][13] , 
	\sa_snapshot[5][12] , \sa_snapshot[5][11] , \sa_snapshot[5][10] , 
	\sa_snapshot[5][9] , \sa_snapshot[5][8] , \sa_snapshot[5][7] , 
	\sa_snapshot[5][6] , \sa_snapshot[5][5] , \sa_snapshot[5][4] , 
	\sa_snapshot[5][3] , \sa_snapshot[5][2] , \sa_snapshot[5][1] , 
	\sa_snapshot[5][0] , \sa_snapshot[4][63] , \sa_snapshot[4][62] , 
	\sa_snapshot[4][61] , \sa_snapshot[4][60] , \sa_snapshot[4][59] , 
	\sa_snapshot[4][58] , \sa_snapshot[4][57] , \sa_snapshot[4][56] , 
	\sa_snapshot[4][55] , \sa_snapshot[4][54] , \sa_snapshot[4][53] , 
	\sa_snapshot[4][52] , \sa_snapshot[4][51] , \sa_snapshot[4][50] , 
	\sa_snapshot[4][49] , \sa_snapshot[4][48] , \sa_snapshot[4][47] , 
	\sa_snapshot[4][46] , \sa_snapshot[4][45] , \sa_snapshot[4][44] , 
	\sa_snapshot[4][43] , \sa_snapshot[4][42] , \sa_snapshot[4][41] , 
	\sa_snapshot[4][40] , \sa_snapshot[4][39] , \sa_snapshot[4][38] , 
	\sa_snapshot[4][37] , \sa_snapshot[4][36] , \sa_snapshot[4][35] , 
	\sa_snapshot[4][34] , \sa_snapshot[4][33] , \sa_snapshot[4][32] , 
	\sa_snapshot[4][31] , \sa_snapshot[4][30] , \sa_snapshot[4][29] , 
	\sa_snapshot[4][28] , \sa_snapshot[4][27] , \sa_snapshot[4][26] , 
	\sa_snapshot[4][25] , \sa_snapshot[4][24] , \sa_snapshot[4][23] , 
	\sa_snapshot[4][22] , \sa_snapshot[4][21] , \sa_snapshot[4][20] , 
	\sa_snapshot[4][19] , \sa_snapshot[4][18] , \sa_snapshot[4][17] , 
	\sa_snapshot[4][16] , \sa_snapshot[4][15] , \sa_snapshot[4][14] , 
	\sa_snapshot[4][13] , \sa_snapshot[4][12] , \sa_snapshot[4][11] , 
	\sa_snapshot[4][10] , \sa_snapshot[4][9] , \sa_snapshot[4][8] , 
	\sa_snapshot[4][7] , \sa_snapshot[4][6] , \sa_snapshot[4][5] , 
	\sa_snapshot[4][4] , \sa_snapshot[4][3] , \sa_snapshot[4][2] , 
	\sa_snapshot[4][1] , \sa_snapshot[4][0] , \sa_snapshot[3][63] , 
	\sa_snapshot[3][62] , \sa_snapshot[3][61] , \sa_snapshot[3][60] , 
	\sa_snapshot[3][59] , \sa_snapshot[3][58] , \sa_snapshot[3][57] , 
	\sa_snapshot[3][56] , \sa_snapshot[3][55] , \sa_snapshot[3][54] , 
	\sa_snapshot[3][53] , \sa_snapshot[3][52] , \sa_snapshot[3][51] , 
	\sa_snapshot[3][50] , \sa_snapshot[3][49] , \sa_snapshot[3][48] , 
	\sa_snapshot[3][47] , \sa_snapshot[3][46] , \sa_snapshot[3][45] , 
	\sa_snapshot[3][44] , \sa_snapshot[3][43] , \sa_snapshot[3][42] , 
	\sa_snapshot[3][41] , \sa_snapshot[3][40] , \sa_snapshot[3][39] , 
	\sa_snapshot[3][38] , \sa_snapshot[3][37] , \sa_snapshot[3][36] , 
	\sa_snapshot[3][35] , \sa_snapshot[3][34] , \sa_snapshot[3][33] , 
	\sa_snapshot[3][32] , \sa_snapshot[3][31] , \sa_snapshot[3][30] , 
	\sa_snapshot[3][29] , \sa_snapshot[3][28] , \sa_snapshot[3][27] , 
	\sa_snapshot[3][26] , \sa_snapshot[3][25] , \sa_snapshot[3][24] , 
	\sa_snapshot[3][23] , \sa_snapshot[3][22] , \sa_snapshot[3][21] , 
	\sa_snapshot[3][20] , \sa_snapshot[3][19] , \sa_snapshot[3][18] , 
	\sa_snapshot[3][17] , \sa_snapshot[3][16] , \sa_snapshot[3][15] , 
	\sa_snapshot[3][14] , \sa_snapshot[3][13] , \sa_snapshot[3][12] , 
	\sa_snapshot[3][11] , \sa_snapshot[3][10] , \sa_snapshot[3][9] , 
	\sa_snapshot[3][8] , \sa_snapshot[3][7] , \sa_snapshot[3][6] , 
	\sa_snapshot[3][5] , \sa_snapshot[3][4] , \sa_snapshot[3][3] , 
	\sa_snapshot[3][2] , \sa_snapshot[3][1] , \sa_snapshot[3][0] , 
	\sa_snapshot[2][63] , \sa_snapshot[2][62] , \sa_snapshot[2][61] , 
	\sa_snapshot[2][60] , \sa_snapshot[2][59] , \sa_snapshot[2][58] , 
	\sa_snapshot[2][57] , \sa_snapshot[2][56] , \sa_snapshot[2][55] , 
	\sa_snapshot[2][54] , \sa_snapshot[2][53] , \sa_snapshot[2][52] , 
	\sa_snapshot[2][51] , \sa_snapshot[2][50] , \sa_snapshot[2][49] , 
	\sa_snapshot[2][48] , \sa_snapshot[2][47] , \sa_snapshot[2][46] , 
	\sa_snapshot[2][45] , \sa_snapshot[2][44] , \sa_snapshot[2][43] , 
	\sa_snapshot[2][42] , \sa_snapshot[2][41] , \sa_snapshot[2][40] , 
	\sa_snapshot[2][39] , \sa_snapshot[2][38] , \sa_snapshot[2][37] , 
	\sa_snapshot[2][36] , \sa_snapshot[2][35] , \sa_snapshot[2][34] , 
	\sa_snapshot[2][33] , \sa_snapshot[2][32] , \sa_snapshot[2][31] , 
	\sa_snapshot[2][30] , \sa_snapshot[2][29] , \sa_snapshot[2][28] , 
	\sa_snapshot[2][27] , \sa_snapshot[2][26] , \sa_snapshot[2][25] , 
	\sa_snapshot[2][24] , \sa_snapshot[2][23] , \sa_snapshot[2][22] , 
	\sa_snapshot[2][21] , \sa_snapshot[2][20] , \sa_snapshot[2][19] , 
	\sa_snapshot[2][18] , \sa_snapshot[2][17] , \sa_snapshot[2][16] , 
	\sa_snapshot[2][15] , \sa_snapshot[2][14] , \sa_snapshot[2][13] , 
	\sa_snapshot[2][12] , \sa_snapshot[2][11] , \sa_snapshot[2][10] , 
	\sa_snapshot[2][9] , \sa_snapshot[2][8] , \sa_snapshot[2][7] , 
	\sa_snapshot[2][6] , \sa_snapshot[2][5] , \sa_snapshot[2][4] , 
	\sa_snapshot[2][3] , \sa_snapshot[2][2] , \sa_snapshot[2][1] , 
	\sa_snapshot[2][0] , \sa_snapshot[1][63] , \sa_snapshot[1][62] , 
	\sa_snapshot[1][61] , \sa_snapshot[1][60] , \sa_snapshot[1][59] , 
	\sa_snapshot[1][58] , \sa_snapshot[1][57] , \sa_snapshot[1][56] , 
	\sa_snapshot[1][55] , \sa_snapshot[1][54] , \sa_snapshot[1][53] , 
	\sa_snapshot[1][52] , \sa_snapshot[1][51] , \sa_snapshot[1][50] , 
	\sa_snapshot[1][49] , \sa_snapshot[1][48] , \sa_snapshot[1][47] , 
	\sa_snapshot[1][46] , \sa_snapshot[1][45] , \sa_snapshot[1][44] , 
	\sa_snapshot[1][43] , \sa_snapshot[1][42] , \sa_snapshot[1][41] , 
	\sa_snapshot[1][40] , \sa_snapshot[1][39] , \sa_snapshot[1][38] , 
	\sa_snapshot[1][37] , \sa_snapshot[1][36] , \sa_snapshot[1][35] , 
	\sa_snapshot[1][34] , \sa_snapshot[1][33] , \sa_snapshot[1][32] , 
	\sa_snapshot[1][31] , \sa_snapshot[1][30] , \sa_snapshot[1][29] , 
	\sa_snapshot[1][28] , \sa_snapshot[1][27] , \sa_snapshot[1][26] , 
	\sa_snapshot[1][25] , \sa_snapshot[1][24] , \sa_snapshot[1][23] , 
	\sa_snapshot[1][22] , \sa_snapshot[1][21] , \sa_snapshot[1][20] , 
	\sa_snapshot[1][19] , \sa_snapshot[1][18] , \sa_snapshot[1][17] , 
	\sa_snapshot[1][16] , \sa_snapshot[1][15] , \sa_snapshot[1][14] , 
	\sa_snapshot[1][13] , \sa_snapshot[1][12] , \sa_snapshot[1][11] , 
	\sa_snapshot[1][10] , \sa_snapshot[1][9] , \sa_snapshot[1][8] , 
	\sa_snapshot[1][7] , \sa_snapshot[1][6] , \sa_snapshot[1][5] , 
	\sa_snapshot[1][4] , \sa_snapshot[1][3] , \sa_snapshot[1][2] , 
	\sa_snapshot[1][1] , \sa_snapshot[1][0] , \sa_snapshot[0][63] , 
	\sa_snapshot[0][62] , \sa_snapshot[0][61] , \sa_snapshot[0][60] , 
	\sa_snapshot[0][59] , \sa_snapshot[0][58] , \sa_snapshot[0][57] , 
	\sa_snapshot[0][56] , \sa_snapshot[0][55] , \sa_snapshot[0][54] , 
	\sa_snapshot[0][53] , \sa_snapshot[0][52] , \sa_snapshot[0][51] , 
	\sa_snapshot[0][50] , \sa_snapshot[0][49] , \sa_snapshot[0][48] , 
	\sa_snapshot[0][47] , \sa_snapshot[0][46] , \sa_snapshot[0][45] , 
	\sa_snapshot[0][44] , \sa_snapshot[0][43] , \sa_snapshot[0][42] , 
	\sa_snapshot[0][41] , \sa_snapshot[0][40] , \sa_snapshot[0][39] , 
	\sa_snapshot[0][38] , \sa_snapshot[0][37] , \sa_snapshot[0][36] , 
	\sa_snapshot[0][35] , \sa_snapshot[0][34] , \sa_snapshot[0][33] , 
	\sa_snapshot[0][32] , \sa_snapshot[0][31] , \sa_snapshot[0][30] , 
	\sa_snapshot[0][29] , \sa_snapshot[0][28] , \sa_snapshot[0][27] , 
	\sa_snapshot[0][26] , \sa_snapshot[0][25] , \sa_snapshot[0][24] , 
	\sa_snapshot[0][23] , \sa_snapshot[0][22] , \sa_snapshot[0][21] , 
	\sa_snapshot[0][20] , \sa_snapshot[0][19] , \sa_snapshot[0][18] , 
	\sa_snapshot[0][17] , \sa_snapshot[0][16] , \sa_snapshot[0][15] , 
	\sa_snapshot[0][14] , \sa_snapshot[0][13] , \sa_snapshot[0][12] , 
	\sa_snapshot[0][11] , \sa_snapshot[0][10] , \sa_snapshot[0][9] , 
	\sa_snapshot[0][8] , \sa_snapshot[0][7] , \sa_snapshot[0][6] , 
	\sa_snapshot[0][5] , \sa_snapshot[0][4] , \sa_snapshot[0][3] , 
	\sa_snapshot[0][2] , \sa_snapshot[0][1] , \sa_snapshot[0][0] }), 
	.sa_count( { \sa_count[31][63] , \sa_count[31][62] , 
	\sa_count[31][61] , \sa_count[31][60] , \sa_count[31][59] , 
	\sa_count[31][58] , \sa_count[31][57] , \sa_count[31][56] , 
	\sa_count[31][55] , \sa_count[31][54] , \sa_count[31][53] , 
	\sa_count[31][52] , \sa_count[31][51] , \sa_count[31][50] , 
	\sa_count[31][49] , \sa_count[31][48] , \sa_count[31][47] , 
	\sa_count[31][46] , \sa_count[31][45] , \sa_count[31][44] , 
	\sa_count[31][43] , \sa_count[31][42] , \sa_count[31][41] , 
	\sa_count[31][40] , \sa_count[31][39] , \sa_count[31][38] , 
	\sa_count[31][37] , \sa_count[31][36] , \sa_count[31][35] , 
	\sa_count[31][34] , \sa_count[31][33] , \sa_count[31][32] , 
	\sa_count[31][31] , \sa_count[31][30] , \sa_count[31][29] , 
	\sa_count[31][28] , \sa_count[31][27] , \sa_count[31][26] , 
	\sa_count[31][25] , \sa_count[31][24] , \sa_count[31][23] , 
	\sa_count[31][22] , \sa_count[31][21] , \sa_count[31][20] , 
	\sa_count[31][19] , \sa_count[31][18] , \sa_count[31][17] , 
	\sa_count[31][16] , \sa_count[31][15] , \sa_count[31][14] , 
	\sa_count[31][13] , \sa_count[31][12] , \sa_count[31][11] , 
	\sa_count[31][10] , \sa_count[31][9] , \sa_count[31][8] , 
	\sa_count[31][7] , \sa_count[31][6] , \sa_count[31][5] , 
	\sa_count[31][4] , \sa_count[31][3] , \sa_count[31][2] , 
	\sa_count[31][1] , \sa_count[31][0] , \sa_count[30][63] , 
	\sa_count[30][62] , \sa_count[30][61] , \sa_count[30][60] , 
	\sa_count[30][59] , \sa_count[30][58] , \sa_count[30][57] , 
	\sa_count[30][56] , \sa_count[30][55] , \sa_count[30][54] , 
	\sa_count[30][53] , \sa_count[30][52] , \sa_count[30][51] , 
	\sa_count[30][50] , \sa_count[30][49] , \sa_count[30][48] , 
	\sa_count[30][47] , \sa_count[30][46] , \sa_count[30][45] , 
	\sa_count[30][44] , \sa_count[30][43] , \sa_count[30][42] , 
	\sa_count[30][41] , \sa_count[30][40] , \sa_count[30][39] , 
	\sa_count[30][38] , \sa_count[30][37] , \sa_count[30][36] , 
	\sa_count[30][35] , \sa_count[30][34] , \sa_count[30][33] , 
	\sa_count[30][32] , \sa_count[30][31] , \sa_count[30][30] , 
	\sa_count[30][29] , \sa_count[30][28] , \sa_count[30][27] , 
	\sa_count[30][26] , \sa_count[30][25] , \sa_count[30][24] , 
	\sa_count[30][23] , \sa_count[30][22] , \sa_count[30][21] , 
	\sa_count[30][20] , \sa_count[30][19] , \sa_count[30][18] , 
	\sa_count[30][17] , \sa_count[30][16] , \sa_count[30][15] , 
	\sa_count[30][14] , \sa_count[30][13] , \sa_count[30][12] , 
	\sa_count[30][11] , \sa_count[30][10] , \sa_count[30][9] , 
	\sa_count[30][8] , \sa_count[30][7] , \sa_count[30][6] , 
	\sa_count[30][5] , \sa_count[30][4] , \sa_count[30][3] , 
	\sa_count[30][2] , \sa_count[30][1] , \sa_count[30][0] , 
	\sa_count[29][63] , \sa_count[29][62] , \sa_count[29][61] , 
	\sa_count[29][60] , \sa_count[29][59] , \sa_count[29][58] , 
	\sa_count[29][57] , \sa_count[29][56] , \sa_count[29][55] , 
	\sa_count[29][54] , \sa_count[29][53] , \sa_count[29][52] , 
	\sa_count[29][51] , \sa_count[29][50] , \sa_count[29][49] , 
	\sa_count[29][48] , \sa_count[29][47] , \sa_count[29][46] , 
	\sa_count[29][45] , \sa_count[29][44] , \sa_count[29][43] , 
	\sa_count[29][42] , \sa_count[29][41] , \sa_count[29][40] , 
	\sa_count[29][39] , \sa_count[29][38] , \sa_count[29][37] , 
	\sa_count[29][36] , \sa_count[29][35] , \sa_count[29][34] , 
	\sa_count[29][33] , \sa_count[29][32] , \sa_count[29][31] , 
	\sa_count[29][30] , \sa_count[29][29] , \sa_count[29][28] , 
	\sa_count[29][27] , \sa_count[29][26] , \sa_count[29][25] , 
	\sa_count[29][24] , \sa_count[29][23] , \sa_count[29][22] , 
	\sa_count[29][21] , \sa_count[29][20] , \sa_count[29][19] , 
	\sa_count[29][18] , \sa_count[29][17] , \sa_count[29][16] , 
	\sa_count[29][15] , \sa_count[29][14] , \sa_count[29][13] , 
	\sa_count[29][12] , \sa_count[29][11] , \sa_count[29][10] , 
	\sa_count[29][9] , \sa_count[29][8] , \sa_count[29][7] , 
	\sa_count[29][6] , \sa_count[29][5] , \sa_count[29][4] , 
	\sa_count[29][3] , \sa_count[29][2] , \sa_count[29][1] , 
	\sa_count[29][0] , \sa_count[28][63] , \sa_count[28][62] , 
	\sa_count[28][61] , \sa_count[28][60] , \sa_count[28][59] , 
	\sa_count[28][58] , \sa_count[28][57] , \sa_count[28][56] , 
	\sa_count[28][55] , \sa_count[28][54] , \sa_count[28][53] , 
	\sa_count[28][52] , \sa_count[28][51] , \sa_count[28][50] , 
	\sa_count[28][49] , \sa_count[28][48] , \sa_count[28][47] , 
	\sa_count[28][46] , \sa_count[28][45] , \sa_count[28][44] , 
	\sa_count[28][43] , \sa_count[28][42] , \sa_count[28][41] , 
	\sa_count[28][40] , \sa_count[28][39] , \sa_count[28][38] , 
	\sa_count[28][37] , \sa_count[28][36] , \sa_count[28][35] , 
	\sa_count[28][34] , \sa_count[28][33] , \sa_count[28][32] , 
	\sa_count[28][31] , \sa_count[28][30] , \sa_count[28][29] , 
	\sa_count[28][28] , \sa_count[28][27] , \sa_count[28][26] , 
	\sa_count[28][25] , \sa_count[28][24] , \sa_count[28][23] , 
	\sa_count[28][22] , \sa_count[28][21] , \sa_count[28][20] , 
	\sa_count[28][19] , \sa_count[28][18] , \sa_count[28][17] , 
	\sa_count[28][16] , \sa_count[28][15] , \sa_count[28][14] , 
	\sa_count[28][13] , \sa_count[28][12] , \sa_count[28][11] , 
	\sa_count[28][10] , \sa_count[28][9] , \sa_count[28][8] , 
	\sa_count[28][7] , \sa_count[28][6] , \sa_count[28][5] , 
	\sa_count[28][4] , \sa_count[28][3] , \sa_count[28][2] , 
	\sa_count[28][1] , \sa_count[28][0] , \sa_count[27][63] , 
	\sa_count[27][62] , \sa_count[27][61] , \sa_count[27][60] , 
	\sa_count[27][59] , \sa_count[27][58] , \sa_count[27][57] , 
	\sa_count[27][56] , \sa_count[27][55] , \sa_count[27][54] , 
	\sa_count[27][53] , \sa_count[27][52] , \sa_count[27][51] , 
	\sa_count[27][50] , \sa_count[27][49] , \sa_count[27][48] , 
	\sa_count[27][47] , \sa_count[27][46] , \sa_count[27][45] , 
	\sa_count[27][44] , \sa_count[27][43] , \sa_count[27][42] , 
	\sa_count[27][41] , \sa_count[27][40] , \sa_count[27][39] , 
	\sa_count[27][38] , \sa_count[27][37] , \sa_count[27][36] , 
	\sa_count[27][35] , \sa_count[27][34] , \sa_count[27][33] , 
	\sa_count[27][32] , \sa_count[27][31] , \sa_count[27][30] , 
	\sa_count[27][29] , \sa_count[27][28] , \sa_count[27][27] , 
	\sa_count[27][26] , \sa_count[27][25] , \sa_count[27][24] , 
	\sa_count[27][23] , \sa_count[27][22] , \sa_count[27][21] , 
	\sa_count[27][20] , \sa_count[27][19] , \sa_count[27][18] , 
	\sa_count[27][17] , \sa_count[27][16] , \sa_count[27][15] , 
	\sa_count[27][14] , \sa_count[27][13] , \sa_count[27][12] , 
	\sa_count[27][11] , \sa_count[27][10] , \sa_count[27][9] , 
	\sa_count[27][8] , \sa_count[27][7] , \sa_count[27][6] , 
	\sa_count[27][5] , \sa_count[27][4] , \sa_count[27][3] , 
	\sa_count[27][2] , \sa_count[27][1] , \sa_count[27][0] , 
	\sa_count[26][63] , \sa_count[26][62] , \sa_count[26][61] , 
	\sa_count[26][60] , \sa_count[26][59] , \sa_count[26][58] , 
	\sa_count[26][57] , \sa_count[26][56] , \sa_count[26][55] , 
	\sa_count[26][54] , \sa_count[26][53] , \sa_count[26][52] , 
	\sa_count[26][51] , \sa_count[26][50] , \sa_count[26][49] , 
	\sa_count[26][48] , \sa_count[26][47] , \sa_count[26][46] , 
	\sa_count[26][45] , \sa_count[26][44] , \sa_count[26][43] , 
	\sa_count[26][42] , \sa_count[26][41] , \sa_count[26][40] , 
	\sa_count[26][39] , \sa_count[26][38] , \sa_count[26][37] , 
	\sa_count[26][36] , \sa_count[26][35] , \sa_count[26][34] , 
	\sa_count[26][33] , \sa_count[26][32] , \sa_count[26][31] , 
	\sa_count[26][30] , \sa_count[26][29] , \sa_count[26][28] , 
	\sa_count[26][27] , \sa_count[26][26] , \sa_count[26][25] , 
	\sa_count[26][24] , \sa_count[26][23] , \sa_count[26][22] , 
	\sa_count[26][21] , \sa_count[26][20] , \sa_count[26][19] , 
	\sa_count[26][18] , \sa_count[26][17] , \sa_count[26][16] , 
	\sa_count[26][15] , \sa_count[26][14] , \sa_count[26][13] , 
	\sa_count[26][12] , \sa_count[26][11] , \sa_count[26][10] , 
	\sa_count[26][9] , \sa_count[26][8] , \sa_count[26][7] , 
	\sa_count[26][6] , \sa_count[26][5] , \sa_count[26][4] , 
	\sa_count[26][3] , \sa_count[26][2] , \sa_count[26][1] , 
	\sa_count[26][0] , \sa_count[25][63] , \sa_count[25][62] , 
	\sa_count[25][61] , \sa_count[25][60] , \sa_count[25][59] , 
	\sa_count[25][58] , \sa_count[25][57] , \sa_count[25][56] , 
	\sa_count[25][55] , \sa_count[25][54] , \sa_count[25][53] , 
	\sa_count[25][52] , \sa_count[25][51] , \sa_count[25][50] , 
	\sa_count[25][49] , \sa_count[25][48] , \sa_count[25][47] , 
	\sa_count[25][46] , \sa_count[25][45] , \sa_count[25][44] , 
	\sa_count[25][43] , \sa_count[25][42] , \sa_count[25][41] , 
	\sa_count[25][40] , \sa_count[25][39] , \sa_count[25][38] , 
	\sa_count[25][37] , \sa_count[25][36] , \sa_count[25][35] , 
	\sa_count[25][34] , \sa_count[25][33] , \sa_count[25][32] , 
	\sa_count[25][31] , \sa_count[25][30] , \sa_count[25][29] , 
	\sa_count[25][28] , \sa_count[25][27] , \sa_count[25][26] , 
	\sa_count[25][25] , \sa_count[25][24] , \sa_count[25][23] , 
	\sa_count[25][22] , \sa_count[25][21] , \sa_count[25][20] , 
	\sa_count[25][19] , \sa_count[25][18] , \sa_count[25][17] , 
	\sa_count[25][16] , \sa_count[25][15] , \sa_count[25][14] , 
	\sa_count[25][13] , \sa_count[25][12] , \sa_count[25][11] , 
	\sa_count[25][10] , \sa_count[25][9] , \sa_count[25][8] , 
	\sa_count[25][7] , \sa_count[25][6] , \sa_count[25][5] , 
	\sa_count[25][4] , \sa_count[25][3] , \sa_count[25][2] , 
	\sa_count[25][1] , \sa_count[25][0] , \sa_count[24][63] , 
	\sa_count[24][62] , \sa_count[24][61] , \sa_count[24][60] , 
	\sa_count[24][59] , \sa_count[24][58] , \sa_count[24][57] , 
	\sa_count[24][56] , \sa_count[24][55] , \sa_count[24][54] , 
	\sa_count[24][53] , \sa_count[24][52] , \sa_count[24][51] , 
	\sa_count[24][50] , \sa_count[24][49] , \sa_count[24][48] , 
	\sa_count[24][47] , \sa_count[24][46] , \sa_count[24][45] , 
	\sa_count[24][44] , \sa_count[24][43] , \sa_count[24][42] , 
	\sa_count[24][41] , \sa_count[24][40] , \sa_count[24][39] , 
	\sa_count[24][38] , \sa_count[24][37] , \sa_count[24][36] , 
	\sa_count[24][35] , \sa_count[24][34] , \sa_count[24][33] , 
	\sa_count[24][32] , \sa_count[24][31] , \sa_count[24][30] , 
	\sa_count[24][29] , \sa_count[24][28] , \sa_count[24][27] , 
	\sa_count[24][26] , \sa_count[24][25] , \sa_count[24][24] , 
	\sa_count[24][23] , \sa_count[24][22] , \sa_count[24][21] , 
	\sa_count[24][20] , \sa_count[24][19] , \sa_count[24][18] , 
	\sa_count[24][17] , \sa_count[24][16] , \sa_count[24][15] , 
	\sa_count[24][14] , \sa_count[24][13] , \sa_count[24][12] , 
	\sa_count[24][11] , \sa_count[24][10] , \sa_count[24][9] , 
	\sa_count[24][8] , \sa_count[24][7] , \sa_count[24][6] , 
	\sa_count[24][5] , \sa_count[24][4] , \sa_count[24][3] , 
	\sa_count[24][2] , \sa_count[24][1] , \sa_count[24][0] , 
	\sa_count[23][63] , \sa_count[23][62] , \sa_count[23][61] , 
	\sa_count[23][60] , \sa_count[23][59] , \sa_count[23][58] , 
	\sa_count[23][57] , \sa_count[23][56] , \sa_count[23][55] , 
	\sa_count[23][54] , \sa_count[23][53] , \sa_count[23][52] , 
	\sa_count[23][51] , \sa_count[23][50] , \sa_count[23][49] , 
	\sa_count[23][48] , \sa_count[23][47] , \sa_count[23][46] , 
	\sa_count[23][45] , \sa_count[23][44] , \sa_count[23][43] , 
	\sa_count[23][42] , \sa_count[23][41] , \sa_count[23][40] , 
	\sa_count[23][39] , \sa_count[23][38] , \sa_count[23][37] , 
	\sa_count[23][36] , \sa_count[23][35] , \sa_count[23][34] , 
	\sa_count[23][33] , \sa_count[23][32] , \sa_count[23][31] , 
	\sa_count[23][30] , \sa_count[23][29] , \sa_count[23][28] , 
	\sa_count[23][27] , \sa_count[23][26] , \sa_count[23][25] , 
	\sa_count[23][24] , \sa_count[23][23] , \sa_count[23][22] , 
	\sa_count[23][21] , \sa_count[23][20] , \sa_count[23][19] , 
	\sa_count[23][18] , \sa_count[23][17] , \sa_count[23][16] , 
	\sa_count[23][15] , \sa_count[23][14] , \sa_count[23][13] , 
	\sa_count[23][12] , \sa_count[23][11] , \sa_count[23][10] , 
	\sa_count[23][9] , \sa_count[23][8] , \sa_count[23][7] , 
	\sa_count[23][6] , \sa_count[23][5] , \sa_count[23][4] , 
	\sa_count[23][3] , \sa_count[23][2] , \sa_count[23][1] , 
	\sa_count[23][0] , \sa_count[22][63] , \sa_count[22][62] , 
	\sa_count[22][61] , \sa_count[22][60] , \sa_count[22][59] , 
	\sa_count[22][58] , \sa_count[22][57] , \sa_count[22][56] , 
	\sa_count[22][55] , \sa_count[22][54] , \sa_count[22][53] , 
	\sa_count[22][52] , \sa_count[22][51] , \sa_count[22][50] , 
	\sa_count[22][49] , \sa_count[22][48] , \sa_count[22][47] , 
	\sa_count[22][46] , \sa_count[22][45] , \sa_count[22][44] , 
	\sa_count[22][43] , \sa_count[22][42] , \sa_count[22][41] , 
	\sa_count[22][40] , \sa_count[22][39] , \sa_count[22][38] , 
	\sa_count[22][37] , \sa_count[22][36] , \sa_count[22][35] , 
	\sa_count[22][34] , \sa_count[22][33] , \sa_count[22][32] , 
	\sa_count[22][31] , \sa_count[22][30] , \sa_count[22][29] , 
	\sa_count[22][28] , \sa_count[22][27] , \sa_count[22][26] , 
	\sa_count[22][25] , \sa_count[22][24] , \sa_count[22][23] , 
	\sa_count[22][22] , \sa_count[22][21] , \sa_count[22][20] , 
	\sa_count[22][19] , \sa_count[22][18] , \sa_count[22][17] , 
	\sa_count[22][16] , \sa_count[22][15] , \sa_count[22][14] , 
	\sa_count[22][13] , \sa_count[22][12] , \sa_count[22][11] , 
	\sa_count[22][10] , \sa_count[22][9] , \sa_count[22][8] , 
	\sa_count[22][7] , \sa_count[22][6] , \sa_count[22][5] , 
	\sa_count[22][4] , \sa_count[22][3] , \sa_count[22][2] , 
	\sa_count[22][1] , \sa_count[22][0] , \sa_count[21][63] , 
	\sa_count[21][62] , \sa_count[21][61] , \sa_count[21][60] , 
	\sa_count[21][59] , \sa_count[21][58] , \sa_count[21][57] , 
	\sa_count[21][56] , \sa_count[21][55] , \sa_count[21][54] , 
	\sa_count[21][53] , \sa_count[21][52] , \sa_count[21][51] , 
	\sa_count[21][50] , \sa_count[21][49] , \sa_count[21][48] , 
	\sa_count[21][47] , \sa_count[21][46] , \sa_count[21][45] , 
	\sa_count[21][44] , \sa_count[21][43] , \sa_count[21][42] , 
	\sa_count[21][41] , \sa_count[21][40] , \sa_count[21][39] , 
	\sa_count[21][38] , \sa_count[21][37] , \sa_count[21][36] , 
	\sa_count[21][35] , \sa_count[21][34] , \sa_count[21][33] , 
	\sa_count[21][32] , \sa_count[21][31] , \sa_count[21][30] , 
	\sa_count[21][29] , \sa_count[21][28] , \sa_count[21][27] , 
	\sa_count[21][26] , \sa_count[21][25] , \sa_count[21][24] , 
	\sa_count[21][23] , \sa_count[21][22] , \sa_count[21][21] , 
	\sa_count[21][20] , \sa_count[21][19] , \sa_count[21][18] , 
	\sa_count[21][17] , \sa_count[21][16] , \sa_count[21][15] , 
	\sa_count[21][14] , \sa_count[21][13] , \sa_count[21][12] , 
	\sa_count[21][11] , \sa_count[21][10] , \sa_count[21][9] , 
	\sa_count[21][8] , \sa_count[21][7] , \sa_count[21][6] , 
	\sa_count[21][5] , \sa_count[21][4] , \sa_count[21][3] , 
	\sa_count[21][2] , \sa_count[21][1] , \sa_count[21][0] , 
	\sa_count[20][63] , \sa_count[20][62] , \sa_count[20][61] , 
	\sa_count[20][60] , \sa_count[20][59] , \sa_count[20][58] , 
	\sa_count[20][57] , \sa_count[20][56] , \sa_count[20][55] , 
	\sa_count[20][54] , \sa_count[20][53] , \sa_count[20][52] , 
	\sa_count[20][51] , \sa_count[20][50] , \sa_count[20][49] , 
	\sa_count[20][48] , \sa_count[20][47] , \sa_count[20][46] , 
	\sa_count[20][45] , \sa_count[20][44] , \sa_count[20][43] , 
	\sa_count[20][42] , \sa_count[20][41] , \sa_count[20][40] , 
	\sa_count[20][39] , \sa_count[20][38] , \sa_count[20][37] , 
	\sa_count[20][36] , \sa_count[20][35] , \sa_count[20][34] , 
	\sa_count[20][33] , \sa_count[20][32] , \sa_count[20][31] , 
	\sa_count[20][30] , \sa_count[20][29] , \sa_count[20][28] , 
	\sa_count[20][27] , \sa_count[20][26] , \sa_count[20][25] , 
	\sa_count[20][24] , \sa_count[20][23] , \sa_count[20][22] , 
	\sa_count[20][21] , \sa_count[20][20] , \sa_count[20][19] , 
	\sa_count[20][18] , \sa_count[20][17] , \sa_count[20][16] , 
	\sa_count[20][15] , \sa_count[20][14] , \sa_count[20][13] , 
	\sa_count[20][12] , \sa_count[20][11] , \sa_count[20][10] , 
	\sa_count[20][9] , \sa_count[20][8] , \sa_count[20][7] , 
	\sa_count[20][6] , \sa_count[20][5] , \sa_count[20][4] , 
	\sa_count[20][3] , \sa_count[20][2] , \sa_count[20][1] , 
	\sa_count[20][0] , \sa_count[19][63] , \sa_count[19][62] , 
	\sa_count[19][61] , \sa_count[19][60] , \sa_count[19][59] , 
	\sa_count[19][58] , \sa_count[19][57] , \sa_count[19][56] , 
	\sa_count[19][55] , \sa_count[19][54] , \sa_count[19][53] , 
	\sa_count[19][52] , \sa_count[19][51] , \sa_count[19][50] , 
	\sa_count[19][49] , \sa_count[19][48] , \sa_count[19][47] , 
	\sa_count[19][46] , \sa_count[19][45] , \sa_count[19][44] , 
	\sa_count[19][43] , \sa_count[19][42] , \sa_count[19][41] , 
	\sa_count[19][40] , \sa_count[19][39] , \sa_count[19][38] , 
	\sa_count[19][37] , \sa_count[19][36] , \sa_count[19][35] , 
	\sa_count[19][34] , \sa_count[19][33] , \sa_count[19][32] , 
	\sa_count[19][31] , \sa_count[19][30] , \sa_count[19][29] , 
	\sa_count[19][28] , \sa_count[19][27] , \sa_count[19][26] , 
	\sa_count[19][25] , \sa_count[19][24] , \sa_count[19][23] , 
	\sa_count[19][22] , \sa_count[19][21] , \sa_count[19][20] , 
	\sa_count[19][19] , \sa_count[19][18] , \sa_count[19][17] , 
	\sa_count[19][16] , \sa_count[19][15] , \sa_count[19][14] , 
	\sa_count[19][13] , \sa_count[19][12] , \sa_count[19][11] , 
	\sa_count[19][10] , \sa_count[19][9] , \sa_count[19][8] , 
	\sa_count[19][7] , \sa_count[19][6] , \sa_count[19][5] , 
	\sa_count[19][4] , \sa_count[19][3] , \sa_count[19][2] , 
	\sa_count[19][1] , \sa_count[19][0] , \sa_count[18][63] , 
	\sa_count[18][62] , \sa_count[18][61] , \sa_count[18][60] , 
	\sa_count[18][59] , \sa_count[18][58] , \sa_count[18][57] , 
	\sa_count[18][56] , \sa_count[18][55] , \sa_count[18][54] , 
	\sa_count[18][53] , \sa_count[18][52] , \sa_count[18][51] , 
	\sa_count[18][50] , \sa_count[18][49] , \sa_count[18][48] , 
	\sa_count[18][47] , \sa_count[18][46] , \sa_count[18][45] , 
	\sa_count[18][44] , \sa_count[18][43] , \sa_count[18][42] , 
	\sa_count[18][41] , \sa_count[18][40] , \sa_count[18][39] , 
	\sa_count[18][38] , \sa_count[18][37] , \sa_count[18][36] , 
	\sa_count[18][35] , \sa_count[18][34] , \sa_count[18][33] , 
	\sa_count[18][32] , \sa_count[18][31] , \sa_count[18][30] , 
	\sa_count[18][29] , \sa_count[18][28] , \sa_count[18][27] , 
	\sa_count[18][26] , \sa_count[18][25] , \sa_count[18][24] , 
	\sa_count[18][23] , \sa_count[18][22] , \sa_count[18][21] , 
	\sa_count[18][20] , \sa_count[18][19] , \sa_count[18][18] , 
	\sa_count[18][17] , \sa_count[18][16] , \sa_count[18][15] , 
	\sa_count[18][14] , \sa_count[18][13] , \sa_count[18][12] , 
	\sa_count[18][11] , \sa_count[18][10] , \sa_count[18][9] , 
	\sa_count[18][8] , \sa_count[18][7] , \sa_count[18][6] , 
	\sa_count[18][5] , \sa_count[18][4] , \sa_count[18][3] , 
	\sa_count[18][2] , \sa_count[18][1] , \sa_count[18][0] , 
	\sa_count[17][63] , \sa_count[17][62] , \sa_count[17][61] , 
	\sa_count[17][60] , \sa_count[17][59] , \sa_count[17][58] , 
	\sa_count[17][57] , \sa_count[17][56] , \sa_count[17][55] , 
	\sa_count[17][54] , \sa_count[17][53] , \sa_count[17][52] , 
	\sa_count[17][51] , \sa_count[17][50] , \sa_count[17][49] , 
	\sa_count[17][48] , \sa_count[17][47] , \sa_count[17][46] , 
	\sa_count[17][45] , \sa_count[17][44] , \sa_count[17][43] , 
	\sa_count[17][42] , \sa_count[17][41] , \sa_count[17][40] , 
	\sa_count[17][39] , \sa_count[17][38] , \sa_count[17][37] , 
	\sa_count[17][36] , \sa_count[17][35] , \sa_count[17][34] , 
	\sa_count[17][33] , \sa_count[17][32] , \sa_count[17][31] , 
	\sa_count[17][30] , \sa_count[17][29] , \sa_count[17][28] , 
	\sa_count[17][27] , \sa_count[17][26] , \sa_count[17][25] , 
	\sa_count[17][24] , \sa_count[17][23] , \sa_count[17][22] , 
	\sa_count[17][21] , \sa_count[17][20] , \sa_count[17][19] , 
	\sa_count[17][18] , \sa_count[17][17] , \sa_count[17][16] , 
	\sa_count[17][15] , \sa_count[17][14] , \sa_count[17][13] , 
	\sa_count[17][12] , \sa_count[17][11] , \sa_count[17][10] , 
	\sa_count[17][9] , \sa_count[17][8] , \sa_count[17][7] , 
	\sa_count[17][6] , \sa_count[17][5] , \sa_count[17][4] , 
	\sa_count[17][3] , \sa_count[17][2] , \sa_count[17][1] , 
	\sa_count[17][0] , \sa_count[16][63] , \sa_count[16][62] , 
	\sa_count[16][61] , \sa_count[16][60] , \sa_count[16][59] , 
	\sa_count[16][58] , \sa_count[16][57] , \sa_count[16][56] , 
	\sa_count[16][55] , \sa_count[16][54] , \sa_count[16][53] , 
	\sa_count[16][52] , \sa_count[16][51] , \sa_count[16][50] , 
	\sa_count[16][49] , \sa_count[16][48] , \sa_count[16][47] , 
	\sa_count[16][46] , \sa_count[16][45] , \sa_count[16][44] , 
	\sa_count[16][43] , \sa_count[16][42] , \sa_count[16][41] , 
	\sa_count[16][40] , \sa_count[16][39] , \sa_count[16][38] , 
	\sa_count[16][37] , \sa_count[16][36] , \sa_count[16][35] , 
	\sa_count[16][34] , \sa_count[16][33] , \sa_count[16][32] , 
	\sa_count[16][31] , \sa_count[16][30] , \sa_count[16][29] , 
	\sa_count[16][28] , \sa_count[16][27] , \sa_count[16][26] , 
	\sa_count[16][25] , \sa_count[16][24] , \sa_count[16][23] , 
	\sa_count[16][22] , \sa_count[16][21] , \sa_count[16][20] , 
	\sa_count[16][19] , \sa_count[16][18] , \sa_count[16][17] , 
	\sa_count[16][16] , \sa_count[16][15] , \sa_count[16][14] , 
	\sa_count[16][13] , \sa_count[16][12] , \sa_count[16][11] , 
	\sa_count[16][10] , \sa_count[16][9] , \sa_count[16][8] , 
	\sa_count[16][7] , \sa_count[16][6] , \sa_count[16][5] , 
	\sa_count[16][4] , \sa_count[16][3] , \sa_count[16][2] , 
	\sa_count[16][1] , \sa_count[16][0] , \sa_count[15][63] , 
	\sa_count[15][62] , \sa_count[15][61] , \sa_count[15][60] , 
	\sa_count[15][59] , \sa_count[15][58] , \sa_count[15][57] , 
	\sa_count[15][56] , \sa_count[15][55] , \sa_count[15][54] , 
	\sa_count[15][53] , \sa_count[15][52] , \sa_count[15][51] , 
	\sa_count[15][50] , \sa_count[15][49] , \sa_count[15][48] , 
	\sa_count[15][47] , \sa_count[15][46] , \sa_count[15][45] , 
	\sa_count[15][44] , \sa_count[15][43] , \sa_count[15][42] , 
	\sa_count[15][41] , \sa_count[15][40] , \sa_count[15][39] , 
	\sa_count[15][38] , \sa_count[15][37] , \sa_count[15][36] , 
	\sa_count[15][35] , \sa_count[15][34] , \sa_count[15][33] , 
	\sa_count[15][32] , \sa_count[15][31] , \sa_count[15][30] , 
	\sa_count[15][29] , \sa_count[15][28] , \sa_count[15][27] , 
	\sa_count[15][26] , \sa_count[15][25] , \sa_count[15][24] , 
	\sa_count[15][23] , \sa_count[15][22] , \sa_count[15][21] , 
	\sa_count[15][20] , \sa_count[15][19] , \sa_count[15][18] , 
	\sa_count[15][17] , \sa_count[15][16] , \sa_count[15][15] , 
	\sa_count[15][14] , \sa_count[15][13] , \sa_count[15][12] , 
	\sa_count[15][11] , \sa_count[15][10] , \sa_count[15][9] , 
	\sa_count[15][8] , \sa_count[15][7] , \sa_count[15][6] , 
	\sa_count[15][5] , \sa_count[15][4] , \sa_count[15][3] , 
	\sa_count[15][2] , \sa_count[15][1] , \sa_count[15][0] , 
	\sa_count[14][63] , \sa_count[14][62] , \sa_count[14][61] , 
	\sa_count[14][60] , \sa_count[14][59] , \sa_count[14][58] , 
	\sa_count[14][57] , \sa_count[14][56] , \sa_count[14][55] , 
	\sa_count[14][54] , \sa_count[14][53] , \sa_count[14][52] , 
	\sa_count[14][51] , \sa_count[14][50] , \sa_count[14][49] , 
	\sa_count[14][48] , \sa_count[14][47] , \sa_count[14][46] , 
	\sa_count[14][45] , \sa_count[14][44] , \sa_count[14][43] , 
	\sa_count[14][42] , \sa_count[14][41] , \sa_count[14][40] , 
	\sa_count[14][39] , \sa_count[14][38] , \sa_count[14][37] , 
	\sa_count[14][36] , \sa_count[14][35] , \sa_count[14][34] , 
	\sa_count[14][33] , \sa_count[14][32] , \sa_count[14][31] , 
	\sa_count[14][30] , \sa_count[14][29] , \sa_count[14][28] , 
	\sa_count[14][27] , \sa_count[14][26] , \sa_count[14][25] , 
	\sa_count[14][24] , \sa_count[14][23] , \sa_count[14][22] , 
	\sa_count[14][21] , \sa_count[14][20] , \sa_count[14][19] , 
	\sa_count[14][18] , \sa_count[14][17] , \sa_count[14][16] , 
	\sa_count[14][15] , \sa_count[14][14] , \sa_count[14][13] , 
	\sa_count[14][12] , \sa_count[14][11] , \sa_count[14][10] , 
	\sa_count[14][9] , \sa_count[14][8] , \sa_count[14][7] , 
	\sa_count[14][6] , \sa_count[14][5] , \sa_count[14][4] , 
	\sa_count[14][3] , \sa_count[14][2] , \sa_count[14][1] , 
	\sa_count[14][0] , \sa_count[13][63] , \sa_count[13][62] , 
	\sa_count[13][61] , \sa_count[13][60] , \sa_count[13][59] , 
	\sa_count[13][58] , \sa_count[13][57] , \sa_count[13][56] , 
	\sa_count[13][55] , \sa_count[13][54] , \sa_count[13][53] , 
	\sa_count[13][52] , \sa_count[13][51] , \sa_count[13][50] , 
	\sa_count[13][49] , \sa_count[13][48] , \sa_count[13][47] , 
	\sa_count[13][46] , \sa_count[13][45] , \sa_count[13][44] , 
	\sa_count[13][43] , \sa_count[13][42] , \sa_count[13][41] , 
	\sa_count[13][40] , \sa_count[13][39] , \sa_count[13][38] , 
	\sa_count[13][37] , \sa_count[13][36] , \sa_count[13][35] , 
	\sa_count[13][34] , \sa_count[13][33] , \sa_count[13][32] , 
	\sa_count[13][31] , \sa_count[13][30] , \sa_count[13][29] , 
	\sa_count[13][28] , \sa_count[13][27] , \sa_count[13][26] , 
	\sa_count[13][25] , \sa_count[13][24] , \sa_count[13][23] , 
	\sa_count[13][22] , \sa_count[13][21] , \sa_count[13][20] , 
	\sa_count[13][19] , \sa_count[13][18] , \sa_count[13][17] , 
	\sa_count[13][16] , \sa_count[13][15] , \sa_count[13][14] , 
	\sa_count[13][13] , \sa_count[13][12] , \sa_count[13][11] , 
	\sa_count[13][10] , \sa_count[13][9] , \sa_count[13][8] , 
	\sa_count[13][7] , \sa_count[13][6] , \sa_count[13][5] , 
	\sa_count[13][4] , \sa_count[13][3] , \sa_count[13][2] , 
	\sa_count[13][1] , \sa_count[13][0] , \sa_count[12][63] , 
	\sa_count[12][62] , \sa_count[12][61] , \sa_count[12][60] , 
	\sa_count[12][59] , \sa_count[12][58] , \sa_count[12][57] , 
	\sa_count[12][56] , \sa_count[12][55] , \sa_count[12][54] , 
	\sa_count[12][53] , \sa_count[12][52] , \sa_count[12][51] , 
	\sa_count[12][50] , \sa_count[12][49] , \sa_count[12][48] , 
	\sa_count[12][47] , \sa_count[12][46] , \sa_count[12][45] , 
	\sa_count[12][44] , \sa_count[12][43] , \sa_count[12][42] , 
	\sa_count[12][41] , \sa_count[12][40] , \sa_count[12][39] , 
	\sa_count[12][38] , \sa_count[12][37] , \sa_count[12][36] , 
	\sa_count[12][35] , \sa_count[12][34] , \sa_count[12][33] , 
	\sa_count[12][32] , \sa_count[12][31] , \sa_count[12][30] , 
	\sa_count[12][29] , \sa_count[12][28] , \sa_count[12][27] , 
	\sa_count[12][26] , \sa_count[12][25] , \sa_count[12][24] , 
	\sa_count[12][23] , \sa_count[12][22] , \sa_count[12][21] , 
	\sa_count[12][20] , \sa_count[12][19] , \sa_count[12][18] , 
	\sa_count[12][17] , \sa_count[12][16] , \sa_count[12][15] , 
	\sa_count[12][14] , \sa_count[12][13] , \sa_count[12][12] , 
	\sa_count[12][11] , \sa_count[12][10] , \sa_count[12][9] , 
	\sa_count[12][8] , \sa_count[12][7] , \sa_count[12][6] , 
	\sa_count[12][5] , \sa_count[12][4] , \sa_count[12][3] , 
	\sa_count[12][2] , \sa_count[12][1] , \sa_count[12][0] , 
	\sa_count[11][63] , \sa_count[11][62] , \sa_count[11][61] , 
	\sa_count[11][60] , \sa_count[11][59] , \sa_count[11][58] , 
	\sa_count[11][57] , \sa_count[11][56] , \sa_count[11][55] , 
	\sa_count[11][54] , \sa_count[11][53] , \sa_count[11][52] , 
	\sa_count[11][51] , \sa_count[11][50] , \sa_count[11][49] , 
	\sa_count[11][48] , \sa_count[11][47] , \sa_count[11][46] , 
	\sa_count[11][45] , \sa_count[11][44] , \sa_count[11][43] , 
	\sa_count[11][42] , \sa_count[11][41] , \sa_count[11][40] , 
	\sa_count[11][39] , \sa_count[11][38] , \sa_count[11][37] , 
	\sa_count[11][36] , \sa_count[11][35] , \sa_count[11][34] , 
	\sa_count[11][33] , \sa_count[11][32] , \sa_count[11][31] , 
	\sa_count[11][30] , \sa_count[11][29] , \sa_count[11][28] , 
	\sa_count[11][27] , \sa_count[11][26] , \sa_count[11][25] , 
	\sa_count[11][24] , \sa_count[11][23] , \sa_count[11][22] , 
	\sa_count[11][21] , \sa_count[11][20] , \sa_count[11][19] , 
	\sa_count[11][18] , \sa_count[11][17] , \sa_count[11][16] , 
	\sa_count[11][15] , \sa_count[11][14] , \sa_count[11][13] , 
	\sa_count[11][12] , \sa_count[11][11] , \sa_count[11][10] , 
	\sa_count[11][9] , \sa_count[11][8] , \sa_count[11][7] , 
	\sa_count[11][6] , \sa_count[11][5] , \sa_count[11][4] , 
	\sa_count[11][3] , \sa_count[11][2] , \sa_count[11][1] , 
	\sa_count[11][0] , \sa_count[10][63] , \sa_count[10][62] , 
	\sa_count[10][61] , \sa_count[10][60] , \sa_count[10][59] , 
	\sa_count[10][58] , \sa_count[10][57] , \sa_count[10][56] , 
	\sa_count[10][55] , \sa_count[10][54] , \sa_count[10][53] , 
	\sa_count[10][52] , \sa_count[10][51] , \sa_count[10][50] , 
	\sa_count[10][49] , \sa_count[10][48] , \sa_count[10][47] , 
	\sa_count[10][46] , \sa_count[10][45] , \sa_count[10][44] , 
	\sa_count[10][43] , \sa_count[10][42] , \sa_count[10][41] , 
	\sa_count[10][40] , \sa_count[10][39] , \sa_count[10][38] , 
	\sa_count[10][37] , \sa_count[10][36] , \sa_count[10][35] , 
	\sa_count[10][34] , \sa_count[10][33] , \sa_count[10][32] , 
	\sa_count[10][31] , \sa_count[10][30] , \sa_count[10][29] , 
	\sa_count[10][28] , \sa_count[10][27] , \sa_count[10][26] , 
	\sa_count[10][25] , \sa_count[10][24] , \sa_count[10][23] , 
	\sa_count[10][22] , \sa_count[10][21] , \sa_count[10][20] , 
	\sa_count[10][19] , \sa_count[10][18] , \sa_count[10][17] , 
	\sa_count[10][16] , \sa_count[10][15] , \sa_count[10][14] , 
	\sa_count[10][13] , \sa_count[10][12] , \sa_count[10][11] , 
	\sa_count[10][10] , \sa_count[10][9] , \sa_count[10][8] , 
	\sa_count[10][7] , \sa_count[10][6] , \sa_count[10][5] , 
	\sa_count[10][4] , \sa_count[10][3] , \sa_count[10][2] , 
	\sa_count[10][1] , \sa_count[10][0] , \sa_count[9][63] , 
	\sa_count[9][62] , \sa_count[9][61] , \sa_count[9][60] , 
	\sa_count[9][59] , \sa_count[9][58] , \sa_count[9][57] , 
	\sa_count[9][56] , \sa_count[9][55] , \sa_count[9][54] , 
	\sa_count[9][53] , \sa_count[9][52] , \sa_count[9][51] , 
	\sa_count[9][50] , \sa_count[9][49] , \sa_count[9][48] , 
	\sa_count[9][47] , \sa_count[9][46] , \sa_count[9][45] , 
	\sa_count[9][44] , \sa_count[9][43] , \sa_count[9][42] , 
	\sa_count[9][41] , \sa_count[9][40] , \sa_count[9][39] , 
	\sa_count[9][38] , \sa_count[9][37] , \sa_count[9][36] , 
	\sa_count[9][35] , \sa_count[9][34] , \sa_count[9][33] , 
	\sa_count[9][32] , \sa_count[9][31] , \sa_count[9][30] , 
	\sa_count[9][29] , \sa_count[9][28] , \sa_count[9][27] , 
	\sa_count[9][26] , \sa_count[9][25] , \sa_count[9][24] , 
	\sa_count[9][23] , \sa_count[9][22] , \sa_count[9][21] , 
	\sa_count[9][20] , \sa_count[9][19] , \sa_count[9][18] , 
	\sa_count[9][17] , \sa_count[9][16] , \sa_count[9][15] , 
	\sa_count[9][14] , \sa_count[9][13] , \sa_count[9][12] , 
	\sa_count[9][11] , \sa_count[9][10] , \sa_count[9][9] , 
	\sa_count[9][8] , \sa_count[9][7] , \sa_count[9][6] , 
	\sa_count[9][5] , \sa_count[9][4] , \sa_count[9][3] , 
	\sa_count[9][2] , \sa_count[9][1] , \sa_count[9][0] , 
	\sa_count[8][63] , \sa_count[8][62] , \sa_count[8][61] , 
	\sa_count[8][60] , \sa_count[8][59] , \sa_count[8][58] , 
	\sa_count[8][57] , \sa_count[8][56] , \sa_count[8][55] , 
	\sa_count[8][54] , \sa_count[8][53] , \sa_count[8][52] , 
	\sa_count[8][51] , \sa_count[8][50] , \sa_count[8][49] , 
	\sa_count[8][48] , \sa_count[8][47] , \sa_count[8][46] , 
	\sa_count[8][45] , \sa_count[8][44] , \sa_count[8][43] , 
	\sa_count[8][42] , \sa_count[8][41] , \sa_count[8][40] , 
	\sa_count[8][39] , \sa_count[8][38] , \sa_count[8][37] , 
	\sa_count[8][36] , \sa_count[8][35] , \sa_count[8][34] , 
	\sa_count[8][33] , \sa_count[8][32] , \sa_count[8][31] , 
	\sa_count[8][30] , \sa_count[8][29] , \sa_count[8][28] , 
	\sa_count[8][27] , \sa_count[8][26] , \sa_count[8][25] , 
	\sa_count[8][24] , \sa_count[8][23] , \sa_count[8][22] , 
	\sa_count[8][21] , \sa_count[8][20] , \sa_count[8][19] , 
	\sa_count[8][18] , \sa_count[8][17] , \sa_count[8][16] , 
	\sa_count[8][15] , \sa_count[8][14] , \sa_count[8][13] , 
	\sa_count[8][12] , \sa_count[8][11] , \sa_count[8][10] , 
	\sa_count[8][9] , \sa_count[8][8] , \sa_count[8][7] , 
	\sa_count[8][6] , \sa_count[8][5] , \sa_count[8][4] , 
	\sa_count[8][3] , \sa_count[8][2] , \sa_count[8][1] , 
	\sa_count[8][0] , \sa_count[7][63] , \sa_count[7][62] , 
	\sa_count[7][61] , \sa_count[7][60] , \sa_count[7][59] , 
	\sa_count[7][58] , \sa_count[7][57] , \sa_count[7][56] , 
	\sa_count[7][55] , \sa_count[7][54] , \sa_count[7][53] , 
	\sa_count[7][52] , \sa_count[7][51] , \sa_count[7][50] , 
	\sa_count[7][49] , \sa_count[7][48] , \sa_count[7][47] , 
	\sa_count[7][46] , \sa_count[7][45] , \sa_count[7][44] , 
	\sa_count[7][43] , \sa_count[7][42] , \sa_count[7][41] , 
	\sa_count[7][40] , \sa_count[7][39] , \sa_count[7][38] , 
	\sa_count[7][37] , \sa_count[7][36] , \sa_count[7][35] , 
	\sa_count[7][34] , \sa_count[7][33] , \sa_count[7][32] , 
	\sa_count[7][31] , \sa_count[7][30] , \sa_count[7][29] , 
	\sa_count[7][28] , \sa_count[7][27] , \sa_count[7][26] , 
	\sa_count[7][25] , \sa_count[7][24] , \sa_count[7][23] , 
	\sa_count[7][22] , \sa_count[7][21] , \sa_count[7][20] , 
	\sa_count[7][19] , \sa_count[7][18] , \sa_count[7][17] , 
	\sa_count[7][16] , \sa_count[7][15] , \sa_count[7][14] , 
	\sa_count[7][13] , \sa_count[7][12] , \sa_count[7][11] , 
	\sa_count[7][10] , \sa_count[7][9] , \sa_count[7][8] , 
	\sa_count[7][7] , \sa_count[7][6] , \sa_count[7][5] , 
	\sa_count[7][4] , \sa_count[7][3] , \sa_count[7][2] , 
	\sa_count[7][1] , \sa_count[7][0] , \sa_count[6][63] , 
	\sa_count[6][62] , \sa_count[6][61] , \sa_count[6][60] , 
	\sa_count[6][59] , \sa_count[6][58] , \sa_count[6][57] , 
	\sa_count[6][56] , \sa_count[6][55] , \sa_count[6][54] , 
	\sa_count[6][53] , \sa_count[6][52] , \sa_count[6][51] , 
	\sa_count[6][50] , \sa_count[6][49] , \sa_count[6][48] , 
	\sa_count[6][47] , \sa_count[6][46] , \sa_count[6][45] , 
	\sa_count[6][44] , \sa_count[6][43] , \sa_count[6][42] , 
	\sa_count[6][41] , \sa_count[6][40] , \sa_count[6][39] , 
	\sa_count[6][38] , \sa_count[6][37] , \sa_count[6][36] , 
	\sa_count[6][35] , \sa_count[6][34] , \sa_count[6][33] , 
	\sa_count[6][32] , \sa_count[6][31] , \sa_count[6][30] , 
	\sa_count[6][29] , \sa_count[6][28] , \sa_count[6][27] , 
	\sa_count[6][26] , \sa_count[6][25] , \sa_count[6][24] , 
	\sa_count[6][23] , \sa_count[6][22] , \sa_count[6][21] , 
	\sa_count[6][20] , \sa_count[6][19] , \sa_count[6][18] , 
	\sa_count[6][17] , \sa_count[6][16] , \sa_count[6][15] , 
	\sa_count[6][14] , \sa_count[6][13] , \sa_count[6][12] , 
	\sa_count[6][11] , \sa_count[6][10] , \sa_count[6][9] , 
	\sa_count[6][8] , \sa_count[6][7] , \sa_count[6][6] , 
	\sa_count[6][5] , \sa_count[6][4] , \sa_count[6][3] , 
	\sa_count[6][2] , \sa_count[6][1] , \sa_count[6][0] , 
	\sa_count[5][63] , \sa_count[5][62] , \sa_count[5][61] , 
	\sa_count[5][60] , \sa_count[5][59] , \sa_count[5][58] , 
	\sa_count[5][57] , \sa_count[5][56] , \sa_count[5][55] , 
	\sa_count[5][54] , \sa_count[5][53] , \sa_count[5][52] , 
	\sa_count[5][51] , \sa_count[5][50] , \sa_count[5][49] , 
	\sa_count[5][48] , \sa_count[5][47] , \sa_count[5][46] , 
	\sa_count[5][45] , \sa_count[5][44] , \sa_count[5][43] , 
	\sa_count[5][42] , \sa_count[5][41] , \sa_count[5][40] , 
	\sa_count[5][39] , \sa_count[5][38] , \sa_count[5][37] , 
	\sa_count[5][36] , \sa_count[5][35] , \sa_count[5][34] , 
	\sa_count[5][33] , \sa_count[5][32] , \sa_count[5][31] , 
	\sa_count[5][30] , \sa_count[5][29] , \sa_count[5][28] , 
	\sa_count[5][27] , \sa_count[5][26] , \sa_count[5][25] , 
	\sa_count[5][24] , \sa_count[5][23] , \sa_count[5][22] , 
	\sa_count[5][21] , \sa_count[5][20] , \sa_count[5][19] , 
	\sa_count[5][18] , \sa_count[5][17] , \sa_count[5][16] , 
	\sa_count[5][15] , \sa_count[5][14] , \sa_count[5][13] , 
	\sa_count[5][12] , \sa_count[5][11] , \sa_count[5][10] , 
	\sa_count[5][9] , \sa_count[5][8] , \sa_count[5][7] , 
	\sa_count[5][6] , \sa_count[5][5] , \sa_count[5][4] , 
	\sa_count[5][3] , \sa_count[5][2] , \sa_count[5][1] , 
	\sa_count[5][0] , \sa_count[4][63] , \sa_count[4][62] , 
	\sa_count[4][61] , \sa_count[4][60] , \sa_count[4][59] , 
	\sa_count[4][58] , \sa_count[4][57] , \sa_count[4][56] , 
	\sa_count[4][55] , \sa_count[4][54] , \sa_count[4][53] , 
	\sa_count[4][52] , \sa_count[4][51] , \sa_count[4][50] , 
	\sa_count[4][49] , \sa_count[4][48] , \sa_count[4][47] , 
	\sa_count[4][46] , \sa_count[4][45] , \sa_count[4][44] , 
	\sa_count[4][43] , \sa_count[4][42] , \sa_count[4][41] , 
	\sa_count[4][40] , \sa_count[4][39] , \sa_count[4][38] , 
	\sa_count[4][37] , \sa_count[4][36] , \sa_count[4][35] , 
	\sa_count[4][34] , \sa_count[4][33] , \sa_count[4][32] , 
	\sa_count[4][31] , \sa_count[4][30] , \sa_count[4][29] , 
	\sa_count[4][28] , \sa_count[4][27] , \sa_count[4][26] , 
	\sa_count[4][25] , \sa_count[4][24] , \sa_count[4][23] , 
	\sa_count[4][22] , \sa_count[4][21] , \sa_count[4][20] , 
	\sa_count[4][19] , \sa_count[4][18] , \sa_count[4][17] , 
	\sa_count[4][16] , \sa_count[4][15] , \sa_count[4][14] , 
	\sa_count[4][13] , \sa_count[4][12] , \sa_count[4][11] , 
	\sa_count[4][10] , \sa_count[4][9] , \sa_count[4][8] , 
	\sa_count[4][7] , \sa_count[4][6] , \sa_count[4][5] , 
	\sa_count[4][4] , \sa_count[4][3] , \sa_count[4][2] , 
	\sa_count[4][1] , \sa_count[4][0] , \sa_count[3][63] , 
	\sa_count[3][62] , \sa_count[3][61] , \sa_count[3][60] , 
	\sa_count[3][59] , \sa_count[3][58] , \sa_count[3][57] , 
	\sa_count[3][56] , \sa_count[3][55] , \sa_count[3][54] , 
	\sa_count[3][53] , \sa_count[3][52] , \sa_count[3][51] , 
	\sa_count[3][50] , \sa_count[3][49] , \sa_count[3][48] , 
	\sa_count[3][47] , \sa_count[3][46] , \sa_count[3][45] , 
	\sa_count[3][44] , \sa_count[3][43] , \sa_count[3][42] , 
	\sa_count[3][41] , \sa_count[3][40] , \sa_count[3][39] , 
	\sa_count[3][38] , \sa_count[3][37] , \sa_count[3][36] , 
	\sa_count[3][35] , \sa_count[3][34] , \sa_count[3][33] , 
	\sa_count[3][32] , \sa_count[3][31] , \sa_count[3][30] , 
	\sa_count[3][29] , \sa_count[3][28] , \sa_count[3][27] , 
	\sa_count[3][26] , \sa_count[3][25] , \sa_count[3][24] , 
	\sa_count[3][23] , \sa_count[3][22] , \sa_count[3][21] , 
	\sa_count[3][20] , \sa_count[3][19] , \sa_count[3][18] , 
	\sa_count[3][17] , \sa_count[3][16] , \sa_count[3][15] , 
	\sa_count[3][14] , \sa_count[3][13] , \sa_count[3][12] , 
	\sa_count[3][11] , \sa_count[3][10] , \sa_count[3][9] , 
	\sa_count[3][8] , \sa_count[3][7] , \sa_count[3][6] , 
	\sa_count[3][5] , \sa_count[3][4] , \sa_count[3][3] , 
	\sa_count[3][2] , \sa_count[3][1] , \sa_count[3][0] , 
	\sa_count[2][63] , \sa_count[2][62] , \sa_count[2][61] , 
	\sa_count[2][60] , \sa_count[2][59] , \sa_count[2][58] , 
	\sa_count[2][57] , \sa_count[2][56] , \sa_count[2][55] , 
	\sa_count[2][54] , \sa_count[2][53] , \sa_count[2][52] , 
	\sa_count[2][51] , \sa_count[2][50] , \sa_count[2][49] , 
	\sa_count[2][48] , \sa_count[2][47] , \sa_count[2][46] , 
	\sa_count[2][45] , \sa_count[2][44] , \sa_count[2][43] , 
	\sa_count[2][42] , \sa_count[2][41] , \sa_count[2][40] , 
	\sa_count[2][39] , \sa_count[2][38] , \sa_count[2][37] , 
	\sa_count[2][36] , \sa_count[2][35] , \sa_count[2][34] , 
	\sa_count[2][33] , \sa_count[2][32] , \sa_count[2][31] , 
	\sa_count[2][30] , \sa_count[2][29] , \sa_count[2][28] , 
	\sa_count[2][27] , \sa_count[2][26] , \sa_count[2][25] , 
	\sa_count[2][24] , \sa_count[2][23] , \sa_count[2][22] , 
	\sa_count[2][21] , \sa_count[2][20] , \sa_count[2][19] , 
	\sa_count[2][18] , \sa_count[2][17] , \sa_count[2][16] , 
	\sa_count[2][15] , \sa_count[2][14] , \sa_count[2][13] , 
	\sa_count[2][12] , \sa_count[2][11] , \sa_count[2][10] , 
	\sa_count[2][9] , \sa_count[2][8] , \sa_count[2][7] , 
	\sa_count[2][6] , \sa_count[2][5] , \sa_count[2][4] , 
	\sa_count[2][3] , \sa_count[2][2] , \sa_count[2][1] , 
	\sa_count[2][0] , \sa_count[1][63] , \sa_count[1][62] , 
	\sa_count[1][61] , \sa_count[1][60] , \sa_count[1][59] , 
	\sa_count[1][58] , \sa_count[1][57] , \sa_count[1][56] , 
	\sa_count[1][55] , \sa_count[1][54] , \sa_count[1][53] , 
	\sa_count[1][52] , \sa_count[1][51] , \sa_count[1][50] , 
	\sa_count[1][49] , \sa_count[1][48] , \sa_count[1][47] , 
	\sa_count[1][46] , \sa_count[1][45] , \sa_count[1][44] , 
	\sa_count[1][43] , \sa_count[1][42] , \sa_count[1][41] , 
	\sa_count[1][40] , \sa_count[1][39] , \sa_count[1][38] , 
	\sa_count[1][37] , \sa_count[1][36] , \sa_count[1][35] , 
	\sa_count[1][34] , \sa_count[1][33] , \sa_count[1][32] , 
	\sa_count[1][31] , \sa_count[1][30] , \sa_count[1][29] , 
	\sa_count[1][28] , \sa_count[1][27] , \sa_count[1][26] , 
	\sa_count[1][25] , \sa_count[1][24] , \sa_count[1][23] , 
	\sa_count[1][22] , \sa_count[1][21] , \sa_count[1][20] , 
	\sa_count[1][19] , \sa_count[1][18] , \sa_count[1][17] , 
	\sa_count[1][16] , \sa_count[1][15] , \sa_count[1][14] , 
	\sa_count[1][13] , \sa_count[1][12] , \sa_count[1][11] , 
	\sa_count[1][10] , \sa_count[1][9] , \sa_count[1][8] , 
	\sa_count[1][7] , \sa_count[1][6] , \sa_count[1][5] , 
	\sa_count[1][4] , \sa_count[1][3] , \sa_count[1][2] , 
	\sa_count[1][1] , \sa_count[1][0] , \sa_count[0][63] , 
	\sa_count[0][62] , \sa_count[0][61] , \sa_count[0][60] , 
	\sa_count[0][59] , \sa_count[0][58] , \sa_count[0][57] , 
	\sa_count[0][56] , \sa_count[0][55] , \sa_count[0][54] , 
	\sa_count[0][53] , \sa_count[0][52] , \sa_count[0][51] , 
	\sa_count[0][50] , \sa_count[0][49] , \sa_count[0][48] , 
	\sa_count[0][47] , \sa_count[0][46] , \sa_count[0][45] , 
	\sa_count[0][44] , \sa_count[0][43] , \sa_count[0][42] , 
	\sa_count[0][41] , \sa_count[0][40] , \sa_count[0][39] , 
	\sa_count[0][38] , \sa_count[0][37] , \sa_count[0][36] , 
	\sa_count[0][35] , \sa_count[0][34] , \sa_count[0][33] , 
	\sa_count[0][32] , \sa_count[0][31] , \sa_count[0][30] , 
	\sa_count[0][29] , \sa_count[0][28] , \sa_count[0][27] , 
	\sa_count[0][26] , \sa_count[0][25] , \sa_count[0][24] , 
	\sa_count[0][23] , \sa_count[0][22] , \sa_count[0][21] , 
	\sa_count[0][20] , \sa_count[0][19] , \sa_count[0][18] , 
	\sa_count[0][17] , \sa_count[0][16] , \sa_count[0][15] , 
	\sa_count[0][14] , \sa_count[0][13] , \sa_count[0][12] , 
	\sa_count[0][11] , \sa_count[0][10] , \sa_count[0][9] , 
	\sa_count[0][8] , \sa_count[0][7] , \sa_count[0][6] , 
	\sa_count[0][5] , \sa_count[0][4] , \sa_count[0][3] , 
	\sa_count[0][2] , \sa_count[0][1] , \sa_count[0][0] }), 
	.debug_kme_ib_tready( debug_kme_ib_tready));
nx_rbus_apb u_nx_rbus_apb ( .rbus_addr_o( _zy_simnet_rbus_ring_i_26_w$[0:15]), 
	.rbus_wr_strb_o( _zy_simnet_rbus_ring_i_27_w$), .rbus_wr_data_o( 
	_zy_simnet_rbus_ring_i_28_w$[0:31]), .rbus_rd_strb_o( 
	_zy_simnet_rbus_ring_i_29_w$), .apb_prdata( apb_prdata[31:0]), 
	.apb_pready( apb_pready), .apb_pslverr( apb_pslverr), .clk( clk), 
	.rst_n( rst_sync_n), .rbus_rd_data_i( 
	_zy_simnet_rbus_ring_o_30_w$[0:31]), .rbus_ack_i( 
	_zy_simnet_rbus_ring_o_31_w$), .rbus_err_ack_i( 
	_zy_simnet_rbus_ring_o_32_w$), .rbus_wr_strb_i( 
	_zy_simnet_rbus_ring_o_33_w$), .rbus_rd_strb_i( 
	_zy_simnet_rbus_ring_o_34_w$), .apb_paddr( apb_paddr[15:0]), 
	.apb_psel( apb_psel), .apb_penable( apb_penable), .apb_pwrite( 
	apb_pwrite), .apb_pwdata( apb_pwdata[31:0]));
cr_kme_core u_cr_kme_core ( .kme_ib_out( _zy_simnet_kme_ib_out_0_w$), 
	.kme_cceip0_ob_out( _zy_simnet_kme_cceip0_ob_out_pre_1_w$[0:82]), 
	.kme_cceip1_ob_out( _zy_simnet_kme_cceip1_ob_out_pre_2_w$[0:82]), 
	.kme_cceip2_ob_out( _zy_simnet_kme_cceip2_ob_out_pre_3_w$[0:82]), 
	.kme_cceip3_ob_out( _zy_simnet_kme_cceip3_ob_out_pre_4_w$[0:82]), 
	.kme_cddip0_ob_out( _zy_simnet_kme_cddip0_ob_out_pre_5_w$[0:82]), 
	.kme_cddip1_ob_out( _zy_simnet_kme_cddip1_ob_out_pre_6_w$[0:82]), 
	.kme_cddip2_ob_out( _zy_simnet_kme_cddip2_ob_out_pre_7_w$[0:82]), 
	.kme_cddip3_ob_out( _zy_simnet_kme_cddip3_ob_out_pre_8_w$[0:82]), 
	.ckv_rd( ckv_rd), .ckv_addr( ckv_addr[14:0]), .kim_rd( kim_rd), 
	.kim_addr( kim_addr[13:0]), .cceip_encrypt_bimc_osync( 
	cceip_encrypt_bimc_osync), .cceip_encrypt_bimc_odat( 
	cceip_encrypt_bimc_odat), .cceip_encrypt_mbe( cceip_encrypt_mbe), 
	.cceip_validate_bimc_osync( cceip_validate_bimc_osync), 
	.cceip_validate_bimc_odat( cceip_validate_bimc_odat), 
	.cceip_validate_mbe( cceip_validate_mbe), 
	.cddip_decrypt_bimc_osync( cddip_decrypt_bimc_osync), 
	.cddip_decrypt_bimc_odat( cddip_decrypt_bimc_odat), 
	.cddip_decrypt_mbe( cddip_decrypt_mbe), .axi_bimc_osync( 
	axi_bimc_osync), .axi_bimc_odat( axi_bimc_odat), .axi_mbe( axi_mbe), 
	.seed0_invalidate( seed0_invalidate), .seed1_invalidate( 
	seed1_invalidate), .set_txc_bp_int( set_txc_bp_int), 
	.set_gcm_tag_fail_int( set_gcm_tag_fail_int), 
	.set_key_tlv_miscmp_int( set_key_tlv_miscmp_int), 
	.set_tlv_bip2_error_int( set_tlv_bip2_error_int), 
	.set_rsm_is_backpressuring( set_rsm_is_backpressuring[7:0]), 
	.idle_components( _zy_simnet_idle_components_9_w$[0:31]), 
	.sa_snapshot( { \sa_snapshot[31][63] , \sa_snapshot[31][62] , 
	\sa_snapshot[31][61] , \sa_snapshot[31][60] , \sa_snapshot[31][59] , 
	\sa_snapshot[31][58] , \sa_snapshot[31][57] , \sa_snapshot[31][56] , 
	\sa_snapshot[31][55] , \sa_snapshot[31][54] , \sa_snapshot[31][53] , 
	\sa_snapshot[31][52] , \sa_snapshot[31][51] , \sa_snapshot[31][50] , 
	\sa_snapshot[31][49] , \sa_snapshot[31][48] , \sa_snapshot[31][47] , 
	\sa_snapshot[31][46] , \sa_snapshot[31][45] , \sa_snapshot[31][44] , 
	\sa_snapshot[31][43] , \sa_snapshot[31][42] , \sa_snapshot[31][41] , 
	\sa_snapshot[31][40] , \sa_snapshot[31][39] , \sa_snapshot[31][38] , 
	\sa_snapshot[31][37] , \sa_snapshot[31][36] , \sa_snapshot[31][35] , 
	\sa_snapshot[31][34] , \sa_snapshot[31][33] , \sa_snapshot[31][32] , 
	\sa_snapshot[31][31] , \sa_snapshot[31][30] , \sa_snapshot[31][29] , 
	\sa_snapshot[31][28] , \sa_snapshot[31][27] , \sa_snapshot[31][26] , 
	\sa_snapshot[31][25] , \sa_snapshot[31][24] , \sa_snapshot[31][23] , 
	\sa_snapshot[31][22] , \sa_snapshot[31][21] , \sa_snapshot[31][20] , 
	\sa_snapshot[31][19] , \sa_snapshot[31][18] , \sa_snapshot[31][17] , 
	\sa_snapshot[31][16] , \sa_snapshot[31][15] , \sa_snapshot[31][14] , 
	\sa_snapshot[31][13] , \sa_snapshot[31][12] , \sa_snapshot[31][11] , 
	\sa_snapshot[31][10] , \sa_snapshot[31][9] , \sa_snapshot[31][8] , 
	\sa_snapshot[31][7] , \sa_snapshot[31][6] , \sa_snapshot[31][5] , 
	\sa_snapshot[31][4] , \sa_snapshot[31][3] , \sa_snapshot[31][2] , 
	\sa_snapshot[31][1] , \sa_snapshot[31][0] , \sa_snapshot[30][63] , 
	\sa_snapshot[30][62] , \sa_snapshot[30][61] , \sa_snapshot[30][60] , 
	\sa_snapshot[30][59] , \sa_snapshot[30][58] , \sa_snapshot[30][57] , 
	\sa_snapshot[30][56] , \sa_snapshot[30][55] , \sa_snapshot[30][54] , 
	\sa_snapshot[30][53] , \sa_snapshot[30][52] , \sa_snapshot[30][51] , 
	\sa_snapshot[30][50] , \sa_snapshot[30][49] , \sa_snapshot[30][48] , 
	\sa_snapshot[30][47] , \sa_snapshot[30][46] , \sa_snapshot[30][45] , 
	\sa_snapshot[30][44] , \sa_snapshot[30][43] , \sa_snapshot[30][42] , 
	\sa_snapshot[30][41] , \sa_snapshot[30][40] , \sa_snapshot[30][39] , 
	\sa_snapshot[30][38] , \sa_snapshot[30][37] , \sa_snapshot[30][36] , 
	\sa_snapshot[30][35] , \sa_snapshot[30][34] , \sa_snapshot[30][33] , 
	\sa_snapshot[30][32] , \sa_snapshot[30][31] , \sa_snapshot[30][30] , 
	\sa_snapshot[30][29] , \sa_snapshot[30][28] , \sa_snapshot[30][27] , 
	\sa_snapshot[30][26] , \sa_snapshot[30][25] , \sa_snapshot[30][24] , 
	\sa_snapshot[30][23] , \sa_snapshot[30][22] , \sa_snapshot[30][21] , 
	\sa_snapshot[30][20] , \sa_snapshot[30][19] , \sa_snapshot[30][18] , 
	\sa_snapshot[30][17] , \sa_snapshot[30][16] , \sa_snapshot[30][15] , 
	\sa_snapshot[30][14] , \sa_snapshot[30][13] , \sa_snapshot[30][12] , 
	\sa_snapshot[30][11] , \sa_snapshot[30][10] , \sa_snapshot[30][9] , 
	\sa_snapshot[30][8] , \sa_snapshot[30][7] , \sa_snapshot[30][6] , 
	\sa_snapshot[30][5] , \sa_snapshot[30][4] , \sa_snapshot[30][3] , 
	\sa_snapshot[30][2] , \sa_snapshot[30][1] , \sa_snapshot[30][0] , 
	\sa_snapshot[29][63] , \sa_snapshot[29][62] , \sa_snapshot[29][61] , 
	\sa_snapshot[29][60] , \sa_snapshot[29][59] , \sa_snapshot[29][58] , 
	\sa_snapshot[29][57] , \sa_snapshot[29][56] , \sa_snapshot[29][55] , 
	\sa_snapshot[29][54] , \sa_snapshot[29][53] , \sa_snapshot[29][52] , 
	\sa_snapshot[29][51] , \sa_snapshot[29][50] , \sa_snapshot[29][49] , 
	\sa_snapshot[29][48] , \sa_snapshot[29][47] , \sa_snapshot[29][46] , 
	\sa_snapshot[29][45] , \sa_snapshot[29][44] , \sa_snapshot[29][43] , 
	\sa_snapshot[29][42] , \sa_snapshot[29][41] , \sa_snapshot[29][40] , 
	\sa_snapshot[29][39] , \sa_snapshot[29][38] , \sa_snapshot[29][37] , 
	\sa_snapshot[29][36] , \sa_snapshot[29][35] , \sa_snapshot[29][34] , 
	\sa_snapshot[29][33] , \sa_snapshot[29][32] , \sa_snapshot[29][31] , 
	\sa_snapshot[29][30] , \sa_snapshot[29][29] , \sa_snapshot[29][28] , 
	\sa_snapshot[29][27] , \sa_snapshot[29][26] , \sa_snapshot[29][25] , 
	\sa_snapshot[29][24] , \sa_snapshot[29][23] , \sa_snapshot[29][22] , 
	\sa_snapshot[29][21] , \sa_snapshot[29][20] , \sa_snapshot[29][19] , 
	\sa_snapshot[29][18] , \sa_snapshot[29][17] , \sa_snapshot[29][16] , 
	\sa_snapshot[29][15] , \sa_snapshot[29][14] , \sa_snapshot[29][13] , 
	\sa_snapshot[29][12] , \sa_snapshot[29][11] , \sa_snapshot[29][10] , 
	\sa_snapshot[29][9] , \sa_snapshot[29][8] , \sa_snapshot[29][7] , 
	\sa_snapshot[29][6] , \sa_snapshot[29][5] , \sa_snapshot[29][4] , 
	\sa_snapshot[29][3] , \sa_snapshot[29][2] , \sa_snapshot[29][1] , 
	\sa_snapshot[29][0] , \sa_snapshot[28][63] , \sa_snapshot[28][62] , 
	\sa_snapshot[28][61] , \sa_snapshot[28][60] , \sa_snapshot[28][59] , 
	\sa_snapshot[28][58] , \sa_snapshot[28][57] , \sa_snapshot[28][56] , 
	\sa_snapshot[28][55] , \sa_snapshot[28][54] , \sa_snapshot[28][53] , 
	\sa_snapshot[28][52] , \sa_snapshot[28][51] , \sa_snapshot[28][50] , 
	\sa_snapshot[28][49] , \sa_snapshot[28][48] , \sa_snapshot[28][47] , 
	\sa_snapshot[28][46] , \sa_snapshot[28][45] , \sa_snapshot[28][44] , 
	\sa_snapshot[28][43] , \sa_snapshot[28][42] , \sa_snapshot[28][41] , 
	\sa_snapshot[28][40] , \sa_snapshot[28][39] , \sa_snapshot[28][38] , 
	\sa_snapshot[28][37] , \sa_snapshot[28][36] , \sa_snapshot[28][35] , 
	\sa_snapshot[28][34] , \sa_snapshot[28][33] , \sa_snapshot[28][32] , 
	\sa_snapshot[28][31] , \sa_snapshot[28][30] , \sa_snapshot[28][29] , 
	\sa_snapshot[28][28] , \sa_snapshot[28][27] , \sa_snapshot[28][26] , 
	\sa_snapshot[28][25] , \sa_snapshot[28][24] , \sa_snapshot[28][23] , 
	\sa_snapshot[28][22] , \sa_snapshot[28][21] , \sa_snapshot[28][20] , 
	\sa_snapshot[28][19] , \sa_snapshot[28][18] , \sa_snapshot[28][17] , 
	\sa_snapshot[28][16] , \sa_snapshot[28][15] , \sa_snapshot[28][14] , 
	\sa_snapshot[28][13] , \sa_snapshot[28][12] , \sa_snapshot[28][11] , 
	\sa_snapshot[28][10] , \sa_snapshot[28][9] , \sa_snapshot[28][8] , 
	\sa_snapshot[28][7] , \sa_snapshot[28][6] , \sa_snapshot[28][5] , 
	\sa_snapshot[28][4] , \sa_snapshot[28][3] , \sa_snapshot[28][2] , 
	\sa_snapshot[28][1] , \sa_snapshot[28][0] , \sa_snapshot[27][63] , 
	\sa_snapshot[27][62] , \sa_snapshot[27][61] , \sa_snapshot[27][60] , 
	\sa_snapshot[27][59] , \sa_snapshot[27][58] , \sa_snapshot[27][57] , 
	\sa_snapshot[27][56] , \sa_snapshot[27][55] , \sa_snapshot[27][54] , 
	\sa_snapshot[27][53] , \sa_snapshot[27][52] , \sa_snapshot[27][51] , 
	\sa_snapshot[27][50] , \sa_snapshot[27][49] , \sa_snapshot[27][48] , 
	\sa_snapshot[27][47] , \sa_snapshot[27][46] , \sa_snapshot[27][45] , 
	\sa_snapshot[27][44] , \sa_snapshot[27][43] , \sa_snapshot[27][42] , 
	\sa_snapshot[27][41] , \sa_snapshot[27][40] , \sa_snapshot[27][39] , 
	\sa_snapshot[27][38] , \sa_snapshot[27][37] , \sa_snapshot[27][36] , 
	\sa_snapshot[27][35] , \sa_snapshot[27][34] , \sa_snapshot[27][33] , 
	\sa_snapshot[27][32] , \sa_snapshot[27][31] , \sa_snapshot[27][30] , 
	\sa_snapshot[27][29] , \sa_snapshot[27][28] , \sa_snapshot[27][27] , 
	\sa_snapshot[27][26] , \sa_snapshot[27][25] , \sa_snapshot[27][24] , 
	\sa_snapshot[27][23] , \sa_snapshot[27][22] , \sa_snapshot[27][21] , 
	\sa_snapshot[27][20] , \sa_snapshot[27][19] , \sa_snapshot[27][18] , 
	\sa_snapshot[27][17] , \sa_snapshot[27][16] , \sa_snapshot[27][15] , 
	\sa_snapshot[27][14] , \sa_snapshot[27][13] , \sa_snapshot[27][12] , 
	\sa_snapshot[27][11] , \sa_snapshot[27][10] , \sa_snapshot[27][9] , 
	\sa_snapshot[27][8] , \sa_snapshot[27][7] , \sa_snapshot[27][6] , 
	\sa_snapshot[27][5] , \sa_snapshot[27][4] , \sa_snapshot[27][3] , 
	\sa_snapshot[27][2] , \sa_snapshot[27][1] , \sa_snapshot[27][0] , 
	\sa_snapshot[26][63] , \sa_snapshot[26][62] , \sa_snapshot[26][61] , 
	\sa_snapshot[26][60] , \sa_snapshot[26][59] , \sa_snapshot[26][58] , 
	\sa_snapshot[26][57] , \sa_snapshot[26][56] , \sa_snapshot[26][55] , 
	\sa_snapshot[26][54] , \sa_snapshot[26][53] , \sa_snapshot[26][52] , 
	\sa_snapshot[26][51] , \sa_snapshot[26][50] , \sa_snapshot[26][49] , 
	\sa_snapshot[26][48] , \sa_snapshot[26][47] , \sa_snapshot[26][46] , 
	\sa_snapshot[26][45] , \sa_snapshot[26][44] , \sa_snapshot[26][43] , 
	\sa_snapshot[26][42] , \sa_snapshot[26][41] , \sa_snapshot[26][40] , 
	\sa_snapshot[26][39] , \sa_snapshot[26][38] , \sa_snapshot[26][37] , 
	\sa_snapshot[26][36] , \sa_snapshot[26][35] , \sa_snapshot[26][34] , 
	\sa_snapshot[26][33] , \sa_snapshot[26][32] , \sa_snapshot[26][31] , 
	\sa_snapshot[26][30] , \sa_snapshot[26][29] , \sa_snapshot[26][28] , 
	\sa_snapshot[26][27] , \sa_snapshot[26][26] , \sa_snapshot[26][25] , 
	\sa_snapshot[26][24] , \sa_snapshot[26][23] , \sa_snapshot[26][22] , 
	\sa_snapshot[26][21] , \sa_snapshot[26][20] , \sa_snapshot[26][19] , 
	\sa_snapshot[26][18] , \sa_snapshot[26][17] , \sa_snapshot[26][16] , 
	\sa_snapshot[26][15] , \sa_snapshot[26][14] , \sa_snapshot[26][13] , 
	\sa_snapshot[26][12] , \sa_snapshot[26][11] , \sa_snapshot[26][10] , 
	\sa_snapshot[26][9] , \sa_snapshot[26][8] , \sa_snapshot[26][7] , 
	\sa_snapshot[26][6] , \sa_snapshot[26][5] , \sa_snapshot[26][4] , 
	\sa_snapshot[26][3] , \sa_snapshot[26][2] , \sa_snapshot[26][1] , 
	\sa_snapshot[26][0] , \sa_snapshot[25][63] , \sa_snapshot[25][62] , 
	\sa_snapshot[25][61] , \sa_snapshot[25][60] , \sa_snapshot[25][59] , 
	\sa_snapshot[25][58] , \sa_snapshot[25][57] , \sa_snapshot[25][56] , 
	\sa_snapshot[25][55] , \sa_snapshot[25][54] , \sa_snapshot[25][53] , 
	\sa_snapshot[25][52] , \sa_snapshot[25][51] , \sa_snapshot[25][50] , 
	\sa_snapshot[25][49] , \sa_snapshot[25][48] , \sa_snapshot[25][47] , 
	\sa_snapshot[25][46] , \sa_snapshot[25][45] , \sa_snapshot[25][44] , 
	\sa_snapshot[25][43] , \sa_snapshot[25][42] , \sa_snapshot[25][41] , 
	\sa_snapshot[25][40] , \sa_snapshot[25][39] , \sa_snapshot[25][38] , 
	\sa_snapshot[25][37] , \sa_snapshot[25][36] , \sa_snapshot[25][35] , 
	\sa_snapshot[25][34] , \sa_snapshot[25][33] , \sa_snapshot[25][32] , 
	\sa_snapshot[25][31] , \sa_snapshot[25][30] , \sa_snapshot[25][29] , 
	\sa_snapshot[25][28] , \sa_snapshot[25][27] , \sa_snapshot[25][26] , 
	\sa_snapshot[25][25] , \sa_snapshot[25][24] , \sa_snapshot[25][23] , 
	\sa_snapshot[25][22] , \sa_snapshot[25][21] , \sa_snapshot[25][20] , 
	\sa_snapshot[25][19] , \sa_snapshot[25][18] , \sa_snapshot[25][17] , 
	\sa_snapshot[25][16] , \sa_snapshot[25][15] , \sa_snapshot[25][14] , 
	\sa_snapshot[25][13] , \sa_snapshot[25][12] , \sa_snapshot[25][11] , 
	\sa_snapshot[25][10] , \sa_snapshot[25][9] , \sa_snapshot[25][8] , 
	\sa_snapshot[25][7] , \sa_snapshot[25][6] , \sa_snapshot[25][5] , 
	\sa_snapshot[25][4] , \sa_snapshot[25][3] , \sa_snapshot[25][2] , 
	\sa_snapshot[25][1] , \sa_snapshot[25][0] , \sa_snapshot[24][63] , 
	\sa_snapshot[24][62] , \sa_snapshot[24][61] , \sa_snapshot[24][60] , 
	\sa_snapshot[24][59] , \sa_snapshot[24][58] , \sa_snapshot[24][57] , 
	\sa_snapshot[24][56] , \sa_snapshot[24][55] , \sa_snapshot[24][54] , 
	\sa_snapshot[24][53] , \sa_snapshot[24][52] , \sa_snapshot[24][51] , 
	\sa_snapshot[24][50] , \sa_snapshot[24][49] , \sa_snapshot[24][48] , 
	\sa_snapshot[24][47] , \sa_snapshot[24][46] , \sa_snapshot[24][45] , 
	\sa_snapshot[24][44] , \sa_snapshot[24][43] , \sa_snapshot[24][42] , 
	\sa_snapshot[24][41] , \sa_snapshot[24][40] , \sa_snapshot[24][39] , 
	\sa_snapshot[24][38] , \sa_snapshot[24][37] , \sa_snapshot[24][36] , 
	\sa_snapshot[24][35] , \sa_snapshot[24][34] , \sa_snapshot[24][33] , 
	\sa_snapshot[24][32] , \sa_snapshot[24][31] , \sa_snapshot[24][30] , 
	\sa_snapshot[24][29] , \sa_snapshot[24][28] , \sa_snapshot[24][27] , 
	\sa_snapshot[24][26] , \sa_snapshot[24][25] , \sa_snapshot[24][24] , 
	\sa_snapshot[24][23] , \sa_snapshot[24][22] , \sa_snapshot[24][21] , 
	\sa_snapshot[24][20] , \sa_snapshot[24][19] , \sa_snapshot[24][18] , 
	\sa_snapshot[24][17] , \sa_snapshot[24][16] , \sa_snapshot[24][15] , 
	\sa_snapshot[24][14] , \sa_snapshot[24][13] , \sa_snapshot[24][12] , 
	\sa_snapshot[24][11] , \sa_snapshot[24][10] , \sa_snapshot[24][9] , 
	\sa_snapshot[24][8] , \sa_snapshot[24][7] , \sa_snapshot[24][6] , 
	\sa_snapshot[24][5] , \sa_snapshot[24][4] , \sa_snapshot[24][3] , 
	\sa_snapshot[24][2] , \sa_snapshot[24][1] , \sa_snapshot[24][0] , 
	\sa_snapshot[23][63] , \sa_snapshot[23][62] , \sa_snapshot[23][61] , 
	\sa_snapshot[23][60] , \sa_snapshot[23][59] , \sa_snapshot[23][58] , 
	\sa_snapshot[23][57] , \sa_snapshot[23][56] , \sa_snapshot[23][55] , 
	\sa_snapshot[23][54] , \sa_snapshot[23][53] , \sa_snapshot[23][52] , 
	\sa_snapshot[23][51] , \sa_snapshot[23][50] , \sa_snapshot[23][49] , 
	\sa_snapshot[23][48] , \sa_snapshot[23][47] , \sa_snapshot[23][46] , 
	\sa_snapshot[23][45] , \sa_snapshot[23][44] , \sa_snapshot[23][43] , 
	\sa_snapshot[23][42] , \sa_snapshot[23][41] , \sa_snapshot[23][40] , 
	\sa_snapshot[23][39] , \sa_snapshot[23][38] , \sa_snapshot[23][37] , 
	\sa_snapshot[23][36] , \sa_snapshot[23][35] , \sa_snapshot[23][34] , 
	\sa_snapshot[23][33] , \sa_snapshot[23][32] , \sa_snapshot[23][31] , 
	\sa_snapshot[23][30] , \sa_snapshot[23][29] , \sa_snapshot[23][28] , 
	\sa_snapshot[23][27] , \sa_snapshot[23][26] , \sa_snapshot[23][25] , 
	\sa_snapshot[23][24] , \sa_snapshot[23][23] , \sa_snapshot[23][22] , 
	\sa_snapshot[23][21] , \sa_snapshot[23][20] , \sa_snapshot[23][19] , 
	\sa_snapshot[23][18] , \sa_snapshot[23][17] , \sa_snapshot[23][16] , 
	\sa_snapshot[23][15] , \sa_snapshot[23][14] , \sa_snapshot[23][13] , 
	\sa_snapshot[23][12] , \sa_snapshot[23][11] , \sa_snapshot[23][10] , 
	\sa_snapshot[23][9] , \sa_snapshot[23][8] , \sa_snapshot[23][7] , 
	\sa_snapshot[23][6] , \sa_snapshot[23][5] , \sa_snapshot[23][4] , 
	\sa_snapshot[23][3] , \sa_snapshot[23][2] , \sa_snapshot[23][1] , 
	\sa_snapshot[23][0] , \sa_snapshot[22][63] , \sa_snapshot[22][62] , 
	\sa_snapshot[22][61] , \sa_snapshot[22][60] , \sa_snapshot[22][59] , 
	\sa_snapshot[22][58] , \sa_snapshot[22][57] , \sa_snapshot[22][56] , 
	\sa_snapshot[22][55] , \sa_snapshot[22][54] , \sa_snapshot[22][53] , 
	\sa_snapshot[22][52] , \sa_snapshot[22][51] , \sa_snapshot[22][50] , 
	\sa_snapshot[22][49] , \sa_snapshot[22][48] , \sa_snapshot[22][47] , 
	\sa_snapshot[22][46] , \sa_snapshot[22][45] , \sa_snapshot[22][44] , 
	\sa_snapshot[22][43] , \sa_snapshot[22][42] , \sa_snapshot[22][41] , 
	\sa_snapshot[22][40] , \sa_snapshot[22][39] , \sa_snapshot[22][38] , 
	\sa_snapshot[22][37] , \sa_snapshot[22][36] , \sa_snapshot[22][35] , 
	\sa_snapshot[22][34] , \sa_snapshot[22][33] , \sa_snapshot[22][32] , 
	\sa_snapshot[22][31] , \sa_snapshot[22][30] , \sa_snapshot[22][29] , 
	\sa_snapshot[22][28] , \sa_snapshot[22][27] , \sa_snapshot[22][26] , 
	\sa_snapshot[22][25] , \sa_snapshot[22][24] , \sa_snapshot[22][23] , 
	\sa_snapshot[22][22] , \sa_snapshot[22][21] , \sa_snapshot[22][20] , 
	\sa_snapshot[22][19] , \sa_snapshot[22][18] , \sa_snapshot[22][17] , 
	\sa_snapshot[22][16] , \sa_snapshot[22][15] , \sa_snapshot[22][14] , 
	\sa_snapshot[22][13] , \sa_snapshot[22][12] , \sa_snapshot[22][11] , 
	\sa_snapshot[22][10] , \sa_snapshot[22][9] , \sa_snapshot[22][8] , 
	\sa_snapshot[22][7] , \sa_snapshot[22][6] , \sa_snapshot[22][5] , 
	\sa_snapshot[22][4] , \sa_snapshot[22][3] , \sa_snapshot[22][2] , 
	\sa_snapshot[22][1] , \sa_snapshot[22][0] , \sa_snapshot[21][63] , 
	\sa_snapshot[21][62] , \sa_snapshot[21][61] , \sa_snapshot[21][60] , 
	\sa_snapshot[21][59] , \sa_snapshot[21][58] , \sa_snapshot[21][57] , 
	\sa_snapshot[21][56] , \sa_snapshot[21][55] , \sa_snapshot[21][54] , 
	\sa_snapshot[21][53] , \sa_snapshot[21][52] , \sa_snapshot[21][51] , 
	\sa_snapshot[21][50] , \sa_snapshot[21][49] , \sa_snapshot[21][48] , 
	\sa_snapshot[21][47] , \sa_snapshot[21][46] , \sa_snapshot[21][45] , 
	\sa_snapshot[21][44] , \sa_snapshot[21][43] , \sa_snapshot[21][42] , 
	\sa_snapshot[21][41] , \sa_snapshot[21][40] , \sa_snapshot[21][39] , 
	\sa_snapshot[21][38] , \sa_snapshot[21][37] , \sa_snapshot[21][36] , 
	\sa_snapshot[21][35] , \sa_snapshot[21][34] , \sa_snapshot[21][33] , 
	\sa_snapshot[21][32] , \sa_snapshot[21][31] , \sa_snapshot[21][30] , 
	\sa_snapshot[21][29] , \sa_snapshot[21][28] , \sa_snapshot[21][27] , 
	\sa_snapshot[21][26] , \sa_snapshot[21][25] , \sa_snapshot[21][24] , 
	\sa_snapshot[21][23] , \sa_snapshot[21][22] , \sa_snapshot[21][21] , 
	\sa_snapshot[21][20] , \sa_snapshot[21][19] , \sa_snapshot[21][18] , 
	\sa_snapshot[21][17] , \sa_snapshot[21][16] , \sa_snapshot[21][15] , 
	\sa_snapshot[21][14] , \sa_snapshot[21][13] , \sa_snapshot[21][12] , 
	\sa_snapshot[21][11] , \sa_snapshot[21][10] , \sa_snapshot[21][9] , 
	\sa_snapshot[21][8] , \sa_snapshot[21][7] , \sa_snapshot[21][6] , 
	\sa_snapshot[21][5] , \sa_snapshot[21][4] , \sa_snapshot[21][3] , 
	\sa_snapshot[21][2] , \sa_snapshot[21][1] , \sa_snapshot[21][0] , 
	\sa_snapshot[20][63] , \sa_snapshot[20][62] , \sa_snapshot[20][61] , 
	\sa_snapshot[20][60] , \sa_snapshot[20][59] , \sa_snapshot[20][58] , 
	\sa_snapshot[20][57] , \sa_snapshot[20][56] , \sa_snapshot[20][55] , 
	\sa_snapshot[20][54] , \sa_snapshot[20][53] , \sa_snapshot[20][52] , 
	\sa_snapshot[20][51] , \sa_snapshot[20][50] , \sa_snapshot[20][49] , 
	\sa_snapshot[20][48] , \sa_snapshot[20][47] , \sa_snapshot[20][46] , 
	\sa_snapshot[20][45] , \sa_snapshot[20][44] , \sa_snapshot[20][43] , 
	\sa_snapshot[20][42] , \sa_snapshot[20][41] , \sa_snapshot[20][40] , 
	\sa_snapshot[20][39] , \sa_snapshot[20][38] , \sa_snapshot[20][37] , 
	\sa_snapshot[20][36] , \sa_snapshot[20][35] , \sa_snapshot[20][34] , 
	\sa_snapshot[20][33] , \sa_snapshot[20][32] , \sa_snapshot[20][31] , 
	\sa_snapshot[20][30] , \sa_snapshot[20][29] , \sa_snapshot[20][28] , 
	\sa_snapshot[20][27] , \sa_snapshot[20][26] , \sa_snapshot[20][25] , 
	\sa_snapshot[20][24] , \sa_snapshot[20][23] , \sa_snapshot[20][22] , 
	\sa_snapshot[20][21] , \sa_snapshot[20][20] , \sa_snapshot[20][19] , 
	\sa_snapshot[20][18] , \sa_snapshot[20][17] , \sa_snapshot[20][16] , 
	\sa_snapshot[20][15] , \sa_snapshot[20][14] , \sa_snapshot[20][13] , 
	\sa_snapshot[20][12] , \sa_snapshot[20][11] , \sa_snapshot[20][10] , 
	\sa_snapshot[20][9] , \sa_snapshot[20][8] , \sa_snapshot[20][7] , 
	\sa_snapshot[20][6] , \sa_snapshot[20][5] , \sa_snapshot[20][4] , 
	\sa_snapshot[20][3] , \sa_snapshot[20][2] , \sa_snapshot[20][1] , 
	\sa_snapshot[20][0] , \sa_snapshot[19][63] , \sa_snapshot[19][62] , 
	\sa_snapshot[19][61] , \sa_snapshot[19][60] , \sa_snapshot[19][59] , 
	\sa_snapshot[19][58] , \sa_snapshot[19][57] , \sa_snapshot[19][56] , 
	\sa_snapshot[19][55] , \sa_snapshot[19][54] , \sa_snapshot[19][53] , 
	\sa_snapshot[19][52] , \sa_snapshot[19][51] , \sa_snapshot[19][50] , 
	\sa_snapshot[19][49] , \sa_snapshot[19][48] , \sa_snapshot[19][47] , 
	\sa_snapshot[19][46] , \sa_snapshot[19][45] , \sa_snapshot[19][44] , 
	\sa_snapshot[19][43] , \sa_snapshot[19][42] , \sa_snapshot[19][41] , 
	\sa_snapshot[19][40] , \sa_snapshot[19][39] , \sa_snapshot[19][38] , 
	\sa_snapshot[19][37] , \sa_snapshot[19][36] , \sa_snapshot[19][35] , 
	\sa_snapshot[19][34] , \sa_snapshot[19][33] , \sa_snapshot[19][32] , 
	\sa_snapshot[19][31] , \sa_snapshot[19][30] , \sa_snapshot[19][29] , 
	\sa_snapshot[19][28] , \sa_snapshot[19][27] , \sa_snapshot[19][26] , 
	\sa_snapshot[19][25] , \sa_snapshot[19][24] , \sa_snapshot[19][23] , 
	\sa_snapshot[19][22] , \sa_snapshot[19][21] , \sa_snapshot[19][20] , 
	\sa_snapshot[19][19] , \sa_snapshot[19][18] , \sa_snapshot[19][17] , 
	\sa_snapshot[19][16] , \sa_snapshot[19][15] , \sa_snapshot[19][14] , 
	\sa_snapshot[19][13] , \sa_snapshot[19][12] , \sa_snapshot[19][11] , 
	\sa_snapshot[19][10] , \sa_snapshot[19][9] , \sa_snapshot[19][8] , 
	\sa_snapshot[19][7] , \sa_snapshot[19][6] , \sa_snapshot[19][5] , 
	\sa_snapshot[19][4] , \sa_snapshot[19][3] , \sa_snapshot[19][2] , 
	\sa_snapshot[19][1] , \sa_snapshot[19][0] , \sa_snapshot[18][63] , 
	\sa_snapshot[18][62] , \sa_snapshot[18][61] , \sa_snapshot[18][60] , 
	\sa_snapshot[18][59] , \sa_snapshot[18][58] , \sa_snapshot[18][57] , 
	\sa_snapshot[18][56] , \sa_snapshot[18][55] , \sa_snapshot[18][54] , 
	\sa_snapshot[18][53] , \sa_snapshot[18][52] , \sa_snapshot[18][51] , 
	\sa_snapshot[18][50] , \sa_snapshot[18][49] , \sa_snapshot[18][48] , 
	\sa_snapshot[18][47] , \sa_snapshot[18][46] , \sa_snapshot[18][45] , 
	\sa_snapshot[18][44] , \sa_snapshot[18][43] , \sa_snapshot[18][42] , 
	\sa_snapshot[18][41] , \sa_snapshot[18][40] , \sa_snapshot[18][39] , 
	\sa_snapshot[18][38] , \sa_snapshot[18][37] , \sa_snapshot[18][36] , 
	\sa_snapshot[18][35] , \sa_snapshot[18][34] , \sa_snapshot[18][33] , 
	\sa_snapshot[18][32] , \sa_snapshot[18][31] , \sa_snapshot[18][30] , 
	\sa_snapshot[18][29] , \sa_snapshot[18][28] , \sa_snapshot[18][27] , 
	\sa_snapshot[18][26] , \sa_snapshot[18][25] , \sa_snapshot[18][24] , 
	\sa_snapshot[18][23] , \sa_snapshot[18][22] , \sa_snapshot[18][21] , 
	\sa_snapshot[18][20] , \sa_snapshot[18][19] , \sa_snapshot[18][18] , 
	\sa_snapshot[18][17] , \sa_snapshot[18][16] , \sa_snapshot[18][15] , 
	\sa_snapshot[18][14] , \sa_snapshot[18][13] , \sa_snapshot[18][12] , 
	\sa_snapshot[18][11] , \sa_snapshot[18][10] , \sa_snapshot[18][9] , 
	\sa_snapshot[18][8] , \sa_snapshot[18][7] , \sa_snapshot[18][6] , 
	\sa_snapshot[18][5] , \sa_snapshot[18][4] , \sa_snapshot[18][3] , 
	\sa_snapshot[18][2] , \sa_snapshot[18][1] , \sa_snapshot[18][0] , 
	\sa_snapshot[17][63] , \sa_snapshot[17][62] , \sa_snapshot[17][61] , 
	\sa_snapshot[17][60] , \sa_snapshot[17][59] , \sa_snapshot[17][58] , 
	\sa_snapshot[17][57] , \sa_snapshot[17][56] , \sa_snapshot[17][55] , 
	\sa_snapshot[17][54] , \sa_snapshot[17][53] , \sa_snapshot[17][52] , 
	\sa_snapshot[17][51] , \sa_snapshot[17][50] , \sa_snapshot[17][49] , 
	\sa_snapshot[17][48] , \sa_snapshot[17][47] , \sa_snapshot[17][46] , 
	\sa_snapshot[17][45] , \sa_snapshot[17][44] , \sa_snapshot[17][43] , 
	\sa_snapshot[17][42] , \sa_snapshot[17][41] , \sa_snapshot[17][40] , 
	\sa_snapshot[17][39] , \sa_snapshot[17][38] , \sa_snapshot[17][37] , 
	\sa_snapshot[17][36] , \sa_snapshot[17][35] , \sa_snapshot[17][34] , 
	\sa_snapshot[17][33] , \sa_snapshot[17][32] , \sa_snapshot[17][31] , 
	\sa_snapshot[17][30] , \sa_snapshot[17][29] , \sa_snapshot[17][28] , 
	\sa_snapshot[17][27] , \sa_snapshot[17][26] , \sa_snapshot[17][25] , 
	\sa_snapshot[17][24] , \sa_snapshot[17][23] , \sa_snapshot[17][22] , 
	\sa_snapshot[17][21] , \sa_snapshot[17][20] , \sa_snapshot[17][19] , 
	\sa_snapshot[17][18] , \sa_snapshot[17][17] , \sa_snapshot[17][16] , 
	\sa_snapshot[17][15] , \sa_snapshot[17][14] , \sa_snapshot[17][13] , 
	\sa_snapshot[17][12] , \sa_snapshot[17][11] , \sa_snapshot[17][10] , 
	\sa_snapshot[17][9] , \sa_snapshot[17][8] , \sa_snapshot[17][7] , 
	\sa_snapshot[17][6] , \sa_snapshot[17][5] , \sa_snapshot[17][4] , 
	\sa_snapshot[17][3] , \sa_snapshot[17][2] , \sa_snapshot[17][1] , 
	\sa_snapshot[17][0] , \sa_snapshot[16][63] , \sa_snapshot[16][62] , 
	\sa_snapshot[16][61] , \sa_snapshot[16][60] , \sa_snapshot[16][59] , 
	\sa_snapshot[16][58] , \sa_snapshot[16][57] , \sa_snapshot[16][56] , 
	\sa_snapshot[16][55] , \sa_snapshot[16][54] , \sa_snapshot[16][53] , 
	\sa_snapshot[16][52] , \sa_snapshot[16][51] , \sa_snapshot[16][50] , 
	\sa_snapshot[16][49] , \sa_snapshot[16][48] , \sa_snapshot[16][47] , 
	\sa_snapshot[16][46] , \sa_snapshot[16][45] , \sa_snapshot[16][44] , 
	\sa_snapshot[16][43] , \sa_snapshot[16][42] , \sa_snapshot[16][41] , 
	\sa_snapshot[16][40] , \sa_snapshot[16][39] , \sa_snapshot[16][38] , 
	\sa_snapshot[16][37] , \sa_snapshot[16][36] , \sa_snapshot[16][35] , 
	\sa_snapshot[16][34] , \sa_snapshot[16][33] , \sa_snapshot[16][32] , 
	\sa_snapshot[16][31] , \sa_snapshot[16][30] , \sa_snapshot[16][29] , 
	\sa_snapshot[16][28] , \sa_snapshot[16][27] , \sa_snapshot[16][26] , 
	\sa_snapshot[16][25] , \sa_snapshot[16][24] , \sa_snapshot[16][23] , 
	\sa_snapshot[16][22] , \sa_snapshot[16][21] , \sa_snapshot[16][20] , 
	\sa_snapshot[16][19] , \sa_snapshot[16][18] , \sa_snapshot[16][17] , 
	\sa_snapshot[16][16] , \sa_snapshot[16][15] , \sa_snapshot[16][14] , 
	\sa_snapshot[16][13] , \sa_snapshot[16][12] , \sa_snapshot[16][11] , 
	\sa_snapshot[16][10] , \sa_snapshot[16][9] , \sa_snapshot[16][8] , 
	\sa_snapshot[16][7] , \sa_snapshot[16][6] , \sa_snapshot[16][5] , 
	\sa_snapshot[16][4] , \sa_snapshot[16][3] , \sa_snapshot[16][2] , 
	\sa_snapshot[16][1] , \sa_snapshot[16][0] , \sa_snapshot[15][63] , 
	\sa_snapshot[15][62] , \sa_snapshot[15][61] , \sa_snapshot[15][60] , 
	\sa_snapshot[15][59] , \sa_snapshot[15][58] , \sa_snapshot[15][57] , 
	\sa_snapshot[15][56] , \sa_snapshot[15][55] , \sa_snapshot[15][54] , 
	\sa_snapshot[15][53] , \sa_snapshot[15][52] , \sa_snapshot[15][51] , 
	\sa_snapshot[15][50] , \sa_snapshot[15][49] , \sa_snapshot[15][48] , 
	\sa_snapshot[15][47] , \sa_snapshot[15][46] , \sa_snapshot[15][45] , 
	\sa_snapshot[15][44] , \sa_snapshot[15][43] , \sa_snapshot[15][42] , 
	\sa_snapshot[15][41] , \sa_snapshot[15][40] , \sa_snapshot[15][39] , 
	\sa_snapshot[15][38] , \sa_snapshot[15][37] , \sa_snapshot[15][36] , 
	\sa_snapshot[15][35] , \sa_snapshot[15][34] , \sa_snapshot[15][33] , 
	\sa_snapshot[15][32] , \sa_snapshot[15][31] , \sa_snapshot[15][30] , 
	\sa_snapshot[15][29] , \sa_snapshot[15][28] , \sa_snapshot[15][27] , 
	\sa_snapshot[15][26] , \sa_snapshot[15][25] , \sa_snapshot[15][24] , 
	\sa_snapshot[15][23] , \sa_snapshot[15][22] , \sa_snapshot[15][21] , 
	\sa_snapshot[15][20] , \sa_snapshot[15][19] , \sa_snapshot[15][18] , 
	\sa_snapshot[15][17] , \sa_snapshot[15][16] , \sa_snapshot[15][15] , 
	\sa_snapshot[15][14] , \sa_snapshot[15][13] , \sa_snapshot[15][12] , 
	\sa_snapshot[15][11] , \sa_snapshot[15][10] , \sa_snapshot[15][9] , 
	\sa_snapshot[15][8] , \sa_snapshot[15][7] , \sa_snapshot[15][6] , 
	\sa_snapshot[15][5] , \sa_snapshot[15][4] , \sa_snapshot[15][3] , 
	\sa_snapshot[15][2] , \sa_snapshot[15][1] , \sa_snapshot[15][0] , 
	\sa_snapshot[14][63] , \sa_snapshot[14][62] , \sa_snapshot[14][61] , 
	\sa_snapshot[14][60] , \sa_snapshot[14][59] , \sa_snapshot[14][58] , 
	\sa_snapshot[14][57] , \sa_snapshot[14][56] , \sa_snapshot[14][55] , 
	\sa_snapshot[14][54] , \sa_snapshot[14][53] , \sa_snapshot[14][52] , 
	\sa_snapshot[14][51] , \sa_snapshot[14][50] , \sa_snapshot[14][49] , 
	\sa_snapshot[14][48] , \sa_snapshot[14][47] , \sa_snapshot[14][46] , 
	\sa_snapshot[14][45] , \sa_snapshot[14][44] , \sa_snapshot[14][43] , 
	\sa_snapshot[14][42] , \sa_snapshot[14][41] , \sa_snapshot[14][40] , 
	\sa_snapshot[14][39] , \sa_snapshot[14][38] , \sa_snapshot[14][37] , 
	\sa_snapshot[14][36] , \sa_snapshot[14][35] , \sa_snapshot[14][34] , 
	\sa_snapshot[14][33] , \sa_snapshot[14][32] , \sa_snapshot[14][31] , 
	\sa_snapshot[14][30] , \sa_snapshot[14][29] , \sa_snapshot[14][28] , 
	\sa_snapshot[14][27] , \sa_snapshot[14][26] , \sa_snapshot[14][25] , 
	\sa_snapshot[14][24] , \sa_snapshot[14][23] , \sa_snapshot[14][22] , 
	\sa_snapshot[14][21] , \sa_snapshot[14][20] , \sa_snapshot[14][19] , 
	\sa_snapshot[14][18] , \sa_snapshot[14][17] , \sa_snapshot[14][16] , 
	\sa_snapshot[14][15] , \sa_snapshot[14][14] , \sa_snapshot[14][13] , 
	\sa_snapshot[14][12] , \sa_snapshot[14][11] , \sa_snapshot[14][10] , 
	\sa_snapshot[14][9] , \sa_snapshot[14][8] , \sa_snapshot[14][7] , 
	\sa_snapshot[14][6] , \sa_snapshot[14][5] , \sa_snapshot[14][4] , 
	\sa_snapshot[14][3] , \sa_snapshot[14][2] , \sa_snapshot[14][1] , 
	\sa_snapshot[14][0] , \sa_snapshot[13][63] , \sa_snapshot[13][62] , 
	\sa_snapshot[13][61] , \sa_snapshot[13][60] , \sa_snapshot[13][59] , 
	\sa_snapshot[13][58] , \sa_snapshot[13][57] , \sa_snapshot[13][56] , 
	\sa_snapshot[13][55] , \sa_snapshot[13][54] , \sa_snapshot[13][53] , 
	\sa_snapshot[13][52] , \sa_snapshot[13][51] , \sa_snapshot[13][50] , 
	\sa_snapshot[13][49] , \sa_snapshot[13][48] , \sa_snapshot[13][47] , 
	\sa_snapshot[13][46] , \sa_snapshot[13][45] , \sa_snapshot[13][44] , 
	\sa_snapshot[13][43] , \sa_snapshot[13][42] , \sa_snapshot[13][41] , 
	\sa_snapshot[13][40] , \sa_snapshot[13][39] , \sa_snapshot[13][38] , 
	\sa_snapshot[13][37] , \sa_snapshot[13][36] , \sa_snapshot[13][35] , 
	\sa_snapshot[13][34] , \sa_snapshot[13][33] , \sa_snapshot[13][32] , 
	\sa_snapshot[13][31] , \sa_snapshot[13][30] , \sa_snapshot[13][29] , 
	\sa_snapshot[13][28] , \sa_snapshot[13][27] , \sa_snapshot[13][26] , 
	\sa_snapshot[13][25] , \sa_snapshot[13][24] , \sa_snapshot[13][23] , 
	\sa_snapshot[13][22] , \sa_snapshot[13][21] , \sa_snapshot[13][20] , 
	\sa_snapshot[13][19] , \sa_snapshot[13][18] , \sa_snapshot[13][17] , 
	\sa_snapshot[13][16] , \sa_snapshot[13][15] , \sa_snapshot[13][14] , 
	\sa_snapshot[13][13] , \sa_snapshot[13][12] , \sa_snapshot[13][11] , 
	\sa_snapshot[13][10] , \sa_snapshot[13][9] , \sa_snapshot[13][8] , 
	\sa_snapshot[13][7] , \sa_snapshot[13][6] , \sa_snapshot[13][5] , 
	\sa_snapshot[13][4] , \sa_snapshot[13][3] , \sa_snapshot[13][2] , 
	\sa_snapshot[13][1] , \sa_snapshot[13][0] , \sa_snapshot[12][63] , 
	\sa_snapshot[12][62] , \sa_snapshot[12][61] , \sa_snapshot[12][60] , 
	\sa_snapshot[12][59] , \sa_snapshot[12][58] , \sa_snapshot[12][57] , 
	\sa_snapshot[12][56] , \sa_snapshot[12][55] , \sa_snapshot[12][54] , 
	\sa_snapshot[12][53] , \sa_snapshot[12][52] , \sa_snapshot[12][51] , 
	\sa_snapshot[12][50] , \sa_snapshot[12][49] , \sa_snapshot[12][48] , 
	\sa_snapshot[12][47] , \sa_snapshot[12][46] , \sa_snapshot[12][45] , 
	\sa_snapshot[12][44] , \sa_snapshot[12][43] , \sa_snapshot[12][42] , 
	\sa_snapshot[12][41] , \sa_snapshot[12][40] , \sa_snapshot[12][39] , 
	\sa_snapshot[12][38] , \sa_snapshot[12][37] , \sa_snapshot[12][36] , 
	\sa_snapshot[12][35] , \sa_snapshot[12][34] , \sa_snapshot[12][33] , 
	\sa_snapshot[12][32] , \sa_snapshot[12][31] , \sa_snapshot[12][30] , 
	\sa_snapshot[12][29] , \sa_snapshot[12][28] , \sa_snapshot[12][27] , 
	\sa_snapshot[12][26] , \sa_snapshot[12][25] , \sa_snapshot[12][24] , 
	\sa_snapshot[12][23] , \sa_snapshot[12][22] , \sa_snapshot[12][21] , 
	\sa_snapshot[12][20] , \sa_snapshot[12][19] , \sa_snapshot[12][18] , 
	\sa_snapshot[12][17] , \sa_snapshot[12][16] , \sa_snapshot[12][15] , 
	\sa_snapshot[12][14] , \sa_snapshot[12][13] , \sa_snapshot[12][12] , 
	\sa_snapshot[12][11] , \sa_snapshot[12][10] , \sa_snapshot[12][9] , 
	\sa_snapshot[12][8] , \sa_snapshot[12][7] , \sa_snapshot[12][6] , 
	\sa_snapshot[12][5] , \sa_snapshot[12][4] , \sa_snapshot[12][3] , 
	\sa_snapshot[12][2] , \sa_snapshot[12][1] , \sa_snapshot[12][0] , 
	\sa_snapshot[11][63] , \sa_snapshot[11][62] , \sa_snapshot[11][61] , 
	\sa_snapshot[11][60] , \sa_snapshot[11][59] , \sa_snapshot[11][58] , 
	\sa_snapshot[11][57] , \sa_snapshot[11][56] , \sa_snapshot[11][55] , 
	\sa_snapshot[11][54] , \sa_snapshot[11][53] , \sa_snapshot[11][52] , 
	\sa_snapshot[11][51] , \sa_snapshot[11][50] , \sa_snapshot[11][49] , 
	\sa_snapshot[11][48] , \sa_snapshot[11][47] , \sa_snapshot[11][46] , 
	\sa_snapshot[11][45] , \sa_snapshot[11][44] , \sa_snapshot[11][43] , 
	\sa_snapshot[11][42] , \sa_snapshot[11][41] , \sa_snapshot[11][40] , 
	\sa_snapshot[11][39] , \sa_snapshot[11][38] , \sa_snapshot[11][37] , 
	\sa_snapshot[11][36] , \sa_snapshot[11][35] , \sa_snapshot[11][34] , 
	\sa_snapshot[11][33] , \sa_snapshot[11][32] , \sa_snapshot[11][31] , 
	\sa_snapshot[11][30] , \sa_snapshot[11][29] , \sa_snapshot[11][28] , 
	\sa_snapshot[11][27] , \sa_snapshot[11][26] , \sa_snapshot[11][25] , 
	\sa_snapshot[11][24] , \sa_snapshot[11][23] , \sa_snapshot[11][22] , 
	\sa_snapshot[11][21] , \sa_snapshot[11][20] , \sa_snapshot[11][19] , 
	\sa_snapshot[11][18] , \sa_snapshot[11][17] , \sa_snapshot[11][16] , 
	\sa_snapshot[11][15] , \sa_snapshot[11][14] , \sa_snapshot[11][13] , 
	\sa_snapshot[11][12] , \sa_snapshot[11][11] , \sa_snapshot[11][10] , 
	\sa_snapshot[11][9] , \sa_snapshot[11][8] , \sa_snapshot[11][7] , 
	\sa_snapshot[11][6] , \sa_snapshot[11][5] , \sa_snapshot[11][4] , 
	\sa_snapshot[11][3] , \sa_snapshot[11][2] , \sa_snapshot[11][1] , 
	\sa_snapshot[11][0] , \sa_snapshot[10][63] , \sa_snapshot[10][62] , 
	\sa_snapshot[10][61] , \sa_snapshot[10][60] , \sa_snapshot[10][59] , 
	\sa_snapshot[10][58] , \sa_snapshot[10][57] , \sa_snapshot[10][56] , 
	\sa_snapshot[10][55] , \sa_snapshot[10][54] , \sa_snapshot[10][53] , 
	\sa_snapshot[10][52] , \sa_snapshot[10][51] , \sa_snapshot[10][50] , 
	\sa_snapshot[10][49] , \sa_snapshot[10][48] , \sa_snapshot[10][47] , 
	\sa_snapshot[10][46] , \sa_snapshot[10][45] , \sa_snapshot[10][44] , 
	\sa_snapshot[10][43] , \sa_snapshot[10][42] , \sa_snapshot[10][41] , 
	\sa_snapshot[10][40] , \sa_snapshot[10][39] , \sa_snapshot[10][38] , 
	\sa_snapshot[10][37] , \sa_snapshot[10][36] , \sa_snapshot[10][35] , 
	\sa_snapshot[10][34] , \sa_snapshot[10][33] , \sa_snapshot[10][32] , 
	\sa_snapshot[10][31] , \sa_snapshot[10][30] , \sa_snapshot[10][29] , 
	\sa_snapshot[10][28] , \sa_snapshot[10][27] , \sa_snapshot[10][26] , 
	\sa_snapshot[10][25] , \sa_snapshot[10][24] , \sa_snapshot[10][23] , 
	\sa_snapshot[10][22] , \sa_snapshot[10][21] , \sa_snapshot[10][20] , 
	\sa_snapshot[10][19] , \sa_snapshot[10][18] , \sa_snapshot[10][17] , 
	\sa_snapshot[10][16] , \sa_snapshot[10][15] , \sa_snapshot[10][14] , 
	\sa_snapshot[10][13] , \sa_snapshot[10][12] , \sa_snapshot[10][11] , 
	\sa_snapshot[10][10] , \sa_snapshot[10][9] , \sa_snapshot[10][8] , 
	\sa_snapshot[10][7] , \sa_snapshot[10][6] , \sa_snapshot[10][5] , 
	\sa_snapshot[10][4] , \sa_snapshot[10][3] , \sa_snapshot[10][2] , 
	\sa_snapshot[10][1] , \sa_snapshot[10][0] , \sa_snapshot[9][63] , 
	\sa_snapshot[9][62] , \sa_snapshot[9][61] , \sa_snapshot[9][60] , 
	\sa_snapshot[9][59] , \sa_snapshot[9][58] , \sa_snapshot[9][57] , 
	\sa_snapshot[9][56] , \sa_snapshot[9][55] , \sa_snapshot[9][54] , 
	\sa_snapshot[9][53] , \sa_snapshot[9][52] , \sa_snapshot[9][51] , 
	\sa_snapshot[9][50] , \sa_snapshot[9][49] , \sa_snapshot[9][48] , 
	\sa_snapshot[9][47] , \sa_snapshot[9][46] , \sa_snapshot[9][45] , 
	\sa_snapshot[9][44] , \sa_snapshot[9][43] , \sa_snapshot[9][42] , 
	\sa_snapshot[9][41] , \sa_snapshot[9][40] , \sa_snapshot[9][39] , 
	\sa_snapshot[9][38] , \sa_snapshot[9][37] , \sa_snapshot[9][36] , 
	\sa_snapshot[9][35] , \sa_snapshot[9][34] , \sa_snapshot[9][33] , 
	\sa_snapshot[9][32] , \sa_snapshot[9][31] , \sa_snapshot[9][30] , 
	\sa_snapshot[9][29] , \sa_snapshot[9][28] , \sa_snapshot[9][27] , 
	\sa_snapshot[9][26] , \sa_snapshot[9][25] , \sa_snapshot[9][24] , 
	\sa_snapshot[9][23] , \sa_snapshot[9][22] , \sa_snapshot[9][21] , 
	\sa_snapshot[9][20] , \sa_snapshot[9][19] , \sa_snapshot[9][18] , 
	\sa_snapshot[9][17] , \sa_snapshot[9][16] , \sa_snapshot[9][15] , 
	\sa_snapshot[9][14] , \sa_snapshot[9][13] , \sa_snapshot[9][12] , 
	\sa_snapshot[9][11] , \sa_snapshot[9][10] , \sa_snapshot[9][9] , 
	\sa_snapshot[9][8] , \sa_snapshot[9][7] , \sa_snapshot[9][6] , 
	\sa_snapshot[9][5] , \sa_snapshot[9][4] , \sa_snapshot[9][3] , 
	\sa_snapshot[9][2] , \sa_snapshot[9][1] , \sa_snapshot[9][0] , 
	\sa_snapshot[8][63] , \sa_snapshot[8][62] , \sa_snapshot[8][61] , 
	\sa_snapshot[8][60] , \sa_snapshot[8][59] , \sa_snapshot[8][58] , 
	\sa_snapshot[8][57] , \sa_snapshot[8][56] , \sa_snapshot[8][55] , 
	\sa_snapshot[8][54] , \sa_snapshot[8][53] , \sa_snapshot[8][52] , 
	\sa_snapshot[8][51] , \sa_snapshot[8][50] , \sa_snapshot[8][49] , 
	\sa_snapshot[8][48] , \sa_snapshot[8][47] , \sa_snapshot[8][46] , 
	\sa_snapshot[8][45] , \sa_snapshot[8][44] , \sa_snapshot[8][43] , 
	\sa_snapshot[8][42] , \sa_snapshot[8][41] , \sa_snapshot[8][40] , 
	\sa_snapshot[8][39] , \sa_snapshot[8][38] , \sa_snapshot[8][37] , 
	\sa_snapshot[8][36] , \sa_snapshot[8][35] , \sa_snapshot[8][34] , 
	\sa_snapshot[8][33] , \sa_snapshot[8][32] , \sa_snapshot[8][31] , 
	\sa_snapshot[8][30] , \sa_snapshot[8][29] , \sa_snapshot[8][28] , 
	\sa_snapshot[8][27] , \sa_snapshot[8][26] , \sa_snapshot[8][25] , 
	\sa_snapshot[8][24] , \sa_snapshot[8][23] , \sa_snapshot[8][22] , 
	\sa_snapshot[8][21] , \sa_snapshot[8][20] , \sa_snapshot[8][19] , 
	\sa_snapshot[8][18] , \sa_snapshot[8][17] , \sa_snapshot[8][16] , 
	\sa_snapshot[8][15] , \sa_snapshot[8][14] , \sa_snapshot[8][13] , 
	\sa_snapshot[8][12] , \sa_snapshot[8][11] , \sa_snapshot[8][10] , 
	\sa_snapshot[8][9] , \sa_snapshot[8][8] , \sa_snapshot[8][7] , 
	\sa_snapshot[8][6] , \sa_snapshot[8][5] , \sa_snapshot[8][4] , 
	\sa_snapshot[8][3] , \sa_snapshot[8][2] , \sa_snapshot[8][1] , 
	\sa_snapshot[8][0] , \sa_snapshot[7][63] , \sa_snapshot[7][62] , 
	\sa_snapshot[7][61] , \sa_snapshot[7][60] , \sa_snapshot[7][59] , 
	\sa_snapshot[7][58] , \sa_snapshot[7][57] , \sa_snapshot[7][56] , 
	\sa_snapshot[7][55] , \sa_snapshot[7][54] , \sa_snapshot[7][53] , 
	\sa_snapshot[7][52] , \sa_snapshot[7][51] , \sa_snapshot[7][50] , 
	\sa_snapshot[7][49] , \sa_snapshot[7][48] , \sa_snapshot[7][47] , 
	\sa_snapshot[7][46] , \sa_snapshot[7][45] , \sa_snapshot[7][44] , 
	\sa_snapshot[7][43] , \sa_snapshot[7][42] , \sa_snapshot[7][41] , 
	\sa_snapshot[7][40] , \sa_snapshot[7][39] , \sa_snapshot[7][38] , 
	\sa_snapshot[7][37] , \sa_snapshot[7][36] , \sa_snapshot[7][35] , 
	\sa_snapshot[7][34] , \sa_snapshot[7][33] , \sa_snapshot[7][32] , 
	\sa_snapshot[7][31] , \sa_snapshot[7][30] , \sa_snapshot[7][29] , 
	\sa_snapshot[7][28] , \sa_snapshot[7][27] , \sa_snapshot[7][26] , 
	\sa_snapshot[7][25] , \sa_snapshot[7][24] , \sa_snapshot[7][23] , 
	\sa_snapshot[7][22] , \sa_snapshot[7][21] , \sa_snapshot[7][20] , 
	\sa_snapshot[7][19] , \sa_snapshot[7][18] , \sa_snapshot[7][17] , 
	\sa_snapshot[7][16] , \sa_snapshot[7][15] , \sa_snapshot[7][14] , 
	\sa_snapshot[7][13] , \sa_snapshot[7][12] , \sa_snapshot[7][11] , 
	\sa_snapshot[7][10] , \sa_snapshot[7][9] , \sa_snapshot[7][8] , 
	\sa_snapshot[7][7] , \sa_snapshot[7][6] , \sa_snapshot[7][5] , 
	\sa_snapshot[7][4] , \sa_snapshot[7][3] , \sa_snapshot[7][2] , 
	\sa_snapshot[7][1] , \sa_snapshot[7][0] , \sa_snapshot[6][63] , 
	\sa_snapshot[6][62] , \sa_snapshot[6][61] , \sa_snapshot[6][60] , 
	\sa_snapshot[6][59] , \sa_snapshot[6][58] , \sa_snapshot[6][57] , 
	\sa_snapshot[6][56] , \sa_snapshot[6][55] , \sa_snapshot[6][54] , 
	\sa_snapshot[6][53] , \sa_snapshot[6][52] , \sa_snapshot[6][51] , 
	\sa_snapshot[6][50] , \sa_snapshot[6][49] , \sa_snapshot[6][48] , 
	\sa_snapshot[6][47] , \sa_snapshot[6][46] , \sa_snapshot[6][45] , 
	\sa_snapshot[6][44] , \sa_snapshot[6][43] , \sa_snapshot[6][42] , 
	\sa_snapshot[6][41] , \sa_snapshot[6][40] , \sa_snapshot[6][39] , 
	\sa_snapshot[6][38] , \sa_snapshot[6][37] , \sa_snapshot[6][36] , 
	\sa_snapshot[6][35] , \sa_snapshot[6][34] , \sa_snapshot[6][33] , 
	\sa_snapshot[6][32] , \sa_snapshot[6][31] , \sa_snapshot[6][30] , 
	\sa_snapshot[6][29] , \sa_snapshot[6][28] , \sa_snapshot[6][27] , 
	\sa_snapshot[6][26] , \sa_snapshot[6][25] , \sa_snapshot[6][24] , 
	\sa_snapshot[6][23] , \sa_snapshot[6][22] , \sa_snapshot[6][21] , 
	\sa_snapshot[6][20] , \sa_snapshot[6][19] , \sa_snapshot[6][18] , 
	\sa_snapshot[6][17] , \sa_snapshot[6][16] , \sa_snapshot[6][15] , 
	\sa_snapshot[6][14] , \sa_snapshot[6][13] , \sa_snapshot[6][12] , 
	\sa_snapshot[6][11] , \sa_snapshot[6][10] , \sa_snapshot[6][9] , 
	\sa_snapshot[6][8] , \sa_snapshot[6][7] , \sa_snapshot[6][6] , 
	\sa_snapshot[6][5] , \sa_snapshot[6][4] , \sa_snapshot[6][3] , 
	\sa_snapshot[6][2] , \sa_snapshot[6][1] , \sa_snapshot[6][0] , 
	\sa_snapshot[5][63] , \sa_snapshot[5][62] , \sa_snapshot[5][61] , 
	\sa_snapshot[5][60] , \sa_snapshot[5][59] , \sa_snapshot[5][58] , 
	\sa_snapshot[5][57] , \sa_snapshot[5][56] , \sa_snapshot[5][55] , 
	\sa_snapshot[5][54] , \sa_snapshot[5][53] , \sa_snapshot[5][52] , 
	\sa_snapshot[5][51] , \sa_snapshot[5][50] , \sa_snapshot[5][49] , 
	\sa_snapshot[5][48] , \sa_snapshot[5][47] , \sa_snapshot[5][46] , 
	\sa_snapshot[5][45] , \sa_snapshot[5][44] , \sa_snapshot[5][43] , 
	\sa_snapshot[5][42] , \sa_snapshot[5][41] , \sa_snapshot[5][40] , 
	\sa_snapshot[5][39] , \sa_snapshot[5][38] , \sa_snapshot[5][37] , 
	\sa_snapshot[5][36] , \sa_snapshot[5][35] , \sa_snapshot[5][34] , 
	\sa_snapshot[5][33] , \sa_snapshot[5][32] , \sa_snapshot[5][31] , 
	\sa_snapshot[5][30] , \sa_snapshot[5][29] , \sa_snapshot[5][28] , 
	\sa_snapshot[5][27] , \sa_snapshot[5][26] , \sa_snapshot[5][25] , 
	\sa_snapshot[5][24] , \sa_snapshot[5][23] , \sa_snapshot[5][22] , 
	\sa_snapshot[5][21] , \sa_snapshot[5][20] , \sa_snapshot[5][19] , 
	\sa_snapshot[5][18] , \sa_snapshot[5][17] , \sa_snapshot[5][16] , 
	\sa_snapshot[5][15] , \sa_snapshot[5][14] , \sa_snapshot[5][13] , 
	\sa_snapshot[5][12] , \sa_snapshot[5][11] , \sa_snapshot[5][10] , 
	\sa_snapshot[5][9] , \sa_snapshot[5][8] , \sa_snapshot[5][7] , 
	\sa_snapshot[5][6] , \sa_snapshot[5][5] , \sa_snapshot[5][4] , 
	\sa_snapshot[5][3] , \sa_snapshot[5][2] , \sa_snapshot[5][1] , 
	\sa_snapshot[5][0] , \sa_snapshot[4][63] , \sa_snapshot[4][62] , 
	\sa_snapshot[4][61] , \sa_snapshot[4][60] , \sa_snapshot[4][59] , 
	\sa_snapshot[4][58] , \sa_snapshot[4][57] , \sa_snapshot[4][56] , 
	\sa_snapshot[4][55] , \sa_snapshot[4][54] , \sa_snapshot[4][53] , 
	\sa_snapshot[4][52] , \sa_snapshot[4][51] , \sa_snapshot[4][50] , 
	\sa_snapshot[4][49] , \sa_snapshot[4][48] , \sa_snapshot[4][47] , 
	\sa_snapshot[4][46] , \sa_snapshot[4][45] , \sa_snapshot[4][44] , 
	\sa_snapshot[4][43] , \sa_snapshot[4][42] , \sa_snapshot[4][41] , 
	\sa_snapshot[4][40] , \sa_snapshot[4][39] , \sa_snapshot[4][38] , 
	\sa_snapshot[4][37] , \sa_snapshot[4][36] , \sa_snapshot[4][35] , 
	\sa_snapshot[4][34] , \sa_snapshot[4][33] , \sa_snapshot[4][32] , 
	\sa_snapshot[4][31] , \sa_snapshot[4][30] , \sa_snapshot[4][29] , 
	\sa_snapshot[4][28] , \sa_snapshot[4][27] , \sa_snapshot[4][26] , 
	\sa_snapshot[4][25] , \sa_snapshot[4][24] , \sa_snapshot[4][23] , 
	\sa_snapshot[4][22] , \sa_snapshot[4][21] , \sa_snapshot[4][20] , 
	\sa_snapshot[4][19] , \sa_snapshot[4][18] , \sa_snapshot[4][17] , 
	\sa_snapshot[4][16] , \sa_snapshot[4][15] , \sa_snapshot[4][14] , 
	\sa_snapshot[4][13] , \sa_snapshot[4][12] , \sa_snapshot[4][11] , 
	\sa_snapshot[4][10] , \sa_snapshot[4][9] , \sa_snapshot[4][8] , 
	\sa_snapshot[4][7] , \sa_snapshot[4][6] , \sa_snapshot[4][5] , 
	\sa_snapshot[4][4] , \sa_snapshot[4][3] , \sa_snapshot[4][2] , 
	\sa_snapshot[4][1] , \sa_snapshot[4][0] , \sa_snapshot[3][63] , 
	\sa_snapshot[3][62] , \sa_snapshot[3][61] , \sa_snapshot[3][60] , 
	\sa_snapshot[3][59] , \sa_snapshot[3][58] , \sa_snapshot[3][57] , 
	\sa_snapshot[3][56] , \sa_snapshot[3][55] , \sa_snapshot[3][54] , 
	\sa_snapshot[3][53] , \sa_snapshot[3][52] , \sa_snapshot[3][51] , 
	\sa_snapshot[3][50] , \sa_snapshot[3][49] , \sa_snapshot[3][48] , 
	\sa_snapshot[3][47] , \sa_snapshot[3][46] , \sa_snapshot[3][45] , 
	\sa_snapshot[3][44] , \sa_snapshot[3][43] , \sa_snapshot[3][42] , 
	\sa_snapshot[3][41] , \sa_snapshot[3][40] , \sa_snapshot[3][39] , 
	\sa_snapshot[3][38] , \sa_snapshot[3][37] , \sa_snapshot[3][36] , 
	\sa_snapshot[3][35] , \sa_snapshot[3][34] , \sa_snapshot[3][33] , 
	\sa_snapshot[3][32] , \sa_snapshot[3][31] , \sa_snapshot[3][30] , 
	\sa_snapshot[3][29] , \sa_snapshot[3][28] , \sa_snapshot[3][27] , 
	\sa_snapshot[3][26] , \sa_snapshot[3][25] , \sa_snapshot[3][24] , 
	\sa_snapshot[3][23] , \sa_snapshot[3][22] , \sa_snapshot[3][21] , 
	\sa_snapshot[3][20] , \sa_snapshot[3][19] , \sa_snapshot[3][18] , 
	\sa_snapshot[3][17] , \sa_snapshot[3][16] , \sa_snapshot[3][15] , 
	\sa_snapshot[3][14] , \sa_snapshot[3][13] , \sa_snapshot[3][12] , 
	\sa_snapshot[3][11] , \sa_snapshot[3][10] , \sa_snapshot[3][9] , 
	\sa_snapshot[3][8] , \sa_snapshot[3][7] , \sa_snapshot[3][6] , 
	\sa_snapshot[3][5] , \sa_snapshot[3][4] , \sa_snapshot[3][3] , 
	\sa_snapshot[3][2] , \sa_snapshot[3][1] , \sa_snapshot[3][0] , 
	\sa_snapshot[2][63] , \sa_snapshot[2][62] , \sa_snapshot[2][61] , 
	\sa_snapshot[2][60] , \sa_snapshot[2][59] , \sa_snapshot[2][58] , 
	\sa_snapshot[2][57] , \sa_snapshot[2][56] , \sa_snapshot[2][55] , 
	\sa_snapshot[2][54] , \sa_snapshot[2][53] , \sa_snapshot[2][52] , 
	\sa_snapshot[2][51] , \sa_snapshot[2][50] , \sa_snapshot[2][49] , 
	\sa_snapshot[2][48] , \sa_snapshot[2][47] , \sa_snapshot[2][46] , 
	\sa_snapshot[2][45] , \sa_snapshot[2][44] , \sa_snapshot[2][43] , 
	\sa_snapshot[2][42] , \sa_snapshot[2][41] , \sa_snapshot[2][40] , 
	\sa_snapshot[2][39] , \sa_snapshot[2][38] , \sa_snapshot[2][37] , 
	\sa_snapshot[2][36] , \sa_snapshot[2][35] , \sa_snapshot[2][34] , 
	\sa_snapshot[2][33] , \sa_snapshot[2][32] , \sa_snapshot[2][31] , 
	\sa_snapshot[2][30] , \sa_snapshot[2][29] , \sa_snapshot[2][28] , 
	\sa_snapshot[2][27] , \sa_snapshot[2][26] , \sa_snapshot[2][25] , 
	\sa_snapshot[2][24] , \sa_snapshot[2][23] , \sa_snapshot[2][22] , 
	\sa_snapshot[2][21] , \sa_snapshot[2][20] , \sa_snapshot[2][19] , 
	\sa_snapshot[2][18] , \sa_snapshot[2][17] , \sa_snapshot[2][16] , 
	\sa_snapshot[2][15] , \sa_snapshot[2][14] , \sa_snapshot[2][13] , 
	\sa_snapshot[2][12] , \sa_snapshot[2][11] , \sa_snapshot[2][10] , 
	\sa_snapshot[2][9] , \sa_snapshot[2][8] , \sa_snapshot[2][7] , 
	\sa_snapshot[2][6] , \sa_snapshot[2][5] , \sa_snapshot[2][4] , 
	\sa_snapshot[2][3] , \sa_snapshot[2][2] , \sa_snapshot[2][1] , 
	\sa_snapshot[2][0] , \sa_snapshot[1][63] , \sa_snapshot[1][62] , 
	\sa_snapshot[1][61] , \sa_snapshot[1][60] , \sa_snapshot[1][59] , 
	\sa_snapshot[1][58] , \sa_snapshot[1][57] , \sa_snapshot[1][56] , 
	\sa_snapshot[1][55] , \sa_snapshot[1][54] , \sa_snapshot[1][53] , 
	\sa_snapshot[1][52] , \sa_snapshot[1][51] , \sa_snapshot[1][50] , 
	\sa_snapshot[1][49] , \sa_snapshot[1][48] , \sa_snapshot[1][47] , 
	\sa_snapshot[1][46] , \sa_snapshot[1][45] , \sa_snapshot[1][44] , 
	\sa_snapshot[1][43] , \sa_snapshot[1][42] , \sa_snapshot[1][41] , 
	\sa_snapshot[1][40] , \sa_snapshot[1][39] , \sa_snapshot[1][38] , 
	\sa_snapshot[1][37] , \sa_snapshot[1][36] , \sa_snapshot[1][35] , 
	\sa_snapshot[1][34] , \sa_snapshot[1][33] , \sa_snapshot[1][32] , 
	\sa_snapshot[1][31] , \sa_snapshot[1][30] , \sa_snapshot[1][29] , 
	\sa_snapshot[1][28] , \sa_snapshot[1][27] , \sa_snapshot[1][26] , 
	\sa_snapshot[1][25] , \sa_snapshot[1][24] , \sa_snapshot[1][23] , 
	\sa_snapshot[1][22] , \sa_snapshot[1][21] , \sa_snapshot[1][20] , 
	\sa_snapshot[1][19] , \sa_snapshot[1][18] , \sa_snapshot[1][17] , 
	\sa_snapshot[1][16] , \sa_snapshot[1][15] , \sa_snapshot[1][14] , 
	\sa_snapshot[1][13] , \sa_snapshot[1][12] , \sa_snapshot[1][11] , 
	\sa_snapshot[1][10] , \sa_snapshot[1][9] , \sa_snapshot[1][8] , 
	\sa_snapshot[1][7] , \sa_snapshot[1][6] , \sa_snapshot[1][5] , 
	\sa_snapshot[1][4] , \sa_snapshot[1][3] , \sa_snapshot[1][2] , 
	\sa_snapshot[1][1] , \sa_snapshot[1][0] , \sa_snapshot[0][63] , 
	\sa_snapshot[0][62] , \sa_snapshot[0][61] , \sa_snapshot[0][60] , 
	\sa_snapshot[0][59] , \sa_snapshot[0][58] , \sa_snapshot[0][57] , 
	\sa_snapshot[0][56] , \sa_snapshot[0][55] , \sa_snapshot[0][54] , 
	\sa_snapshot[0][53] , \sa_snapshot[0][52] , \sa_snapshot[0][51] , 
	\sa_snapshot[0][50] , \sa_snapshot[0][49] , \sa_snapshot[0][48] , 
	\sa_snapshot[0][47] , \sa_snapshot[0][46] , \sa_snapshot[0][45] , 
	\sa_snapshot[0][44] , \sa_snapshot[0][43] , \sa_snapshot[0][42] , 
	\sa_snapshot[0][41] , \sa_snapshot[0][40] , \sa_snapshot[0][39] , 
	\sa_snapshot[0][38] , \sa_snapshot[0][37] , \sa_snapshot[0][36] , 
	\sa_snapshot[0][35] , \sa_snapshot[0][34] , \sa_snapshot[0][33] , 
	\sa_snapshot[0][32] , \sa_snapshot[0][31] , \sa_snapshot[0][30] , 
	\sa_snapshot[0][29] , \sa_snapshot[0][28] , \sa_snapshot[0][27] , 
	\sa_snapshot[0][26] , \sa_snapshot[0][25] , \sa_snapshot[0][24] , 
	\sa_snapshot[0][23] , \sa_snapshot[0][22] , \sa_snapshot[0][21] , 
	\sa_snapshot[0][20] , \sa_snapshot[0][19] , \sa_snapshot[0][18] , 
	\sa_snapshot[0][17] , \sa_snapshot[0][16] , \sa_snapshot[0][15] , 
	\sa_snapshot[0][14] , \sa_snapshot[0][13] , \sa_snapshot[0][12] , 
	\sa_snapshot[0][11] , \sa_snapshot[0][10] , \sa_snapshot[0][9] , 
	\sa_snapshot[0][8] , \sa_snapshot[0][7] , \sa_snapshot[0][6] , 
	\sa_snapshot[0][5] , \sa_snapshot[0][4] , \sa_snapshot[0][3] , 
	\sa_snapshot[0][2] , \sa_snapshot[0][1] , \sa_snapshot[0][0] }), 
	.sa_count( { \sa_count[31][63] , \sa_count[31][62] , 
	\sa_count[31][61] , \sa_count[31][60] , \sa_count[31][59] , 
	\sa_count[31][58] , \sa_count[31][57] , \sa_count[31][56] , 
	\sa_count[31][55] , \sa_count[31][54] , \sa_count[31][53] , 
	\sa_count[31][52] , \sa_count[31][51] , \sa_count[31][50] , 
	\sa_count[31][49] , \sa_count[31][48] , \sa_count[31][47] , 
	\sa_count[31][46] , \sa_count[31][45] , \sa_count[31][44] , 
	\sa_count[31][43] , \sa_count[31][42] , \sa_count[31][41] , 
	\sa_count[31][40] , \sa_count[31][39] , \sa_count[31][38] , 
	\sa_count[31][37] , \sa_count[31][36] , \sa_count[31][35] , 
	\sa_count[31][34] , \sa_count[31][33] , \sa_count[31][32] , 
	\sa_count[31][31] , \sa_count[31][30] , \sa_count[31][29] , 
	\sa_count[31][28] , \sa_count[31][27] , \sa_count[31][26] , 
	\sa_count[31][25] , \sa_count[31][24] , \sa_count[31][23] , 
	\sa_count[31][22] , \sa_count[31][21] , \sa_count[31][20] , 
	\sa_count[31][19] , \sa_count[31][18] , \sa_count[31][17] , 
	\sa_count[31][16] , \sa_count[31][15] , \sa_count[31][14] , 
	\sa_count[31][13] , \sa_count[31][12] , \sa_count[31][11] , 
	\sa_count[31][10] , \sa_count[31][9] , \sa_count[31][8] , 
	\sa_count[31][7] , \sa_count[31][6] , \sa_count[31][5] , 
	\sa_count[31][4] , \sa_count[31][3] , \sa_count[31][2] , 
	\sa_count[31][1] , \sa_count[31][0] , \sa_count[30][63] , 
	\sa_count[30][62] , \sa_count[30][61] , \sa_count[30][60] , 
	\sa_count[30][59] , \sa_count[30][58] , \sa_count[30][57] , 
	\sa_count[30][56] , \sa_count[30][55] , \sa_count[30][54] , 
	\sa_count[30][53] , \sa_count[30][52] , \sa_count[30][51] , 
	\sa_count[30][50] , \sa_count[30][49] , \sa_count[30][48] , 
	\sa_count[30][47] , \sa_count[30][46] , \sa_count[30][45] , 
	\sa_count[30][44] , \sa_count[30][43] , \sa_count[30][42] , 
	\sa_count[30][41] , \sa_count[30][40] , \sa_count[30][39] , 
	\sa_count[30][38] , \sa_count[30][37] , \sa_count[30][36] , 
	\sa_count[30][35] , \sa_count[30][34] , \sa_count[30][33] , 
	\sa_count[30][32] , \sa_count[30][31] , \sa_count[30][30] , 
	\sa_count[30][29] , \sa_count[30][28] , \sa_count[30][27] , 
	\sa_count[30][26] , \sa_count[30][25] , \sa_count[30][24] , 
	\sa_count[30][23] , \sa_count[30][22] , \sa_count[30][21] , 
	\sa_count[30][20] , \sa_count[30][19] , \sa_count[30][18] , 
	\sa_count[30][17] , \sa_count[30][16] , \sa_count[30][15] , 
	\sa_count[30][14] , \sa_count[30][13] , \sa_count[30][12] , 
	\sa_count[30][11] , \sa_count[30][10] , \sa_count[30][9] , 
	\sa_count[30][8] , \sa_count[30][7] , \sa_count[30][6] , 
	\sa_count[30][5] , \sa_count[30][4] , \sa_count[30][3] , 
	\sa_count[30][2] , \sa_count[30][1] , \sa_count[30][0] , 
	\sa_count[29][63] , \sa_count[29][62] , \sa_count[29][61] , 
	\sa_count[29][60] , \sa_count[29][59] , \sa_count[29][58] , 
	\sa_count[29][57] , \sa_count[29][56] , \sa_count[29][55] , 
	\sa_count[29][54] , \sa_count[29][53] , \sa_count[29][52] , 
	\sa_count[29][51] , \sa_count[29][50] , \sa_count[29][49] , 
	\sa_count[29][48] , \sa_count[29][47] , \sa_count[29][46] , 
	\sa_count[29][45] , \sa_count[29][44] , \sa_count[29][43] , 
	\sa_count[29][42] , \sa_count[29][41] , \sa_count[29][40] , 
	\sa_count[29][39] , \sa_count[29][38] , \sa_count[29][37] , 
	\sa_count[29][36] , \sa_count[29][35] , \sa_count[29][34] , 
	\sa_count[29][33] , \sa_count[29][32] , \sa_count[29][31] , 
	\sa_count[29][30] , \sa_count[29][29] , \sa_count[29][28] , 
	\sa_count[29][27] , \sa_count[29][26] , \sa_count[29][25] , 
	\sa_count[29][24] , \sa_count[29][23] , \sa_count[29][22] , 
	\sa_count[29][21] , \sa_count[29][20] , \sa_count[29][19] , 
	\sa_count[29][18] , \sa_count[29][17] , \sa_count[29][16] , 
	\sa_count[29][15] , \sa_count[29][14] , \sa_count[29][13] , 
	\sa_count[29][12] , \sa_count[29][11] , \sa_count[29][10] , 
	\sa_count[29][9] , \sa_count[29][8] , \sa_count[29][7] , 
	\sa_count[29][6] , \sa_count[29][5] , \sa_count[29][4] , 
	\sa_count[29][3] , \sa_count[29][2] , \sa_count[29][1] , 
	\sa_count[29][0] , \sa_count[28][63] , \sa_count[28][62] , 
	\sa_count[28][61] , \sa_count[28][60] , \sa_count[28][59] , 
	\sa_count[28][58] , \sa_count[28][57] , \sa_count[28][56] , 
	\sa_count[28][55] , \sa_count[28][54] , \sa_count[28][53] , 
	\sa_count[28][52] , \sa_count[28][51] , \sa_count[28][50] , 
	\sa_count[28][49] , \sa_count[28][48] , \sa_count[28][47] , 
	\sa_count[28][46] , \sa_count[28][45] , \sa_count[28][44] , 
	\sa_count[28][43] , \sa_count[28][42] , \sa_count[28][41] , 
	\sa_count[28][40] , \sa_count[28][39] , \sa_count[28][38] , 
	\sa_count[28][37] , \sa_count[28][36] , \sa_count[28][35] , 
	\sa_count[28][34] , \sa_count[28][33] , \sa_count[28][32] , 
	\sa_count[28][31] , \sa_count[28][30] , \sa_count[28][29] , 
	\sa_count[28][28] , \sa_count[28][27] , \sa_count[28][26] , 
	\sa_count[28][25] , \sa_count[28][24] , \sa_count[28][23] , 
	\sa_count[28][22] , \sa_count[28][21] , \sa_count[28][20] , 
	\sa_count[28][19] , \sa_count[28][18] , \sa_count[28][17] , 
	\sa_count[28][16] , \sa_count[28][15] , \sa_count[28][14] , 
	\sa_count[28][13] , \sa_count[28][12] , \sa_count[28][11] , 
	\sa_count[28][10] , \sa_count[28][9] , \sa_count[28][8] , 
	\sa_count[28][7] , \sa_count[28][6] , \sa_count[28][5] , 
	\sa_count[28][4] , \sa_count[28][3] , \sa_count[28][2] , 
	\sa_count[28][1] , \sa_count[28][0] , \sa_count[27][63] , 
	\sa_count[27][62] , \sa_count[27][61] , \sa_count[27][60] , 
	\sa_count[27][59] , \sa_count[27][58] , \sa_count[27][57] , 
	\sa_count[27][56] , \sa_count[27][55] , \sa_count[27][54] , 
	\sa_count[27][53] , \sa_count[27][52] , \sa_count[27][51] , 
	\sa_count[27][50] , \sa_count[27][49] , \sa_count[27][48] , 
	\sa_count[27][47] , \sa_count[27][46] , \sa_count[27][45] , 
	\sa_count[27][44] , \sa_count[27][43] , \sa_count[27][42] , 
	\sa_count[27][41] , \sa_count[27][40] , \sa_count[27][39] , 
	\sa_count[27][38] , \sa_count[27][37] , \sa_count[27][36] , 
	\sa_count[27][35] , \sa_count[27][34] , \sa_count[27][33] , 
	\sa_count[27][32] , \sa_count[27][31] , \sa_count[27][30] , 
	\sa_count[27][29] , \sa_count[27][28] , \sa_count[27][27] , 
	\sa_count[27][26] , \sa_count[27][25] , \sa_count[27][24] , 
	\sa_count[27][23] , \sa_count[27][22] , \sa_count[27][21] , 
	\sa_count[27][20] , \sa_count[27][19] , \sa_count[27][18] , 
	\sa_count[27][17] , \sa_count[27][16] , \sa_count[27][15] , 
	\sa_count[27][14] , \sa_count[27][13] , \sa_count[27][12] , 
	\sa_count[27][11] , \sa_count[27][10] , \sa_count[27][9] , 
	\sa_count[27][8] , \sa_count[27][7] , \sa_count[27][6] , 
	\sa_count[27][5] , \sa_count[27][4] , \sa_count[27][3] , 
	\sa_count[27][2] , \sa_count[27][1] , \sa_count[27][0] , 
	\sa_count[26][63] , \sa_count[26][62] , \sa_count[26][61] , 
	\sa_count[26][60] , \sa_count[26][59] , \sa_count[26][58] , 
	\sa_count[26][57] , \sa_count[26][56] , \sa_count[26][55] , 
	\sa_count[26][54] , \sa_count[26][53] , \sa_count[26][52] , 
	\sa_count[26][51] , \sa_count[26][50] , \sa_count[26][49] , 
	\sa_count[26][48] , \sa_count[26][47] , \sa_count[26][46] , 
	\sa_count[26][45] , \sa_count[26][44] , \sa_count[26][43] , 
	\sa_count[26][42] , \sa_count[26][41] , \sa_count[26][40] , 
	\sa_count[26][39] , \sa_count[26][38] , \sa_count[26][37] , 
	\sa_count[26][36] , \sa_count[26][35] , \sa_count[26][34] , 
	\sa_count[26][33] , \sa_count[26][32] , \sa_count[26][31] , 
	\sa_count[26][30] , \sa_count[26][29] , \sa_count[26][28] , 
	\sa_count[26][27] , \sa_count[26][26] , \sa_count[26][25] , 
	\sa_count[26][24] , \sa_count[26][23] , \sa_count[26][22] , 
	\sa_count[26][21] , \sa_count[26][20] , \sa_count[26][19] , 
	\sa_count[26][18] , \sa_count[26][17] , \sa_count[26][16] , 
	\sa_count[26][15] , \sa_count[26][14] , \sa_count[26][13] , 
	\sa_count[26][12] , \sa_count[26][11] , \sa_count[26][10] , 
	\sa_count[26][9] , \sa_count[26][8] , \sa_count[26][7] , 
	\sa_count[26][6] , \sa_count[26][5] , \sa_count[26][4] , 
	\sa_count[26][3] , \sa_count[26][2] , \sa_count[26][1] , 
	\sa_count[26][0] , \sa_count[25][63] , \sa_count[25][62] , 
	\sa_count[25][61] , \sa_count[25][60] , \sa_count[25][59] , 
	\sa_count[25][58] , \sa_count[25][57] , \sa_count[25][56] , 
	\sa_count[25][55] , \sa_count[25][54] , \sa_count[25][53] , 
	\sa_count[25][52] , \sa_count[25][51] , \sa_count[25][50] , 
	\sa_count[25][49] , \sa_count[25][48] , \sa_count[25][47] , 
	\sa_count[25][46] , \sa_count[25][45] , \sa_count[25][44] , 
	\sa_count[25][43] , \sa_count[25][42] , \sa_count[25][41] , 
	\sa_count[25][40] , \sa_count[25][39] , \sa_count[25][38] , 
	\sa_count[25][37] , \sa_count[25][36] , \sa_count[25][35] , 
	\sa_count[25][34] , \sa_count[25][33] , \sa_count[25][32] , 
	\sa_count[25][31] , \sa_count[25][30] , \sa_count[25][29] , 
	\sa_count[25][28] , \sa_count[25][27] , \sa_count[25][26] , 
	\sa_count[25][25] , \sa_count[25][24] , \sa_count[25][23] , 
	\sa_count[25][22] , \sa_count[25][21] , \sa_count[25][20] , 
	\sa_count[25][19] , \sa_count[25][18] , \sa_count[25][17] , 
	\sa_count[25][16] , \sa_count[25][15] , \sa_count[25][14] , 
	\sa_count[25][13] , \sa_count[25][12] , \sa_count[25][11] , 
	\sa_count[25][10] , \sa_count[25][9] , \sa_count[25][8] , 
	\sa_count[25][7] , \sa_count[25][6] , \sa_count[25][5] , 
	\sa_count[25][4] , \sa_count[25][3] , \sa_count[25][2] , 
	\sa_count[25][1] , \sa_count[25][0] , \sa_count[24][63] , 
	\sa_count[24][62] , \sa_count[24][61] , \sa_count[24][60] , 
	\sa_count[24][59] , \sa_count[24][58] , \sa_count[24][57] , 
	\sa_count[24][56] , \sa_count[24][55] , \sa_count[24][54] , 
	\sa_count[24][53] , \sa_count[24][52] , \sa_count[24][51] , 
	\sa_count[24][50] , \sa_count[24][49] , \sa_count[24][48] , 
	\sa_count[24][47] , \sa_count[24][46] , \sa_count[24][45] , 
	\sa_count[24][44] , \sa_count[24][43] , \sa_count[24][42] , 
	\sa_count[24][41] , \sa_count[24][40] , \sa_count[24][39] , 
	\sa_count[24][38] , \sa_count[24][37] , \sa_count[24][36] , 
	\sa_count[24][35] , \sa_count[24][34] , \sa_count[24][33] , 
	\sa_count[24][32] , \sa_count[24][31] , \sa_count[24][30] , 
	\sa_count[24][29] , \sa_count[24][28] , \sa_count[24][27] , 
	\sa_count[24][26] , \sa_count[24][25] , \sa_count[24][24] , 
	\sa_count[24][23] , \sa_count[24][22] , \sa_count[24][21] , 
	\sa_count[24][20] , \sa_count[24][19] , \sa_count[24][18] , 
	\sa_count[24][17] , \sa_count[24][16] , \sa_count[24][15] , 
	\sa_count[24][14] , \sa_count[24][13] , \sa_count[24][12] , 
	\sa_count[24][11] , \sa_count[24][10] , \sa_count[24][9] , 
	\sa_count[24][8] , \sa_count[24][7] , \sa_count[24][6] , 
	\sa_count[24][5] , \sa_count[24][4] , \sa_count[24][3] , 
	\sa_count[24][2] , \sa_count[24][1] , \sa_count[24][0] , 
	\sa_count[23][63] , \sa_count[23][62] , \sa_count[23][61] , 
	\sa_count[23][60] , \sa_count[23][59] , \sa_count[23][58] , 
	\sa_count[23][57] , \sa_count[23][56] , \sa_count[23][55] , 
	\sa_count[23][54] , \sa_count[23][53] , \sa_count[23][52] , 
	\sa_count[23][51] , \sa_count[23][50] , \sa_count[23][49] , 
	\sa_count[23][48] , \sa_count[23][47] , \sa_count[23][46] , 
	\sa_count[23][45] , \sa_count[23][44] , \sa_count[23][43] , 
	\sa_count[23][42] , \sa_count[23][41] , \sa_count[23][40] , 
	\sa_count[23][39] , \sa_count[23][38] , \sa_count[23][37] , 
	\sa_count[23][36] , \sa_count[23][35] , \sa_count[23][34] , 
	\sa_count[23][33] , \sa_count[23][32] , \sa_count[23][31] , 
	\sa_count[23][30] , \sa_count[23][29] , \sa_count[23][28] , 
	\sa_count[23][27] , \sa_count[23][26] , \sa_count[23][25] , 
	\sa_count[23][24] , \sa_count[23][23] , \sa_count[23][22] , 
	\sa_count[23][21] , \sa_count[23][20] , \sa_count[23][19] , 
	\sa_count[23][18] , \sa_count[23][17] , \sa_count[23][16] , 
	\sa_count[23][15] , \sa_count[23][14] , \sa_count[23][13] , 
	\sa_count[23][12] , \sa_count[23][11] , \sa_count[23][10] , 
	\sa_count[23][9] , \sa_count[23][8] , \sa_count[23][7] , 
	\sa_count[23][6] , \sa_count[23][5] , \sa_count[23][4] , 
	\sa_count[23][3] , \sa_count[23][2] , \sa_count[23][1] , 
	\sa_count[23][0] , \sa_count[22][63] , \sa_count[22][62] , 
	\sa_count[22][61] , \sa_count[22][60] , \sa_count[22][59] , 
	\sa_count[22][58] , \sa_count[22][57] , \sa_count[22][56] , 
	\sa_count[22][55] , \sa_count[22][54] , \sa_count[22][53] , 
	\sa_count[22][52] , \sa_count[22][51] , \sa_count[22][50] , 
	\sa_count[22][49] , \sa_count[22][48] , \sa_count[22][47] , 
	\sa_count[22][46] , \sa_count[22][45] , \sa_count[22][44] , 
	\sa_count[22][43] , \sa_count[22][42] , \sa_count[22][41] , 
	\sa_count[22][40] , \sa_count[22][39] , \sa_count[22][38] , 
	\sa_count[22][37] , \sa_count[22][36] , \sa_count[22][35] , 
	\sa_count[22][34] , \sa_count[22][33] , \sa_count[22][32] , 
	\sa_count[22][31] , \sa_count[22][30] , \sa_count[22][29] , 
	\sa_count[22][28] , \sa_count[22][27] , \sa_count[22][26] , 
	\sa_count[22][25] , \sa_count[22][24] , \sa_count[22][23] , 
	\sa_count[22][22] , \sa_count[22][21] , \sa_count[22][20] , 
	\sa_count[22][19] , \sa_count[22][18] , \sa_count[22][17] , 
	\sa_count[22][16] , \sa_count[22][15] , \sa_count[22][14] , 
	\sa_count[22][13] , \sa_count[22][12] , \sa_count[22][11] , 
	\sa_count[22][10] , \sa_count[22][9] , \sa_count[22][8] , 
	\sa_count[22][7] , \sa_count[22][6] , \sa_count[22][5] , 
	\sa_count[22][4] , \sa_count[22][3] , \sa_count[22][2] , 
	\sa_count[22][1] , \sa_count[22][0] , \sa_count[21][63] , 
	\sa_count[21][62] , \sa_count[21][61] , \sa_count[21][60] , 
	\sa_count[21][59] , \sa_count[21][58] , \sa_count[21][57] , 
	\sa_count[21][56] , \sa_count[21][55] , \sa_count[21][54] , 
	\sa_count[21][53] , \sa_count[21][52] , \sa_count[21][51] , 
	\sa_count[21][50] , \sa_count[21][49] , \sa_count[21][48] , 
	\sa_count[21][47] , \sa_count[21][46] , \sa_count[21][45] , 
	\sa_count[21][44] , \sa_count[21][43] , \sa_count[21][42] , 
	\sa_count[21][41] , \sa_count[21][40] , \sa_count[21][39] , 
	\sa_count[21][38] , \sa_count[21][37] , \sa_count[21][36] , 
	\sa_count[21][35] , \sa_count[21][34] , \sa_count[21][33] , 
	\sa_count[21][32] , \sa_count[21][31] , \sa_count[21][30] , 
	\sa_count[21][29] , \sa_count[21][28] , \sa_count[21][27] , 
	\sa_count[21][26] , \sa_count[21][25] , \sa_count[21][24] , 
	\sa_count[21][23] , \sa_count[21][22] , \sa_count[21][21] , 
	\sa_count[21][20] , \sa_count[21][19] , \sa_count[21][18] , 
	\sa_count[21][17] , \sa_count[21][16] , \sa_count[21][15] , 
	\sa_count[21][14] , \sa_count[21][13] , \sa_count[21][12] , 
	\sa_count[21][11] , \sa_count[21][10] , \sa_count[21][9] , 
	\sa_count[21][8] , \sa_count[21][7] , \sa_count[21][6] , 
	\sa_count[21][5] , \sa_count[21][4] , \sa_count[21][3] , 
	\sa_count[21][2] , \sa_count[21][1] , \sa_count[21][0] , 
	\sa_count[20][63] , \sa_count[20][62] , \sa_count[20][61] , 
	\sa_count[20][60] , \sa_count[20][59] , \sa_count[20][58] , 
	\sa_count[20][57] , \sa_count[20][56] , \sa_count[20][55] , 
	\sa_count[20][54] , \sa_count[20][53] , \sa_count[20][52] , 
	\sa_count[20][51] , \sa_count[20][50] , \sa_count[20][49] , 
	\sa_count[20][48] , \sa_count[20][47] , \sa_count[20][46] , 
	\sa_count[20][45] , \sa_count[20][44] , \sa_count[20][43] , 
	\sa_count[20][42] , \sa_count[20][41] , \sa_count[20][40] , 
	\sa_count[20][39] , \sa_count[20][38] , \sa_count[20][37] , 
	\sa_count[20][36] , \sa_count[20][35] , \sa_count[20][34] , 
	\sa_count[20][33] , \sa_count[20][32] , \sa_count[20][31] , 
	\sa_count[20][30] , \sa_count[20][29] , \sa_count[20][28] , 
	\sa_count[20][27] , \sa_count[20][26] , \sa_count[20][25] , 
	\sa_count[20][24] , \sa_count[20][23] , \sa_count[20][22] , 
	\sa_count[20][21] , \sa_count[20][20] , \sa_count[20][19] , 
	\sa_count[20][18] , \sa_count[20][17] , \sa_count[20][16] , 
	\sa_count[20][15] , \sa_count[20][14] , \sa_count[20][13] , 
	\sa_count[20][12] , \sa_count[20][11] , \sa_count[20][10] , 
	\sa_count[20][9] , \sa_count[20][8] , \sa_count[20][7] , 
	\sa_count[20][6] , \sa_count[20][5] , \sa_count[20][4] , 
	\sa_count[20][3] , \sa_count[20][2] , \sa_count[20][1] , 
	\sa_count[20][0] , \sa_count[19][63] , \sa_count[19][62] , 
	\sa_count[19][61] , \sa_count[19][60] , \sa_count[19][59] , 
	\sa_count[19][58] , \sa_count[19][57] , \sa_count[19][56] , 
	\sa_count[19][55] , \sa_count[19][54] , \sa_count[19][53] , 
	\sa_count[19][52] , \sa_count[19][51] , \sa_count[19][50] , 
	\sa_count[19][49] , \sa_count[19][48] , \sa_count[19][47] , 
	\sa_count[19][46] , \sa_count[19][45] , \sa_count[19][44] , 
	\sa_count[19][43] , \sa_count[19][42] , \sa_count[19][41] , 
	\sa_count[19][40] , \sa_count[19][39] , \sa_count[19][38] , 
	\sa_count[19][37] , \sa_count[19][36] , \sa_count[19][35] , 
	\sa_count[19][34] , \sa_count[19][33] , \sa_count[19][32] , 
	\sa_count[19][31] , \sa_count[19][30] , \sa_count[19][29] , 
	\sa_count[19][28] , \sa_count[19][27] , \sa_count[19][26] , 
	\sa_count[19][25] , \sa_count[19][24] , \sa_count[19][23] , 
	\sa_count[19][22] , \sa_count[19][21] , \sa_count[19][20] , 
	\sa_count[19][19] , \sa_count[19][18] , \sa_count[19][17] , 
	\sa_count[19][16] , \sa_count[19][15] , \sa_count[19][14] , 
	\sa_count[19][13] , \sa_count[19][12] , \sa_count[19][11] , 
	\sa_count[19][10] , \sa_count[19][9] , \sa_count[19][8] , 
	\sa_count[19][7] , \sa_count[19][6] , \sa_count[19][5] , 
	\sa_count[19][4] , \sa_count[19][3] , \sa_count[19][2] , 
	\sa_count[19][1] , \sa_count[19][0] , \sa_count[18][63] , 
	\sa_count[18][62] , \sa_count[18][61] , \sa_count[18][60] , 
	\sa_count[18][59] , \sa_count[18][58] , \sa_count[18][57] , 
	\sa_count[18][56] , \sa_count[18][55] , \sa_count[18][54] , 
	\sa_count[18][53] , \sa_count[18][52] , \sa_count[18][51] , 
	\sa_count[18][50] , \sa_count[18][49] , \sa_count[18][48] , 
	\sa_count[18][47] , \sa_count[18][46] , \sa_count[18][45] , 
	\sa_count[18][44] , \sa_count[18][43] , \sa_count[18][42] , 
	\sa_count[18][41] , \sa_count[18][40] , \sa_count[18][39] , 
	\sa_count[18][38] , \sa_count[18][37] , \sa_count[18][36] , 
	\sa_count[18][35] , \sa_count[18][34] , \sa_count[18][33] , 
	\sa_count[18][32] , \sa_count[18][31] , \sa_count[18][30] , 
	\sa_count[18][29] , \sa_count[18][28] , \sa_count[18][27] , 
	\sa_count[18][26] , \sa_count[18][25] , \sa_count[18][24] , 
	\sa_count[18][23] , \sa_count[18][22] , \sa_count[18][21] , 
	\sa_count[18][20] , \sa_count[18][19] , \sa_count[18][18] , 
	\sa_count[18][17] , \sa_count[18][16] , \sa_count[18][15] , 
	\sa_count[18][14] , \sa_count[18][13] , \sa_count[18][12] , 
	\sa_count[18][11] , \sa_count[18][10] , \sa_count[18][9] , 
	\sa_count[18][8] , \sa_count[18][7] , \sa_count[18][6] , 
	\sa_count[18][5] , \sa_count[18][4] , \sa_count[18][3] , 
	\sa_count[18][2] , \sa_count[18][1] , \sa_count[18][0] , 
	\sa_count[17][63] , \sa_count[17][62] , \sa_count[17][61] , 
	\sa_count[17][60] , \sa_count[17][59] , \sa_count[17][58] , 
	\sa_count[17][57] , \sa_count[17][56] , \sa_count[17][55] , 
	\sa_count[17][54] , \sa_count[17][53] , \sa_count[17][52] , 
	\sa_count[17][51] , \sa_count[17][50] , \sa_count[17][49] , 
	\sa_count[17][48] , \sa_count[17][47] , \sa_count[17][46] , 
	\sa_count[17][45] , \sa_count[17][44] , \sa_count[17][43] , 
	\sa_count[17][42] , \sa_count[17][41] , \sa_count[17][40] , 
	\sa_count[17][39] , \sa_count[17][38] , \sa_count[17][37] , 
	\sa_count[17][36] , \sa_count[17][35] , \sa_count[17][34] , 
	\sa_count[17][33] , \sa_count[17][32] , \sa_count[17][31] , 
	\sa_count[17][30] , \sa_count[17][29] , \sa_count[17][28] , 
	\sa_count[17][27] , \sa_count[17][26] , \sa_count[17][25] , 
	\sa_count[17][24] , \sa_count[17][23] , \sa_count[17][22] , 
	\sa_count[17][21] , \sa_count[17][20] , \sa_count[17][19] , 
	\sa_count[17][18] , \sa_count[17][17] , \sa_count[17][16] , 
	\sa_count[17][15] , \sa_count[17][14] , \sa_count[17][13] , 
	\sa_count[17][12] , \sa_count[17][11] , \sa_count[17][10] , 
	\sa_count[17][9] , \sa_count[17][8] , \sa_count[17][7] , 
	\sa_count[17][6] , \sa_count[17][5] , \sa_count[17][4] , 
	\sa_count[17][3] , \sa_count[17][2] , \sa_count[17][1] , 
	\sa_count[17][0] , \sa_count[16][63] , \sa_count[16][62] , 
	\sa_count[16][61] , \sa_count[16][60] , \sa_count[16][59] , 
	\sa_count[16][58] , \sa_count[16][57] , \sa_count[16][56] , 
	\sa_count[16][55] , \sa_count[16][54] , \sa_count[16][53] , 
	\sa_count[16][52] , \sa_count[16][51] , \sa_count[16][50] , 
	\sa_count[16][49] , \sa_count[16][48] , \sa_count[16][47] , 
	\sa_count[16][46] , \sa_count[16][45] , \sa_count[16][44] , 
	\sa_count[16][43] , \sa_count[16][42] , \sa_count[16][41] , 
	\sa_count[16][40] , \sa_count[16][39] , \sa_count[16][38] , 
	\sa_count[16][37] , \sa_count[16][36] , \sa_count[16][35] , 
	\sa_count[16][34] , \sa_count[16][33] , \sa_count[16][32] , 
	\sa_count[16][31] , \sa_count[16][30] , \sa_count[16][29] , 
	\sa_count[16][28] , \sa_count[16][27] , \sa_count[16][26] , 
	\sa_count[16][25] , \sa_count[16][24] , \sa_count[16][23] , 
	\sa_count[16][22] , \sa_count[16][21] , \sa_count[16][20] , 
	\sa_count[16][19] , \sa_count[16][18] , \sa_count[16][17] , 
	\sa_count[16][16] , \sa_count[16][15] , \sa_count[16][14] , 
	\sa_count[16][13] , \sa_count[16][12] , \sa_count[16][11] , 
	\sa_count[16][10] , \sa_count[16][9] , \sa_count[16][8] , 
	\sa_count[16][7] , \sa_count[16][6] , \sa_count[16][5] , 
	\sa_count[16][4] , \sa_count[16][3] , \sa_count[16][2] , 
	\sa_count[16][1] , \sa_count[16][0] , \sa_count[15][63] , 
	\sa_count[15][62] , \sa_count[15][61] , \sa_count[15][60] , 
	\sa_count[15][59] , \sa_count[15][58] , \sa_count[15][57] , 
	\sa_count[15][56] , \sa_count[15][55] , \sa_count[15][54] , 
	\sa_count[15][53] , \sa_count[15][52] , \sa_count[15][51] , 
	\sa_count[15][50] , \sa_count[15][49] , \sa_count[15][48] , 
	\sa_count[15][47] , \sa_count[15][46] , \sa_count[15][45] , 
	\sa_count[15][44] , \sa_count[15][43] , \sa_count[15][42] , 
	\sa_count[15][41] , \sa_count[15][40] , \sa_count[15][39] , 
	\sa_count[15][38] , \sa_count[15][37] , \sa_count[15][36] , 
	\sa_count[15][35] , \sa_count[15][34] , \sa_count[15][33] , 
	\sa_count[15][32] , \sa_count[15][31] , \sa_count[15][30] , 
	\sa_count[15][29] , \sa_count[15][28] , \sa_count[15][27] , 
	\sa_count[15][26] , \sa_count[15][25] , \sa_count[15][24] , 
	\sa_count[15][23] , \sa_count[15][22] , \sa_count[15][21] , 
	\sa_count[15][20] , \sa_count[15][19] , \sa_count[15][18] , 
	\sa_count[15][17] , \sa_count[15][16] , \sa_count[15][15] , 
	\sa_count[15][14] , \sa_count[15][13] , \sa_count[15][12] , 
	\sa_count[15][11] , \sa_count[15][10] , \sa_count[15][9] , 
	\sa_count[15][8] , \sa_count[15][7] , \sa_count[15][6] , 
	\sa_count[15][5] , \sa_count[15][4] , \sa_count[15][3] , 
	\sa_count[15][2] , \sa_count[15][1] , \sa_count[15][0] , 
	\sa_count[14][63] , \sa_count[14][62] , \sa_count[14][61] , 
	\sa_count[14][60] , \sa_count[14][59] , \sa_count[14][58] , 
	\sa_count[14][57] , \sa_count[14][56] , \sa_count[14][55] , 
	\sa_count[14][54] , \sa_count[14][53] , \sa_count[14][52] , 
	\sa_count[14][51] , \sa_count[14][50] , \sa_count[14][49] , 
	\sa_count[14][48] , \sa_count[14][47] , \sa_count[14][46] , 
	\sa_count[14][45] , \sa_count[14][44] , \sa_count[14][43] , 
	\sa_count[14][42] , \sa_count[14][41] , \sa_count[14][40] , 
	\sa_count[14][39] , \sa_count[14][38] , \sa_count[14][37] , 
	\sa_count[14][36] , \sa_count[14][35] , \sa_count[14][34] , 
	\sa_count[14][33] , \sa_count[14][32] , \sa_count[14][31] , 
	\sa_count[14][30] , \sa_count[14][29] , \sa_count[14][28] , 
	\sa_count[14][27] , \sa_count[14][26] , \sa_count[14][25] , 
	\sa_count[14][24] , \sa_count[14][23] , \sa_count[14][22] , 
	\sa_count[14][21] , \sa_count[14][20] , \sa_count[14][19] , 
	\sa_count[14][18] , \sa_count[14][17] , \sa_count[14][16] , 
	\sa_count[14][15] , \sa_count[14][14] , \sa_count[14][13] , 
	\sa_count[14][12] , \sa_count[14][11] , \sa_count[14][10] , 
	\sa_count[14][9] , \sa_count[14][8] , \sa_count[14][7] , 
	\sa_count[14][6] , \sa_count[14][5] , \sa_count[14][4] , 
	\sa_count[14][3] , \sa_count[14][2] , \sa_count[14][1] , 
	\sa_count[14][0] , \sa_count[13][63] , \sa_count[13][62] , 
	\sa_count[13][61] , \sa_count[13][60] , \sa_count[13][59] , 
	\sa_count[13][58] , \sa_count[13][57] , \sa_count[13][56] , 
	\sa_count[13][55] , \sa_count[13][54] , \sa_count[13][53] , 
	\sa_count[13][52] , \sa_count[13][51] , \sa_count[13][50] , 
	\sa_count[13][49] , \sa_count[13][48] , \sa_count[13][47] , 
	\sa_count[13][46] , \sa_count[13][45] , \sa_count[13][44] , 
	\sa_count[13][43] , \sa_count[13][42] , \sa_count[13][41] , 
	\sa_count[13][40] , \sa_count[13][39] , \sa_count[13][38] , 
	\sa_count[13][37] , \sa_count[13][36] , \sa_count[13][35] , 
	\sa_count[13][34] , \sa_count[13][33] , \sa_count[13][32] , 
	\sa_count[13][31] , \sa_count[13][30] , \sa_count[13][29] , 
	\sa_count[13][28] , \sa_count[13][27] , \sa_count[13][26] , 
	\sa_count[13][25] , \sa_count[13][24] , \sa_count[13][23] , 
	\sa_count[13][22] , \sa_count[13][21] , \sa_count[13][20] , 
	\sa_count[13][19] , \sa_count[13][18] , \sa_count[13][17] , 
	\sa_count[13][16] , \sa_count[13][15] , \sa_count[13][14] , 
	\sa_count[13][13] , \sa_count[13][12] , \sa_count[13][11] , 
	\sa_count[13][10] , \sa_count[13][9] , \sa_count[13][8] , 
	\sa_count[13][7] , \sa_count[13][6] , \sa_count[13][5] , 
	\sa_count[13][4] , \sa_count[13][3] , \sa_count[13][2] , 
	\sa_count[13][1] , \sa_count[13][0] , \sa_count[12][63] , 
	\sa_count[12][62] , \sa_count[12][61] , \sa_count[12][60] , 
	\sa_count[12][59] , \sa_count[12][58] , \sa_count[12][57] , 
	\sa_count[12][56] , \sa_count[12][55] , \sa_count[12][54] , 
	\sa_count[12][53] , \sa_count[12][52] , \sa_count[12][51] , 
	\sa_count[12][50] , \sa_count[12][49] , \sa_count[12][48] , 
	\sa_count[12][47] , \sa_count[12][46] , \sa_count[12][45] , 
	\sa_count[12][44] , \sa_count[12][43] , \sa_count[12][42] , 
	\sa_count[12][41] , \sa_count[12][40] , \sa_count[12][39] , 
	\sa_count[12][38] , \sa_count[12][37] , \sa_count[12][36] , 
	\sa_count[12][35] , \sa_count[12][34] , \sa_count[12][33] , 
	\sa_count[12][32] , \sa_count[12][31] , \sa_count[12][30] , 
	\sa_count[12][29] , \sa_count[12][28] , \sa_count[12][27] , 
	\sa_count[12][26] , \sa_count[12][25] , \sa_count[12][24] , 
	\sa_count[12][23] , \sa_count[12][22] , \sa_count[12][21] , 
	\sa_count[12][20] , \sa_count[12][19] , \sa_count[12][18] , 
	\sa_count[12][17] , \sa_count[12][16] , \sa_count[12][15] , 
	\sa_count[12][14] , \sa_count[12][13] , \sa_count[12][12] , 
	\sa_count[12][11] , \sa_count[12][10] , \sa_count[12][9] , 
	\sa_count[12][8] , \sa_count[12][7] , \sa_count[12][6] , 
	\sa_count[12][5] , \sa_count[12][4] , \sa_count[12][3] , 
	\sa_count[12][2] , \sa_count[12][1] , \sa_count[12][0] , 
	\sa_count[11][63] , \sa_count[11][62] , \sa_count[11][61] , 
	\sa_count[11][60] , \sa_count[11][59] , \sa_count[11][58] , 
	\sa_count[11][57] , \sa_count[11][56] , \sa_count[11][55] , 
	\sa_count[11][54] , \sa_count[11][53] , \sa_count[11][52] , 
	\sa_count[11][51] , \sa_count[11][50] , \sa_count[11][49] , 
	\sa_count[11][48] , \sa_count[11][47] , \sa_count[11][46] , 
	\sa_count[11][45] , \sa_count[11][44] , \sa_count[11][43] , 
	\sa_count[11][42] , \sa_count[11][41] , \sa_count[11][40] , 
	\sa_count[11][39] , \sa_count[11][38] , \sa_count[11][37] , 
	\sa_count[11][36] , \sa_count[11][35] , \sa_count[11][34] , 
	\sa_count[11][33] , \sa_count[11][32] , \sa_count[11][31] , 
	\sa_count[11][30] , \sa_count[11][29] , \sa_count[11][28] , 
	\sa_count[11][27] , \sa_count[11][26] , \sa_count[11][25] , 
	\sa_count[11][24] , \sa_count[11][23] , \sa_count[11][22] , 
	\sa_count[11][21] , \sa_count[11][20] , \sa_count[11][19] , 
	\sa_count[11][18] , \sa_count[11][17] , \sa_count[11][16] , 
	\sa_count[11][15] , \sa_count[11][14] , \sa_count[11][13] , 
	\sa_count[11][12] , \sa_count[11][11] , \sa_count[11][10] , 
	\sa_count[11][9] , \sa_count[11][8] , \sa_count[11][7] , 
	\sa_count[11][6] , \sa_count[11][5] , \sa_count[11][4] , 
	\sa_count[11][3] , \sa_count[11][2] , \sa_count[11][1] , 
	\sa_count[11][0] , \sa_count[10][63] , \sa_count[10][62] , 
	\sa_count[10][61] , \sa_count[10][60] , \sa_count[10][59] , 
	\sa_count[10][58] , \sa_count[10][57] , \sa_count[10][56] , 
	\sa_count[10][55] , \sa_count[10][54] , \sa_count[10][53] , 
	\sa_count[10][52] , \sa_count[10][51] , \sa_count[10][50] , 
	\sa_count[10][49] , \sa_count[10][48] , \sa_count[10][47] , 
	\sa_count[10][46] , \sa_count[10][45] , \sa_count[10][44] , 
	\sa_count[10][43] , \sa_count[10][42] , \sa_count[10][41] , 
	\sa_count[10][40] , \sa_count[10][39] , \sa_count[10][38] , 
	\sa_count[10][37] , \sa_count[10][36] , \sa_count[10][35] , 
	\sa_count[10][34] , \sa_count[10][33] , \sa_count[10][32] , 
	\sa_count[10][31] , \sa_count[10][30] , \sa_count[10][29] , 
	\sa_count[10][28] , \sa_count[10][27] , \sa_count[10][26] , 
	\sa_count[10][25] , \sa_count[10][24] , \sa_count[10][23] , 
	\sa_count[10][22] , \sa_count[10][21] , \sa_count[10][20] , 
	\sa_count[10][19] , \sa_count[10][18] , \sa_count[10][17] , 
	\sa_count[10][16] , \sa_count[10][15] , \sa_count[10][14] , 
	\sa_count[10][13] , \sa_count[10][12] , \sa_count[10][11] , 
	\sa_count[10][10] , \sa_count[10][9] , \sa_count[10][8] , 
	\sa_count[10][7] , \sa_count[10][6] , \sa_count[10][5] , 
	\sa_count[10][4] , \sa_count[10][3] , \sa_count[10][2] , 
	\sa_count[10][1] , \sa_count[10][0] , \sa_count[9][63] , 
	\sa_count[9][62] , \sa_count[9][61] , \sa_count[9][60] , 
	\sa_count[9][59] , \sa_count[9][58] , \sa_count[9][57] , 
	\sa_count[9][56] , \sa_count[9][55] , \sa_count[9][54] , 
	\sa_count[9][53] , \sa_count[9][52] , \sa_count[9][51] , 
	\sa_count[9][50] , \sa_count[9][49] , \sa_count[9][48] , 
	\sa_count[9][47] , \sa_count[9][46] , \sa_count[9][45] , 
	\sa_count[9][44] , \sa_count[9][43] , \sa_count[9][42] , 
	\sa_count[9][41] , \sa_count[9][40] , \sa_count[9][39] , 
	\sa_count[9][38] , \sa_count[9][37] , \sa_count[9][36] , 
	\sa_count[9][35] , \sa_count[9][34] , \sa_count[9][33] , 
	\sa_count[9][32] , \sa_count[9][31] , \sa_count[9][30] , 
	\sa_count[9][29] , \sa_count[9][28] , \sa_count[9][27] , 
	\sa_count[9][26] , \sa_count[9][25] , \sa_count[9][24] , 
	\sa_count[9][23] , \sa_count[9][22] , \sa_count[9][21] , 
	\sa_count[9][20] , \sa_count[9][19] , \sa_count[9][18] , 
	\sa_count[9][17] , \sa_count[9][16] , \sa_count[9][15] , 
	\sa_count[9][14] , \sa_count[9][13] , \sa_count[9][12] , 
	\sa_count[9][11] , \sa_count[9][10] , \sa_count[9][9] , 
	\sa_count[9][8] , \sa_count[9][7] , \sa_count[9][6] , 
	\sa_count[9][5] , \sa_count[9][4] , \sa_count[9][3] , 
	\sa_count[9][2] , \sa_count[9][1] , \sa_count[9][0] , 
	\sa_count[8][63] , \sa_count[8][62] , \sa_count[8][61] , 
	\sa_count[8][60] , \sa_count[8][59] , \sa_count[8][58] , 
	\sa_count[8][57] , \sa_count[8][56] , \sa_count[8][55] , 
	\sa_count[8][54] , \sa_count[8][53] , \sa_count[8][52] , 
	\sa_count[8][51] , \sa_count[8][50] , \sa_count[8][49] , 
	\sa_count[8][48] , \sa_count[8][47] , \sa_count[8][46] , 
	\sa_count[8][45] , \sa_count[8][44] , \sa_count[8][43] , 
	\sa_count[8][42] , \sa_count[8][41] , \sa_count[8][40] , 
	\sa_count[8][39] , \sa_count[8][38] , \sa_count[8][37] , 
	\sa_count[8][36] , \sa_count[8][35] , \sa_count[8][34] , 
	\sa_count[8][33] , \sa_count[8][32] , \sa_count[8][31] , 
	\sa_count[8][30] , \sa_count[8][29] , \sa_count[8][28] , 
	\sa_count[8][27] , \sa_count[8][26] , \sa_count[8][25] , 
	\sa_count[8][24] , \sa_count[8][23] , \sa_count[8][22] , 
	\sa_count[8][21] , \sa_count[8][20] , \sa_count[8][19] , 
	\sa_count[8][18] , \sa_count[8][17] , \sa_count[8][16] , 
	\sa_count[8][15] , \sa_count[8][14] , \sa_count[8][13] , 
	\sa_count[8][12] , \sa_count[8][11] , \sa_count[8][10] , 
	\sa_count[8][9] , \sa_count[8][8] , \sa_count[8][7] , 
	\sa_count[8][6] , \sa_count[8][5] , \sa_count[8][4] , 
	\sa_count[8][3] , \sa_count[8][2] , \sa_count[8][1] , 
	\sa_count[8][0] , \sa_count[7][63] , \sa_count[7][62] , 
	\sa_count[7][61] , \sa_count[7][60] , \sa_count[7][59] , 
	\sa_count[7][58] , \sa_count[7][57] , \sa_count[7][56] , 
	\sa_count[7][55] , \sa_count[7][54] , \sa_count[7][53] , 
	\sa_count[7][52] , \sa_count[7][51] , \sa_count[7][50] , 
	\sa_count[7][49] , \sa_count[7][48] , \sa_count[7][47] , 
	\sa_count[7][46] , \sa_count[7][45] , \sa_count[7][44] , 
	\sa_count[7][43] , \sa_count[7][42] , \sa_count[7][41] , 
	\sa_count[7][40] , \sa_count[7][39] , \sa_count[7][38] , 
	\sa_count[7][37] , \sa_count[7][36] , \sa_count[7][35] , 
	\sa_count[7][34] , \sa_count[7][33] , \sa_count[7][32] , 
	\sa_count[7][31] , \sa_count[7][30] , \sa_count[7][29] , 
	\sa_count[7][28] , \sa_count[7][27] , \sa_count[7][26] , 
	\sa_count[7][25] , \sa_count[7][24] , \sa_count[7][23] , 
	\sa_count[7][22] , \sa_count[7][21] , \sa_count[7][20] , 
	\sa_count[7][19] , \sa_count[7][18] , \sa_count[7][17] , 
	\sa_count[7][16] , \sa_count[7][15] , \sa_count[7][14] , 
	\sa_count[7][13] , \sa_count[7][12] , \sa_count[7][11] , 
	\sa_count[7][10] , \sa_count[7][9] , \sa_count[7][8] , 
	\sa_count[7][7] , \sa_count[7][6] , \sa_count[7][5] , 
	\sa_count[7][4] , \sa_count[7][3] , \sa_count[7][2] , 
	\sa_count[7][1] , \sa_count[7][0] , \sa_count[6][63] , 
	\sa_count[6][62] , \sa_count[6][61] , \sa_count[6][60] , 
	\sa_count[6][59] , \sa_count[6][58] , \sa_count[6][57] , 
	\sa_count[6][56] , \sa_count[6][55] , \sa_count[6][54] , 
	\sa_count[6][53] , \sa_count[6][52] , \sa_count[6][51] , 
	\sa_count[6][50] , \sa_count[6][49] , \sa_count[6][48] , 
	\sa_count[6][47] , \sa_count[6][46] , \sa_count[6][45] , 
	\sa_count[6][44] , \sa_count[6][43] , \sa_count[6][42] , 
	\sa_count[6][41] , \sa_count[6][40] , \sa_count[6][39] , 
	\sa_count[6][38] , \sa_count[6][37] , \sa_count[6][36] , 
	\sa_count[6][35] , \sa_count[6][34] , \sa_count[6][33] , 
	\sa_count[6][32] , \sa_count[6][31] , \sa_count[6][30] , 
	\sa_count[6][29] , \sa_count[6][28] , \sa_count[6][27] , 
	\sa_count[6][26] , \sa_count[6][25] , \sa_count[6][24] , 
	\sa_count[6][23] , \sa_count[6][22] , \sa_count[6][21] , 
	\sa_count[6][20] , \sa_count[6][19] , \sa_count[6][18] , 
	\sa_count[6][17] , \sa_count[6][16] , \sa_count[6][15] , 
	\sa_count[6][14] , \sa_count[6][13] , \sa_count[6][12] , 
	\sa_count[6][11] , \sa_count[6][10] , \sa_count[6][9] , 
	\sa_count[6][8] , \sa_count[6][7] , \sa_count[6][6] , 
	\sa_count[6][5] , \sa_count[6][4] , \sa_count[6][3] , 
	\sa_count[6][2] , \sa_count[6][1] , \sa_count[6][0] , 
	\sa_count[5][63] , \sa_count[5][62] , \sa_count[5][61] , 
	\sa_count[5][60] , \sa_count[5][59] , \sa_count[5][58] , 
	\sa_count[5][57] , \sa_count[5][56] , \sa_count[5][55] , 
	\sa_count[5][54] , \sa_count[5][53] , \sa_count[5][52] , 
	\sa_count[5][51] , \sa_count[5][50] , \sa_count[5][49] , 
	\sa_count[5][48] , \sa_count[5][47] , \sa_count[5][46] , 
	\sa_count[5][45] , \sa_count[5][44] , \sa_count[5][43] , 
	\sa_count[5][42] , \sa_count[5][41] , \sa_count[5][40] , 
	\sa_count[5][39] , \sa_count[5][38] , \sa_count[5][37] , 
	\sa_count[5][36] , \sa_count[5][35] , \sa_count[5][34] , 
	\sa_count[5][33] , \sa_count[5][32] , \sa_count[5][31] , 
	\sa_count[5][30] , \sa_count[5][29] , \sa_count[5][28] , 
	\sa_count[5][27] , \sa_count[5][26] , \sa_count[5][25] , 
	\sa_count[5][24] , \sa_count[5][23] , \sa_count[5][22] , 
	\sa_count[5][21] , \sa_count[5][20] , \sa_count[5][19] , 
	\sa_count[5][18] , \sa_count[5][17] , \sa_count[5][16] , 
	\sa_count[5][15] , \sa_count[5][14] , \sa_count[5][13] , 
	\sa_count[5][12] , \sa_count[5][11] , \sa_count[5][10] , 
	\sa_count[5][9] , \sa_count[5][8] , \sa_count[5][7] , 
	\sa_count[5][6] , \sa_count[5][5] , \sa_count[5][4] , 
	\sa_count[5][3] , \sa_count[5][2] , \sa_count[5][1] , 
	\sa_count[5][0] , \sa_count[4][63] , \sa_count[4][62] , 
	\sa_count[4][61] , \sa_count[4][60] , \sa_count[4][59] , 
	\sa_count[4][58] , \sa_count[4][57] , \sa_count[4][56] , 
	\sa_count[4][55] , \sa_count[4][54] , \sa_count[4][53] , 
	\sa_count[4][52] , \sa_count[4][51] , \sa_count[4][50] , 
	\sa_count[4][49] , \sa_count[4][48] , \sa_count[4][47] , 
	\sa_count[4][46] , \sa_count[4][45] , \sa_count[4][44] , 
	\sa_count[4][43] , \sa_count[4][42] , \sa_count[4][41] , 
	\sa_count[4][40] , \sa_count[4][39] , \sa_count[4][38] , 
	\sa_count[4][37] , \sa_count[4][36] , \sa_count[4][35] , 
	\sa_count[4][34] , \sa_count[4][33] , \sa_count[4][32] , 
	\sa_count[4][31] , \sa_count[4][30] , \sa_count[4][29] , 
	\sa_count[4][28] , \sa_count[4][27] , \sa_count[4][26] , 
	\sa_count[4][25] , \sa_count[4][24] , \sa_count[4][23] , 
	\sa_count[4][22] , \sa_count[4][21] , \sa_count[4][20] , 
	\sa_count[4][19] , \sa_count[4][18] , \sa_count[4][17] , 
	\sa_count[4][16] , \sa_count[4][15] , \sa_count[4][14] , 
	\sa_count[4][13] , \sa_count[4][12] , \sa_count[4][11] , 
	\sa_count[4][10] , \sa_count[4][9] , \sa_count[4][8] , 
	\sa_count[4][7] , \sa_count[4][6] , \sa_count[4][5] , 
	\sa_count[4][4] , \sa_count[4][3] , \sa_count[4][2] , 
	\sa_count[4][1] , \sa_count[4][0] , \sa_count[3][63] , 
	\sa_count[3][62] , \sa_count[3][61] , \sa_count[3][60] , 
	\sa_count[3][59] , \sa_count[3][58] , \sa_count[3][57] , 
	\sa_count[3][56] , \sa_count[3][55] , \sa_count[3][54] , 
	\sa_count[3][53] , \sa_count[3][52] , \sa_count[3][51] , 
	\sa_count[3][50] , \sa_count[3][49] , \sa_count[3][48] , 
	\sa_count[3][47] , \sa_count[3][46] , \sa_count[3][45] , 
	\sa_count[3][44] , \sa_count[3][43] , \sa_count[3][42] , 
	\sa_count[3][41] , \sa_count[3][40] , \sa_count[3][39] , 
	\sa_count[3][38] , \sa_count[3][37] , \sa_count[3][36] , 
	\sa_count[3][35] , \sa_count[3][34] , \sa_count[3][33] , 
	\sa_count[3][32] , \sa_count[3][31] , \sa_count[3][30] , 
	\sa_count[3][29] , \sa_count[3][28] , \sa_count[3][27] , 
	\sa_count[3][26] , \sa_count[3][25] , \sa_count[3][24] , 
	\sa_count[3][23] , \sa_count[3][22] , \sa_count[3][21] , 
	\sa_count[3][20] , \sa_count[3][19] , \sa_count[3][18] , 
	\sa_count[3][17] , \sa_count[3][16] , \sa_count[3][15] , 
	\sa_count[3][14] , \sa_count[3][13] , \sa_count[3][12] , 
	\sa_count[3][11] , \sa_count[3][10] , \sa_count[3][9] , 
	\sa_count[3][8] , \sa_count[3][7] , \sa_count[3][6] , 
	\sa_count[3][5] , \sa_count[3][4] , \sa_count[3][3] , 
	\sa_count[3][2] , \sa_count[3][1] , \sa_count[3][0] , 
	\sa_count[2][63] , \sa_count[2][62] , \sa_count[2][61] , 
	\sa_count[2][60] , \sa_count[2][59] , \sa_count[2][58] , 
	\sa_count[2][57] , \sa_count[2][56] , \sa_count[2][55] , 
	\sa_count[2][54] , \sa_count[2][53] , \sa_count[2][52] , 
	\sa_count[2][51] , \sa_count[2][50] , \sa_count[2][49] , 
	\sa_count[2][48] , \sa_count[2][47] , \sa_count[2][46] , 
	\sa_count[2][45] , \sa_count[2][44] , \sa_count[2][43] , 
	\sa_count[2][42] , \sa_count[2][41] , \sa_count[2][40] , 
	\sa_count[2][39] , \sa_count[2][38] , \sa_count[2][37] , 
	\sa_count[2][36] , \sa_count[2][35] , \sa_count[2][34] , 
	\sa_count[2][33] , \sa_count[2][32] , \sa_count[2][31] , 
	\sa_count[2][30] , \sa_count[2][29] , \sa_count[2][28] , 
	\sa_count[2][27] , \sa_count[2][26] , \sa_count[2][25] , 
	\sa_count[2][24] , \sa_count[2][23] , \sa_count[2][22] , 
	\sa_count[2][21] , \sa_count[2][20] , \sa_count[2][19] , 
	\sa_count[2][18] , \sa_count[2][17] , \sa_count[2][16] , 
	\sa_count[2][15] , \sa_count[2][14] , \sa_count[2][13] , 
	\sa_count[2][12] , \sa_count[2][11] , \sa_count[2][10] , 
	\sa_count[2][9] , \sa_count[2][8] , \sa_count[2][7] , 
	\sa_count[2][6] , \sa_count[2][5] , \sa_count[2][4] , 
	\sa_count[2][3] , \sa_count[2][2] , \sa_count[2][1] , 
	\sa_count[2][0] , \sa_count[1][63] , \sa_count[1][62] , 
	\sa_count[1][61] , \sa_count[1][60] , \sa_count[1][59] , 
	\sa_count[1][58] , \sa_count[1][57] , \sa_count[1][56] , 
	\sa_count[1][55] , \sa_count[1][54] , \sa_count[1][53] , 
	\sa_count[1][52] , \sa_count[1][51] , \sa_count[1][50] , 
	\sa_count[1][49] , \sa_count[1][48] , \sa_count[1][47] , 
	\sa_count[1][46] , \sa_count[1][45] , \sa_count[1][44] , 
	\sa_count[1][43] , \sa_count[1][42] , \sa_count[1][41] , 
	\sa_count[1][40] , \sa_count[1][39] , \sa_count[1][38] , 
	\sa_count[1][37] , \sa_count[1][36] , \sa_count[1][35] , 
	\sa_count[1][34] , \sa_count[1][33] , \sa_count[1][32] , 
	\sa_count[1][31] , \sa_count[1][30] , \sa_count[1][29] , 
	\sa_count[1][28] , \sa_count[1][27] , \sa_count[1][26] , 
	\sa_count[1][25] , \sa_count[1][24] , \sa_count[1][23] , 
	\sa_count[1][22] , \sa_count[1][21] , \sa_count[1][20] , 
	\sa_count[1][19] , \sa_count[1][18] , \sa_count[1][17] , 
	\sa_count[1][16] , \sa_count[1][15] , \sa_count[1][14] , 
	\sa_count[1][13] , \sa_count[1][12] , \sa_count[1][11] , 
	\sa_count[1][10] , \sa_count[1][9] , \sa_count[1][8] , 
	\sa_count[1][7] , \sa_count[1][6] , \sa_count[1][5] , 
	\sa_count[1][4] , \sa_count[1][3] , \sa_count[1][2] , 
	\sa_count[1][1] , \sa_count[1][0] , \sa_count[0][63] , 
	\sa_count[0][62] , \sa_count[0][61] , \sa_count[0][60] , 
	\sa_count[0][59] , \sa_count[0][58] , \sa_count[0][57] , 
	\sa_count[0][56] , \sa_count[0][55] , \sa_count[0][54] , 
	\sa_count[0][53] , \sa_count[0][52] , \sa_count[0][51] , 
	\sa_count[0][50] , \sa_count[0][49] , \sa_count[0][48] , 
	\sa_count[0][47] , \sa_count[0][46] , \sa_count[0][45] , 
	\sa_count[0][44] , \sa_count[0][43] , \sa_count[0][42] , 
	\sa_count[0][41] , \sa_count[0][40] , \sa_count[0][39] , 
	\sa_count[0][38] , \sa_count[0][37] , \sa_count[0][36] , 
	\sa_count[0][35] , \sa_count[0][34] , \sa_count[0][33] , 
	\sa_count[0][32] , \sa_count[0][31] , \sa_count[0][30] , 
	\sa_count[0][29] , \sa_count[0][28] , \sa_count[0][27] , 
	\sa_count[0][26] , \sa_count[0][25] , \sa_count[0][24] , 
	\sa_count[0][23] , \sa_count[0][22] , \sa_count[0][21] , 
	\sa_count[0][20] , \sa_count[0][19] , \sa_count[0][18] , 
	\sa_count[0][17] , \sa_count[0][16] , \sa_count[0][15] , 
	\sa_count[0][14] , \sa_count[0][13] , \sa_count[0][12] , 
	\sa_count[0][11] , \sa_count[0][10] , \sa_count[0][9] , 
	\sa_count[0][8] , \sa_count[0][7] , \sa_count[0][6] , 
	\sa_count[0][5] , \sa_count[0][4] , \sa_count[0][3] , 
	\sa_count[0][2] , \sa_count[0][1] , \sa_count[0][0] }), .kme_idle( 
	kme_idle), .clk( clk), .rst_n( rst_sync_n), .scan_en( scan_en), 
	.scan_mode( scan_mode), .scan_rst_n( scan_rst_n), 
	.disable_debug_cmd( disable_debug_cmd), .disable_unencrypted_keys( 
	disable_unencrypted_keys), .suppress_key_tlvs( suppress_key_tlvs), 
	.always_validate_kim_ref( always_validate_kim_ref), .kme_ib_in( 
	_zy_simnet_kme_ib_in_10_w$[0:82]), .kme_cceip0_ob_in( 
	_zy_simnet_kme_cceip0_ob_in_mod_11_w$), .kme_cceip1_ob_in( 
	_zy_simnet_kme_cceip1_ob_in_mod_12_w$), .kme_cceip2_ob_in( 
	_zy_simnet_kme_cceip2_ob_in_mod_13_w$), .kme_cceip3_ob_in( 
	_zy_simnet_kme_cceip3_ob_in_mod_14_w$), .kme_cddip0_ob_in( 
	_zy_simnet_kme_cddip0_ob_in_mod_15_w$), .kme_cddip1_ob_in( 
	_zy_simnet_kme_cddip1_ob_in_mod_16_w$), .kme_cddip2_ob_in( 
	_zy_simnet_kme_cddip2_ob_in_mod_17_w$), .kme_cddip3_ob_in( 
	_zy_simnet_kme_cddip3_ob_in_mod_18_w$), .ckv_dout( ckv_dout[63:0]), 
	.ckv_mbe( ckv_mbe), .kim_dout( _zy_simnet_kim_dout_19_w$[0:37]), 
	.kim_mbe( kim_mbe), .bimc_rst_n( bimc_rst_n), 
	.cceip_encrypt_bimc_isync( cceip_encrypt_bimc_isync), 
	.cceip_encrypt_bimc_idat( cceip_encrypt_bimc_idat), 
	.cceip_validate_bimc_isync( cceip_validate_bimc_isync), 
	.cceip_validate_bimc_idat( cceip_validate_bimc_idat), 
	.cddip_decrypt_bimc_isync( cddip_decrypt_bimc_isync), 
	.cddip_decrypt_bimc_idat( cddip_decrypt_bimc_idat), 
	.axi_bimc_isync( axi_bimc_isync), .axi_bimc_idat( axi_bimc_idat), 
	.labels( { \_zy_simnet_tvar_20[7][271] , 
	\_zy_simnet_tvar_20[7][270] , \_zy_simnet_tvar_20[7][269] , 
	\_zy_simnet_tvar_20[7][268] , \_zy_simnet_tvar_20[7][267] , 
	\_zy_simnet_tvar_20[7][266] , \_zy_simnet_tvar_20[7][265] , 
	\_zy_simnet_tvar_20[7][264] , \_zy_simnet_tvar_20[7][263] , 
	\_zy_simnet_tvar_20[7][262] , \_zy_simnet_tvar_20[7][261] , 
	\_zy_simnet_tvar_20[7][260] , \_zy_simnet_tvar_20[7][259] , 
	\_zy_simnet_tvar_20[7][258] , \_zy_simnet_tvar_20[7][257] , 
	\_zy_simnet_tvar_20[7][256] , \_zy_simnet_tvar_20[7][255] , 
	\_zy_simnet_tvar_20[7][254] , \_zy_simnet_tvar_20[7][253] , 
	\_zy_simnet_tvar_20[7][252] , \_zy_simnet_tvar_20[7][251] , 
	\_zy_simnet_tvar_20[7][250] , \_zy_simnet_tvar_20[7][249] , 
	\_zy_simnet_tvar_20[7][248] , \_zy_simnet_tvar_20[7][247] , 
	\_zy_simnet_tvar_20[7][246] , \_zy_simnet_tvar_20[7][245] , 
	\_zy_simnet_tvar_20[7][244] , \_zy_simnet_tvar_20[7][243] , 
	\_zy_simnet_tvar_20[7][242] , \_zy_simnet_tvar_20[7][241] , 
	\_zy_simnet_tvar_20[7][240] , \_zy_simnet_tvar_20[7][239] , 
	\_zy_simnet_tvar_20[7][238] , \_zy_simnet_tvar_20[7][237] , 
	\_zy_simnet_tvar_20[7][236] , \_zy_simnet_tvar_20[7][235] , 
	\_zy_simnet_tvar_20[7][234] , \_zy_simnet_tvar_20[7][233] , 
	\_zy_simnet_tvar_20[7][232] , \_zy_simnet_tvar_20[7][231] , 
	\_zy_simnet_tvar_20[7][230] , \_zy_simnet_tvar_20[7][229] , 
	\_zy_simnet_tvar_20[7][228] , \_zy_simnet_tvar_20[7][227] , 
	\_zy_simnet_tvar_20[7][226] , \_zy_simnet_tvar_20[7][225] , 
	\_zy_simnet_tvar_20[7][224] , \_zy_simnet_tvar_20[7][223] , 
	\_zy_simnet_tvar_20[7][222] , \_zy_simnet_tvar_20[7][221] , 
	\_zy_simnet_tvar_20[7][220] , \_zy_simnet_tvar_20[7][219] , 
	\_zy_simnet_tvar_20[7][218] , \_zy_simnet_tvar_20[7][217] , 
	\_zy_simnet_tvar_20[7][216] , \_zy_simnet_tvar_20[7][215] , 
	\_zy_simnet_tvar_20[7][214] , \_zy_simnet_tvar_20[7][213] , 
	\_zy_simnet_tvar_20[7][212] , \_zy_simnet_tvar_20[7][211] , 
	\_zy_simnet_tvar_20[7][210] , \_zy_simnet_tvar_20[7][209] , 
	\_zy_simnet_tvar_20[7][208] , \_zy_simnet_tvar_20[7][207] , 
	\_zy_simnet_tvar_20[7][206] , \_zy_simnet_tvar_20[7][205] , 
	\_zy_simnet_tvar_20[7][204] , \_zy_simnet_tvar_20[7][203] , 
	\_zy_simnet_tvar_20[7][202] , \_zy_simnet_tvar_20[7][201] , 
	\_zy_simnet_tvar_20[7][200] , \_zy_simnet_tvar_20[7][199] , 
	\_zy_simnet_tvar_20[7][198] , \_zy_simnet_tvar_20[7][197] , 
	\_zy_simnet_tvar_20[7][196] , \_zy_simnet_tvar_20[7][195] , 
	\_zy_simnet_tvar_20[7][194] , \_zy_simnet_tvar_20[7][193] , 
	\_zy_simnet_tvar_20[7][192] , \_zy_simnet_tvar_20[7][191] , 
	\_zy_simnet_tvar_20[7][190] , \_zy_simnet_tvar_20[7][189] , 
	\_zy_simnet_tvar_20[7][188] , \_zy_simnet_tvar_20[7][187] , 
	\_zy_simnet_tvar_20[7][186] , \_zy_simnet_tvar_20[7][185] , 
	\_zy_simnet_tvar_20[7][184] , \_zy_simnet_tvar_20[7][183] , 
	\_zy_simnet_tvar_20[7][182] , \_zy_simnet_tvar_20[7][181] , 
	\_zy_simnet_tvar_20[7][180] , \_zy_simnet_tvar_20[7][179] , 
	\_zy_simnet_tvar_20[7][178] , \_zy_simnet_tvar_20[7][177] , 
	\_zy_simnet_tvar_20[7][176] , \_zy_simnet_tvar_20[7][175] , 
	\_zy_simnet_tvar_20[7][174] , \_zy_simnet_tvar_20[7][173] , 
	\_zy_simnet_tvar_20[7][172] , \_zy_simnet_tvar_20[7][171] , 
	\_zy_simnet_tvar_20[7][170] , \_zy_simnet_tvar_20[7][169] , 
	\_zy_simnet_tvar_20[7][168] , \_zy_simnet_tvar_20[7][167] , 
	\_zy_simnet_tvar_20[7][166] , \_zy_simnet_tvar_20[7][165] , 
	\_zy_simnet_tvar_20[7][164] , \_zy_simnet_tvar_20[7][163] , 
	\_zy_simnet_tvar_20[7][162] , \_zy_simnet_tvar_20[7][161] , 
	\_zy_simnet_tvar_20[7][160] , \_zy_simnet_tvar_20[7][159] , 
	\_zy_simnet_tvar_20[7][158] , \_zy_simnet_tvar_20[7][157] , 
	\_zy_simnet_tvar_20[7][156] , \_zy_simnet_tvar_20[7][155] , 
	\_zy_simnet_tvar_20[7][154] , \_zy_simnet_tvar_20[7][153] , 
	\_zy_simnet_tvar_20[7][152] , \_zy_simnet_tvar_20[7][151] , 
	\_zy_simnet_tvar_20[7][150] , \_zy_simnet_tvar_20[7][149] , 
	\_zy_simnet_tvar_20[7][148] , \_zy_simnet_tvar_20[7][147] , 
	\_zy_simnet_tvar_20[7][146] , \_zy_simnet_tvar_20[7][145] , 
	\_zy_simnet_tvar_20[7][144] , \_zy_simnet_tvar_20[7][143] , 
	\_zy_simnet_tvar_20[7][142] , \_zy_simnet_tvar_20[7][141] , 
	\_zy_simnet_tvar_20[7][140] , \_zy_simnet_tvar_20[7][139] , 
	\_zy_simnet_tvar_20[7][138] , \_zy_simnet_tvar_20[7][137] , 
	\_zy_simnet_tvar_20[7][136] , \_zy_simnet_tvar_20[7][135] , 
	\_zy_simnet_tvar_20[7][134] , \_zy_simnet_tvar_20[7][133] , 
	\_zy_simnet_tvar_20[7][132] , \_zy_simnet_tvar_20[7][131] , 
	\_zy_simnet_tvar_20[7][130] , \_zy_simnet_tvar_20[7][129] , 
	\_zy_simnet_tvar_20[7][128] , \_zy_simnet_tvar_20[7][127] , 
	\_zy_simnet_tvar_20[7][126] , \_zy_simnet_tvar_20[7][125] , 
	\_zy_simnet_tvar_20[7][124] , \_zy_simnet_tvar_20[7][123] , 
	\_zy_simnet_tvar_20[7][122] , \_zy_simnet_tvar_20[7][121] , 
	\_zy_simnet_tvar_20[7][120] , \_zy_simnet_tvar_20[7][119] , 
	\_zy_simnet_tvar_20[7][118] , \_zy_simnet_tvar_20[7][117] , 
	\_zy_simnet_tvar_20[7][116] , \_zy_simnet_tvar_20[7][115] , 
	\_zy_simnet_tvar_20[7][114] , \_zy_simnet_tvar_20[7][113] , 
	\_zy_simnet_tvar_20[7][112] , \_zy_simnet_tvar_20[7][111] , 
	\_zy_simnet_tvar_20[7][110] , \_zy_simnet_tvar_20[7][109] , 
	\_zy_simnet_tvar_20[7][108] , \_zy_simnet_tvar_20[7][107] , 
	\_zy_simnet_tvar_20[7][106] , \_zy_simnet_tvar_20[7][105] , 
	\_zy_simnet_tvar_20[7][104] , \_zy_simnet_tvar_20[7][103] , 
	\_zy_simnet_tvar_20[7][102] , \_zy_simnet_tvar_20[7][101] , 
	\_zy_simnet_tvar_20[7][100] , \_zy_simnet_tvar_20[7][99] , 
	\_zy_simnet_tvar_20[7][98] , \_zy_simnet_tvar_20[7][97] , 
	\_zy_simnet_tvar_20[7][96] , \_zy_simnet_tvar_20[7][95] , 
	\_zy_simnet_tvar_20[7][94] , \_zy_simnet_tvar_20[7][93] , 
	\_zy_simnet_tvar_20[7][92] , \_zy_simnet_tvar_20[7][91] , 
	\_zy_simnet_tvar_20[7][90] , \_zy_simnet_tvar_20[7][89] , 
	\_zy_simnet_tvar_20[7][88] , \_zy_simnet_tvar_20[7][87] , 
	\_zy_simnet_tvar_20[7][86] , \_zy_simnet_tvar_20[7][85] , 
	\_zy_simnet_tvar_20[7][84] , \_zy_simnet_tvar_20[7][83] , 
	\_zy_simnet_tvar_20[7][82] , \_zy_simnet_tvar_20[7][81] , 
	\_zy_simnet_tvar_20[7][80] , \_zy_simnet_tvar_20[7][79] , 
	\_zy_simnet_tvar_20[7][78] , \_zy_simnet_tvar_20[7][77] , 
	\_zy_simnet_tvar_20[7][76] , \_zy_simnet_tvar_20[7][75] , 
	\_zy_simnet_tvar_20[7][74] , \_zy_simnet_tvar_20[7][73] , 
	\_zy_simnet_tvar_20[7][72] , \_zy_simnet_tvar_20[7][71] , 
	\_zy_simnet_tvar_20[7][70] , \_zy_simnet_tvar_20[7][69] , 
	\_zy_simnet_tvar_20[7][68] , \_zy_simnet_tvar_20[7][67] , 
	\_zy_simnet_tvar_20[7][66] , \_zy_simnet_tvar_20[7][65] , 
	\_zy_simnet_tvar_20[7][64] , \_zy_simnet_tvar_20[7][63] , 
	\_zy_simnet_tvar_20[7][62] , \_zy_simnet_tvar_20[7][61] , 
	\_zy_simnet_tvar_20[7][60] , \_zy_simnet_tvar_20[7][59] , 
	\_zy_simnet_tvar_20[7][58] , \_zy_simnet_tvar_20[7][57] , 
	\_zy_simnet_tvar_20[7][56] , \_zy_simnet_tvar_20[7][55] , 
	\_zy_simnet_tvar_20[7][54] , \_zy_simnet_tvar_20[7][53] , 
	\_zy_simnet_tvar_20[7][52] , \_zy_simnet_tvar_20[7][51] , 
	\_zy_simnet_tvar_20[7][50] , \_zy_simnet_tvar_20[7][49] , 
	\_zy_simnet_tvar_20[7][48] , \_zy_simnet_tvar_20[7][47] , 
	\_zy_simnet_tvar_20[7][46] , \_zy_simnet_tvar_20[7][45] , 
	\_zy_simnet_tvar_20[7][44] , \_zy_simnet_tvar_20[7][43] , 
	\_zy_simnet_tvar_20[7][42] , \_zy_simnet_tvar_20[7][41] , 
	\_zy_simnet_tvar_20[7][40] , \_zy_simnet_tvar_20[7][39] , 
	\_zy_simnet_tvar_20[7][38] , \_zy_simnet_tvar_20[7][37] , 
	\_zy_simnet_tvar_20[7][36] , \_zy_simnet_tvar_20[7][35] , 
	\_zy_simnet_tvar_20[7][34] , \_zy_simnet_tvar_20[7][33] , 
	\_zy_simnet_tvar_20[7][32] , \_zy_simnet_tvar_20[7][31] , 
	\_zy_simnet_tvar_20[7][30] , \_zy_simnet_tvar_20[7][29] , 
	\_zy_simnet_tvar_20[7][28] , \_zy_simnet_tvar_20[7][27] , 
	\_zy_simnet_tvar_20[7][26] , \_zy_simnet_tvar_20[7][25] , 
	\_zy_simnet_tvar_20[7][24] , \_zy_simnet_tvar_20[7][23] , 
	\_zy_simnet_tvar_20[7][22] , \_zy_simnet_tvar_20[7][21] , 
	\_zy_simnet_tvar_20[7][20] , \_zy_simnet_tvar_20[7][19] , 
	\_zy_simnet_tvar_20[7][18] , \_zy_simnet_tvar_20[7][17] , 
	\_zy_simnet_tvar_20[7][16] , \_zy_simnet_tvar_20[7][15] , 
	\_zy_simnet_tvar_20[7][14] , \_zy_simnet_tvar_20[7][13] , 
	\_zy_simnet_tvar_20[7][12] , \_zy_simnet_tvar_20[7][11] , 
	\_zy_simnet_tvar_20[7][10] , \_zy_simnet_tvar_20[7][9] , 
	\_zy_simnet_tvar_20[7][8] , \_zy_simnet_tvar_20[7][7] , 
	\_zy_simnet_tvar_20[7][6] , \_zy_simnet_tvar_20[7][5] , 
	\_zy_simnet_tvar_20[7][4] , \_zy_simnet_tvar_20[7][3] , 
	\_zy_simnet_tvar_20[7][2] , \_zy_simnet_tvar_20[7][1] , 
	\_zy_simnet_tvar_20[7][0] , \_zy_simnet_tvar_20[6][271] , 
	\_zy_simnet_tvar_20[6][270] , \_zy_simnet_tvar_20[6][269] , 
	\_zy_simnet_tvar_20[6][268] , \_zy_simnet_tvar_20[6][267] , 
	\_zy_simnet_tvar_20[6][266] , \_zy_simnet_tvar_20[6][265] , 
	\_zy_simnet_tvar_20[6][264] , \_zy_simnet_tvar_20[6][263] , 
	\_zy_simnet_tvar_20[6][262] , \_zy_simnet_tvar_20[6][261] , 
	\_zy_simnet_tvar_20[6][260] , \_zy_simnet_tvar_20[6][259] , 
	\_zy_simnet_tvar_20[6][258] , \_zy_simnet_tvar_20[6][257] , 
	\_zy_simnet_tvar_20[6][256] , \_zy_simnet_tvar_20[6][255] , 
	\_zy_simnet_tvar_20[6][254] , \_zy_simnet_tvar_20[6][253] , 
	\_zy_simnet_tvar_20[6][252] , \_zy_simnet_tvar_20[6][251] , 
	\_zy_simnet_tvar_20[6][250] , \_zy_simnet_tvar_20[6][249] , 
	\_zy_simnet_tvar_20[6][248] , \_zy_simnet_tvar_20[6][247] , 
	\_zy_simnet_tvar_20[6][246] , \_zy_simnet_tvar_20[6][245] , 
	\_zy_simnet_tvar_20[6][244] , \_zy_simnet_tvar_20[6][243] , 
	\_zy_simnet_tvar_20[6][242] , \_zy_simnet_tvar_20[6][241] , 
	\_zy_simnet_tvar_20[6][240] , \_zy_simnet_tvar_20[6][239] , 
	\_zy_simnet_tvar_20[6][238] , \_zy_simnet_tvar_20[6][237] , 
	\_zy_simnet_tvar_20[6][236] , \_zy_simnet_tvar_20[6][235] , 
	\_zy_simnet_tvar_20[6][234] , \_zy_simnet_tvar_20[6][233] , 
	\_zy_simnet_tvar_20[6][232] , \_zy_simnet_tvar_20[6][231] , 
	\_zy_simnet_tvar_20[6][230] , \_zy_simnet_tvar_20[6][229] , 
	\_zy_simnet_tvar_20[6][228] , \_zy_simnet_tvar_20[6][227] , 
	\_zy_simnet_tvar_20[6][226] , \_zy_simnet_tvar_20[6][225] , 
	\_zy_simnet_tvar_20[6][224] , \_zy_simnet_tvar_20[6][223] , 
	\_zy_simnet_tvar_20[6][222] , \_zy_simnet_tvar_20[6][221] , 
	\_zy_simnet_tvar_20[6][220] , \_zy_simnet_tvar_20[6][219] , 
	\_zy_simnet_tvar_20[6][218] , \_zy_simnet_tvar_20[6][217] , 
	\_zy_simnet_tvar_20[6][216] , \_zy_simnet_tvar_20[6][215] , 
	\_zy_simnet_tvar_20[6][214] , \_zy_simnet_tvar_20[6][213] , 
	\_zy_simnet_tvar_20[6][212] , \_zy_simnet_tvar_20[6][211] , 
	\_zy_simnet_tvar_20[6][210] , \_zy_simnet_tvar_20[6][209] , 
	\_zy_simnet_tvar_20[6][208] , \_zy_simnet_tvar_20[6][207] , 
	\_zy_simnet_tvar_20[6][206] , \_zy_simnet_tvar_20[6][205] , 
	\_zy_simnet_tvar_20[6][204] , \_zy_simnet_tvar_20[6][203] , 
	\_zy_simnet_tvar_20[6][202] , \_zy_simnet_tvar_20[6][201] , 
	\_zy_simnet_tvar_20[6][200] , \_zy_simnet_tvar_20[6][199] , 
	\_zy_simnet_tvar_20[6][198] , \_zy_simnet_tvar_20[6][197] , 
	\_zy_simnet_tvar_20[6][196] , \_zy_simnet_tvar_20[6][195] , 
	\_zy_simnet_tvar_20[6][194] , \_zy_simnet_tvar_20[6][193] , 
	\_zy_simnet_tvar_20[6][192] , \_zy_simnet_tvar_20[6][191] , 
	\_zy_simnet_tvar_20[6][190] , \_zy_simnet_tvar_20[6][189] , 
	\_zy_simnet_tvar_20[6][188] , \_zy_simnet_tvar_20[6][187] , 
	\_zy_simnet_tvar_20[6][186] , \_zy_simnet_tvar_20[6][185] , 
	\_zy_simnet_tvar_20[6][184] , \_zy_simnet_tvar_20[6][183] , 
	\_zy_simnet_tvar_20[6][182] , \_zy_simnet_tvar_20[6][181] , 
	\_zy_simnet_tvar_20[6][180] , \_zy_simnet_tvar_20[6][179] , 
	\_zy_simnet_tvar_20[6][178] , \_zy_simnet_tvar_20[6][177] , 
	\_zy_simnet_tvar_20[6][176] , \_zy_simnet_tvar_20[6][175] , 
	\_zy_simnet_tvar_20[6][174] , \_zy_simnet_tvar_20[6][173] , 
	\_zy_simnet_tvar_20[6][172] , \_zy_simnet_tvar_20[6][171] , 
	\_zy_simnet_tvar_20[6][170] , \_zy_simnet_tvar_20[6][169] , 
	\_zy_simnet_tvar_20[6][168] , \_zy_simnet_tvar_20[6][167] , 
	\_zy_simnet_tvar_20[6][166] , \_zy_simnet_tvar_20[6][165] , 
	\_zy_simnet_tvar_20[6][164] , \_zy_simnet_tvar_20[6][163] , 
	\_zy_simnet_tvar_20[6][162] , \_zy_simnet_tvar_20[6][161] , 
	\_zy_simnet_tvar_20[6][160] , \_zy_simnet_tvar_20[6][159] , 
	\_zy_simnet_tvar_20[6][158] , \_zy_simnet_tvar_20[6][157] , 
	\_zy_simnet_tvar_20[6][156] , \_zy_simnet_tvar_20[6][155] , 
	\_zy_simnet_tvar_20[6][154] , \_zy_simnet_tvar_20[6][153] , 
	\_zy_simnet_tvar_20[6][152] , \_zy_simnet_tvar_20[6][151] , 
	\_zy_simnet_tvar_20[6][150] , \_zy_simnet_tvar_20[6][149] , 
	\_zy_simnet_tvar_20[6][148] , \_zy_simnet_tvar_20[6][147] , 
	\_zy_simnet_tvar_20[6][146] , \_zy_simnet_tvar_20[6][145] , 
	\_zy_simnet_tvar_20[6][144] , \_zy_simnet_tvar_20[6][143] , 
	\_zy_simnet_tvar_20[6][142] , \_zy_simnet_tvar_20[6][141] , 
	\_zy_simnet_tvar_20[6][140] , \_zy_simnet_tvar_20[6][139] , 
	\_zy_simnet_tvar_20[6][138] , \_zy_simnet_tvar_20[6][137] , 
	\_zy_simnet_tvar_20[6][136] , \_zy_simnet_tvar_20[6][135] , 
	\_zy_simnet_tvar_20[6][134] , \_zy_simnet_tvar_20[6][133] , 
	\_zy_simnet_tvar_20[6][132] , \_zy_simnet_tvar_20[6][131] , 
	\_zy_simnet_tvar_20[6][130] , \_zy_simnet_tvar_20[6][129] , 
	\_zy_simnet_tvar_20[6][128] , \_zy_simnet_tvar_20[6][127] , 
	\_zy_simnet_tvar_20[6][126] , \_zy_simnet_tvar_20[6][125] , 
	\_zy_simnet_tvar_20[6][124] , \_zy_simnet_tvar_20[6][123] , 
	\_zy_simnet_tvar_20[6][122] , \_zy_simnet_tvar_20[6][121] , 
	\_zy_simnet_tvar_20[6][120] , \_zy_simnet_tvar_20[6][119] , 
	\_zy_simnet_tvar_20[6][118] , \_zy_simnet_tvar_20[6][117] , 
	\_zy_simnet_tvar_20[6][116] , \_zy_simnet_tvar_20[6][115] , 
	\_zy_simnet_tvar_20[6][114] , \_zy_simnet_tvar_20[6][113] , 
	\_zy_simnet_tvar_20[6][112] , \_zy_simnet_tvar_20[6][111] , 
	\_zy_simnet_tvar_20[6][110] , \_zy_simnet_tvar_20[6][109] , 
	\_zy_simnet_tvar_20[6][108] , \_zy_simnet_tvar_20[6][107] , 
	\_zy_simnet_tvar_20[6][106] , \_zy_simnet_tvar_20[6][105] , 
	\_zy_simnet_tvar_20[6][104] , \_zy_simnet_tvar_20[6][103] , 
	\_zy_simnet_tvar_20[6][102] , \_zy_simnet_tvar_20[6][101] , 
	\_zy_simnet_tvar_20[6][100] , \_zy_simnet_tvar_20[6][99] , 
	\_zy_simnet_tvar_20[6][98] , \_zy_simnet_tvar_20[6][97] , 
	\_zy_simnet_tvar_20[6][96] , \_zy_simnet_tvar_20[6][95] , 
	\_zy_simnet_tvar_20[6][94] , \_zy_simnet_tvar_20[6][93] , 
	\_zy_simnet_tvar_20[6][92] , \_zy_simnet_tvar_20[6][91] , 
	\_zy_simnet_tvar_20[6][90] , \_zy_simnet_tvar_20[6][89] , 
	\_zy_simnet_tvar_20[6][88] , \_zy_simnet_tvar_20[6][87] , 
	\_zy_simnet_tvar_20[6][86] , \_zy_simnet_tvar_20[6][85] , 
	\_zy_simnet_tvar_20[6][84] , \_zy_simnet_tvar_20[6][83] , 
	\_zy_simnet_tvar_20[6][82] , \_zy_simnet_tvar_20[6][81] , 
	\_zy_simnet_tvar_20[6][80] , \_zy_simnet_tvar_20[6][79] , 
	\_zy_simnet_tvar_20[6][78] , \_zy_simnet_tvar_20[6][77] , 
	\_zy_simnet_tvar_20[6][76] , \_zy_simnet_tvar_20[6][75] , 
	\_zy_simnet_tvar_20[6][74] , \_zy_simnet_tvar_20[6][73] , 
	\_zy_simnet_tvar_20[6][72] , \_zy_simnet_tvar_20[6][71] , 
	\_zy_simnet_tvar_20[6][70] , \_zy_simnet_tvar_20[6][69] , 
	\_zy_simnet_tvar_20[6][68] , \_zy_simnet_tvar_20[6][67] , 
	\_zy_simnet_tvar_20[6][66] , \_zy_simnet_tvar_20[6][65] , 
	\_zy_simnet_tvar_20[6][64] , \_zy_simnet_tvar_20[6][63] , 
	\_zy_simnet_tvar_20[6][62] , \_zy_simnet_tvar_20[6][61] , 
	\_zy_simnet_tvar_20[6][60] , \_zy_simnet_tvar_20[6][59] , 
	\_zy_simnet_tvar_20[6][58] , \_zy_simnet_tvar_20[6][57] , 
	\_zy_simnet_tvar_20[6][56] , \_zy_simnet_tvar_20[6][55] , 
	\_zy_simnet_tvar_20[6][54] , \_zy_simnet_tvar_20[6][53] , 
	\_zy_simnet_tvar_20[6][52] , \_zy_simnet_tvar_20[6][51] , 
	\_zy_simnet_tvar_20[6][50] , \_zy_simnet_tvar_20[6][49] , 
	\_zy_simnet_tvar_20[6][48] , \_zy_simnet_tvar_20[6][47] , 
	\_zy_simnet_tvar_20[6][46] , \_zy_simnet_tvar_20[6][45] , 
	\_zy_simnet_tvar_20[6][44] , \_zy_simnet_tvar_20[6][43] , 
	\_zy_simnet_tvar_20[6][42] , \_zy_simnet_tvar_20[6][41] , 
	\_zy_simnet_tvar_20[6][40] , \_zy_simnet_tvar_20[6][39] , 
	\_zy_simnet_tvar_20[6][38] , \_zy_simnet_tvar_20[6][37] , 
	\_zy_simnet_tvar_20[6][36] , \_zy_simnet_tvar_20[6][35] , 
	\_zy_simnet_tvar_20[6][34] , \_zy_simnet_tvar_20[6][33] , 
	\_zy_simnet_tvar_20[6][32] , \_zy_simnet_tvar_20[6][31] , 
	\_zy_simnet_tvar_20[6][30] , \_zy_simnet_tvar_20[6][29] , 
	\_zy_simnet_tvar_20[6][28] , \_zy_simnet_tvar_20[6][27] , 
	\_zy_simnet_tvar_20[6][26] , \_zy_simnet_tvar_20[6][25] , 
	\_zy_simnet_tvar_20[6][24] , \_zy_simnet_tvar_20[6][23] , 
	\_zy_simnet_tvar_20[6][22] , \_zy_simnet_tvar_20[6][21] , 
	\_zy_simnet_tvar_20[6][20] , \_zy_simnet_tvar_20[6][19] , 
	\_zy_simnet_tvar_20[6][18] , \_zy_simnet_tvar_20[6][17] , 
	\_zy_simnet_tvar_20[6][16] , \_zy_simnet_tvar_20[6][15] , 
	\_zy_simnet_tvar_20[6][14] , \_zy_simnet_tvar_20[6][13] , 
	\_zy_simnet_tvar_20[6][12] , \_zy_simnet_tvar_20[6][11] , 
	\_zy_simnet_tvar_20[6][10] , \_zy_simnet_tvar_20[6][9] , 
	\_zy_simnet_tvar_20[6][8] , \_zy_simnet_tvar_20[6][7] , 
	\_zy_simnet_tvar_20[6][6] , \_zy_simnet_tvar_20[6][5] , 
	\_zy_simnet_tvar_20[6][4] , \_zy_simnet_tvar_20[6][3] , 
	\_zy_simnet_tvar_20[6][2] , \_zy_simnet_tvar_20[6][1] , 
	\_zy_simnet_tvar_20[6][0] , \_zy_simnet_tvar_20[5][271] , 
	\_zy_simnet_tvar_20[5][270] , \_zy_simnet_tvar_20[5][269] , 
	\_zy_simnet_tvar_20[5][268] , \_zy_simnet_tvar_20[5][267] , 
	\_zy_simnet_tvar_20[5][266] , \_zy_simnet_tvar_20[5][265] , 
	\_zy_simnet_tvar_20[5][264] , \_zy_simnet_tvar_20[5][263] , 
	\_zy_simnet_tvar_20[5][262] , \_zy_simnet_tvar_20[5][261] , 
	\_zy_simnet_tvar_20[5][260] , \_zy_simnet_tvar_20[5][259] , 
	\_zy_simnet_tvar_20[5][258] , \_zy_simnet_tvar_20[5][257] , 
	\_zy_simnet_tvar_20[5][256] , \_zy_simnet_tvar_20[5][255] , 
	\_zy_simnet_tvar_20[5][254] , \_zy_simnet_tvar_20[5][253] , 
	\_zy_simnet_tvar_20[5][252] , \_zy_simnet_tvar_20[5][251] , 
	\_zy_simnet_tvar_20[5][250] , \_zy_simnet_tvar_20[5][249] , 
	\_zy_simnet_tvar_20[5][248] , \_zy_simnet_tvar_20[5][247] , 
	\_zy_simnet_tvar_20[5][246] , \_zy_simnet_tvar_20[5][245] , 
	\_zy_simnet_tvar_20[5][244] , \_zy_simnet_tvar_20[5][243] , 
	\_zy_simnet_tvar_20[5][242] , \_zy_simnet_tvar_20[5][241] , 
	\_zy_simnet_tvar_20[5][240] , \_zy_simnet_tvar_20[5][239] , 
	\_zy_simnet_tvar_20[5][238] , \_zy_simnet_tvar_20[5][237] , 
	\_zy_simnet_tvar_20[5][236] , \_zy_simnet_tvar_20[5][235] , 
	\_zy_simnet_tvar_20[5][234] , \_zy_simnet_tvar_20[5][233] , 
	\_zy_simnet_tvar_20[5][232] , \_zy_simnet_tvar_20[5][231] , 
	\_zy_simnet_tvar_20[5][230] , \_zy_simnet_tvar_20[5][229] , 
	\_zy_simnet_tvar_20[5][228] , \_zy_simnet_tvar_20[5][227] , 
	\_zy_simnet_tvar_20[5][226] , \_zy_simnet_tvar_20[5][225] , 
	\_zy_simnet_tvar_20[5][224] , \_zy_simnet_tvar_20[5][223] , 
	\_zy_simnet_tvar_20[5][222] , \_zy_simnet_tvar_20[5][221] , 
	\_zy_simnet_tvar_20[5][220] , \_zy_simnet_tvar_20[5][219] , 
	\_zy_simnet_tvar_20[5][218] , \_zy_simnet_tvar_20[5][217] , 
	\_zy_simnet_tvar_20[5][216] , \_zy_simnet_tvar_20[5][215] , 
	\_zy_simnet_tvar_20[5][214] , \_zy_simnet_tvar_20[5][213] , 
	\_zy_simnet_tvar_20[5][212] , \_zy_simnet_tvar_20[5][211] , 
	\_zy_simnet_tvar_20[5][210] , \_zy_simnet_tvar_20[5][209] , 
	\_zy_simnet_tvar_20[5][208] , \_zy_simnet_tvar_20[5][207] , 
	\_zy_simnet_tvar_20[5][206] , \_zy_simnet_tvar_20[5][205] , 
	\_zy_simnet_tvar_20[5][204] , \_zy_simnet_tvar_20[5][203] , 
	\_zy_simnet_tvar_20[5][202] , \_zy_simnet_tvar_20[5][201] , 
	\_zy_simnet_tvar_20[5][200] , \_zy_simnet_tvar_20[5][199] , 
	\_zy_simnet_tvar_20[5][198] , \_zy_simnet_tvar_20[5][197] , 
	\_zy_simnet_tvar_20[5][196] , \_zy_simnet_tvar_20[5][195] , 
	\_zy_simnet_tvar_20[5][194] , \_zy_simnet_tvar_20[5][193] , 
	\_zy_simnet_tvar_20[5][192] , \_zy_simnet_tvar_20[5][191] , 
	\_zy_simnet_tvar_20[5][190] , \_zy_simnet_tvar_20[5][189] , 
	\_zy_simnet_tvar_20[5][188] , \_zy_simnet_tvar_20[5][187] , 
	\_zy_simnet_tvar_20[5][186] , \_zy_simnet_tvar_20[5][185] , 
	\_zy_simnet_tvar_20[5][184] , \_zy_simnet_tvar_20[5][183] , 
	\_zy_simnet_tvar_20[5][182] , \_zy_simnet_tvar_20[5][181] , 
	\_zy_simnet_tvar_20[5][180] , \_zy_simnet_tvar_20[5][179] , 
	\_zy_simnet_tvar_20[5][178] , \_zy_simnet_tvar_20[5][177] , 
	\_zy_simnet_tvar_20[5][176] , \_zy_simnet_tvar_20[5][175] , 
	\_zy_simnet_tvar_20[5][174] , \_zy_simnet_tvar_20[5][173] , 
	\_zy_simnet_tvar_20[5][172] , \_zy_simnet_tvar_20[5][171] , 
	\_zy_simnet_tvar_20[5][170] , \_zy_simnet_tvar_20[5][169] , 
	\_zy_simnet_tvar_20[5][168] , \_zy_simnet_tvar_20[5][167] , 
	\_zy_simnet_tvar_20[5][166] , \_zy_simnet_tvar_20[5][165] , 
	\_zy_simnet_tvar_20[5][164] , \_zy_simnet_tvar_20[5][163] , 
	\_zy_simnet_tvar_20[5][162] , \_zy_simnet_tvar_20[5][161] , 
	\_zy_simnet_tvar_20[5][160] , \_zy_simnet_tvar_20[5][159] , 
	\_zy_simnet_tvar_20[5][158] , \_zy_simnet_tvar_20[5][157] , 
	\_zy_simnet_tvar_20[5][156] , \_zy_simnet_tvar_20[5][155] , 
	\_zy_simnet_tvar_20[5][154] , \_zy_simnet_tvar_20[5][153] , 
	\_zy_simnet_tvar_20[5][152] , \_zy_simnet_tvar_20[5][151] , 
	\_zy_simnet_tvar_20[5][150] , \_zy_simnet_tvar_20[5][149] , 
	\_zy_simnet_tvar_20[5][148] , \_zy_simnet_tvar_20[5][147] , 
	\_zy_simnet_tvar_20[5][146] , \_zy_simnet_tvar_20[5][145] , 
	\_zy_simnet_tvar_20[5][144] , \_zy_simnet_tvar_20[5][143] , 
	\_zy_simnet_tvar_20[5][142] , \_zy_simnet_tvar_20[5][141] , 
	\_zy_simnet_tvar_20[5][140] , \_zy_simnet_tvar_20[5][139] , 
	\_zy_simnet_tvar_20[5][138] , \_zy_simnet_tvar_20[5][137] , 
	\_zy_simnet_tvar_20[5][136] , \_zy_simnet_tvar_20[5][135] , 
	\_zy_simnet_tvar_20[5][134] , \_zy_simnet_tvar_20[5][133] , 
	\_zy_simnet_tvar_20[5][132] , \_zy_simnet_tvar_20[5][131] , 
	\_zy_simnet_tvar_20[5][130] , \_zy_simnet_tvar_20[5][129] , 
	\_zy_simnet_tvar_20[5][128] , \_zy_simnet_tvar_20[5][127] , 
	\_zy_simnet_tvar_20[5][126] , \_zy_simnet_tvar_20[5][125] , 
	\_zy_simnet_tvar_20[5][124] , \_zy_simnet_tvar_20[5][123] , 
	\_zy_simnet_tvar_20[5][122] , \_zy_simnet_tvar_20[5][121] , 
	\_zy_simnet_tvar_20[5][120] , \_zy_simnet_tvar_20[5][119] , 
	\_zy_simnet_tvar_20[5][118] , \_zy_simnet_tvar_20[5][117] , 
	\_zy_simnet_tvar_20[5][116] , \_zy_simnet_tvar_20[5][115] , 
	\_zy_simnet_tvar_20[5][114] , \_zy_simnet_tvar_20[5][113] , 
	\_zy_simnet_tvar_20[5][112] , \_zy_simnet_tvar_20[5][111] , 
	\_zy_simnet_tvar_20[5][110] , \_zy_simnet_tvar_20[5][109] , 
	\_zy_simnet_tvar_20[5][108] , \_zy_simnet_tvar_20[5][107] , 
	\_zy_simnet_tvar_20[5][106] , \_zy_simnet_tvar_20[5][105] , 
	\_zy_simnet_tvar_20[5][104] , \_zy_simnet_tvar_20[5][103] , 
	\_zy_simnet_tvar_20[5][102] , \_zy_simnet_tvar_20[5][101] , 
	\_zy_simnet_tvar_20[5][100] , \_zy_simnet_tvar_20[5][99] , 
	\_zy_simnet_tvar_20[5][98] , \_zy_simnet_tvar_20[5][97] , 
	\_zy_simnet_tvar_20[5][96] , \_zy_simnet_tvar_20[5][95] , 
	\_zy_simnet_tvar_20[5][94] , \_zy_simnet_tvar_20[5][93] , 
	\_zy_simnet_tvar_20[5][92] , \_zy_simnet_tvar_20[5][91] , 
	\_zy_simnet_tvar_20[5][90] , \_zy_simnet_tvar_20[5][89] , 
	\_zy_simnet_tvar_20[5][88] , \_zy_simnet_tvar_20[5][87] , 
	\_zy_simnet_tvar_20[5][86] , \_zy_simnet_tvar_20[5][85] , 
	\_zy_simnet_tvar_20[5][84] , \_zy_simnet_tvar_20[5][83] , 
	\_zy_simnet_tvar_20[5][82] , \_zy_simnet_tvar_20[5][81] , 
	\_zy_simnet_tvar_20[5][80] , \_zy_simnet_tvar_20[5][79] , 
	\_zy_simnet_tvar_20[5][78] , \_zy_simnet_tvar_20[5][77] , 
	\_zy_simnet_tvar_20[5][76] , \_zy_simnet_tvar_20[5][75] , 
	\_zy_simnet_tvar_20[5][74] , \_zy_simnet_tvar_20[5][73] , 
	\_zy_simnet_tvar_20[5][72] , \_zy_simnet_tvar_20[5][71] , 
	\_zy_simnet_tvar_20[5][70] , \_zy_simnet_tvar_20[5][69] , 
	\_zy_simnet_tvar_20[5][68] , \_zy_simnet_tvar_20[5][67] , 
	\_zy_simnet_tvar_20[5][66] , \_zy_simnet_tvar_20[5][65] , 
	\_zy_simnet_tvar_20[5][64] , \_zy_simnet_tvar_20[5][63] , 
	\_zy_simnet_tvar_20[5][62] , \_zy_simnet_tvar_20[5][61] , 
	\_zy_simnet_tvar_20[5][60] , \_zy_simnet_tvar_20[5][59] , 
	\_zy_simnet_tvar_20[5][58] , \_zy_simnet_tvar_20[5][57] , 
	\_zy_simnet_tvar_20[5][56] , \_zy_simnet_tvar_20[5][55] , 
	\_zy_simnet_tvar_20[5][54] , \_zy_simnet_tvar_20[5][53] , 
	\_zy_simnet_tvar_20[5][52] , \_zy_simnet_tvar_20[5][51] , 
	\_zy_simnet_tvar_20[5][50] , \_zy_simnet_tvar_20[5][49] , 
	\_zy_simnet_tvar_20[5][48] , \_zy_simnet_tvar_20[5][47] , 
	\_zy_simnet_tvar_20[5][46] , \_zy_simnet_tvar_20[5][45] , 
	\_zy_simnet_tvar_20[5][44] , \_zy_simnet_tvar_20[5][43] , 
	\_zy_simnet_tvar_20[5][42] , \_zy_simnet_tvar_20[5][41] , 
	\_zy_simnet_tvar_20[5][40] , \_zy_simnet_tvar_20[5][39] , 
	\_zy_simnet_tvar_20[5][38] , \_zy_simnet_tvar_20[5][37] , 
	\_zy_simnet_tvar_20[5][36] , \_zy_simnet_tvar_20[5][35] , 
	\_zy_simnet_tvar_20[5][34] , \_zy_simnet_tvar_20[5][33] , 
	\_zy_simnet_tvar_20[5][32] , \_zy_simnet_tvar_20[5][31] , 
	\_zy_simnet_tvar_20[5][30] , \_zy_simnet_tvar_20[5][29] , 
	\_zy_simnet_tvar_20[5][28] , \_zy_simnet_tvar_20[5][27] , 
	\_zy_simnet_tvar_20[5][26] , \_zy_simnet_tvar_20[5][25] , 
	\_zy_simnet_tvar_20[5][24] , \_zy_simnet_tvar_20[5][23] , 
	\_zy_simnet_tvar_20[5][22] , \_zy_simnet_tvar_20[5][21] , 
	\_zy_simnet_tvar_20[5][20] , \_zy_simnet_tvar_20[5][19] , 
	\_zy_simnet_tvar_20[5][18] , \_zy_simnet_tvar_20[5][17] , 
	\_zy_simnet_tvar_20[5][16] , \_zy_simnet_tvar_20[5][15] , 
	\_zy_simnet_tvar_20[5][14] , \_zy_simnet_tvar_20[5][13] , 
	\_zy_simnet_tvar_20[5][12] , \_zy_simnet_tvar_20[5][11] , 
	\_zy_simnet_tvar_20[5][10] , \_zy_simnet_tvar_20[5][9] , 
	\_zy_simnet_tvar_20[5][8] , \_zy_simnet_tvar_20[5][7] , 
	\_zy_simnet_tvar_20[5][6] , \_zy_simnet_tvar_20[5][5] , 
	\_zy_simnet_tvar_20[5][4] , \_zy_simnet_tvar_20[5][3] , 
	\_zy_simnet_tvar_20[5][2] , \_zy_simnet_tvar_20[5][1] , 
	\_zy_simnet_tvar_20[5][0] , \_zy_simnet_tvar_20[4][271] , 
	\_zy_simnet_tvar_20[4][270] , \_zy_simnet_tvar_20[4][269] , 
	\_zy_simnet_tvar_20[4][268] , \_zy_simnet_tvar_20[4][267] , 
	\_zy_simnet_tvar_20[4][266] , \_zy_simnet_tvar_20[4][265] , 
	\_zy_simnet_tvar_20[4][264] , \_zy_simnet_tvar_20[4][263] , 
	\_zy_simnet_tvar_20[4][262] , \_zy_simnet_tvar_20[4][261] , 
	\_zy_simnet_tvar_20[4][260] , \_zy_simnet_tvar_20[4][259] , 
	\_zy_simnet_tvar_20[4][258] , \_zy_simnet_tvar_20[4][257] , 
	\_zy_simnet_tvar_20[4][256] , \_zy_simnet_tvar_20[4][255] , 
	\_zy_simnet_tvar_20[4][254] , \_zy_simnet_tvar_20[4][253] , 
	\_zy_simnet_tvar_20[4][252] , \_zy_simnet_tvar_20[4][251] , 
	\_zy_simnet_tvar_20[4][250] , \_zy_simnet_tvar_20[4][249] , 
	\_zy_simnet_tvar_20[4][248] , \_zy_simnet_tvar_20[4][247] , 
	\_zy_simnet_tvar_20[4][246] , \_zy_simnet_tvar_20[4][245] , 
	\_zy_simnet_tvar_20[4][244] , \_zy_simnet_tvar_20[4][243] , 
	\_zy_simnet_tvar_20[4][242] , \_zy_simnet_tvar_20[4][241] , 
	\_zy_simnet_tvar_20[4][240] , \_zy_simnet_tvar_20[4][239] , 
	\_zy_simnet_tvar_20[4][238] , \_zy_simnet_tvar_20[4][237] , 
	\_zy_simnet_tvar_20[4][236] , \_zy_simnet_tvar_20[4][235] , 
	\_zy_simnet_tvar_20[4][234] , \_zy_simnet_tvar_20[4][233] , 
	\_zy_simnet_tvar_20[4][232] , \_zy_simnet_tvar_20[4][231] , 
	\_zy_simnet_tvar_20[4][230] , \_zy_simnet_tvar_20[4][229] , 
	\_zy_simnet_tvar_20[4][228] , \_zy_simnet_tvar_20[4][227] , 
	\_zy_simnet_tvar_20[4][226] , \_zy_simnet_tvar_20[4][225] , 
	\_zy_simnet_tvar_20[4][224] , \_zy_simnet_tvar_20[4][223] , 
	\_zy_simnet_tvar_20[4][222] , \_zy_simnet_tvar_20[4][221] , 
	\_zy_simnet_tvar_20[4][220] , \_zy_simnet_tvar_20[4][219] , 
	\_zy_simnet_tvar_20[4][218] , \_zy_simnet_tvar_20[4][217] , 
	\_zy_simnet_tvar_20[4][216] , \_zy_simnet_tvar_20[4][215] , 
	\_zy_simnet_tvar_20[4][214] , \_zy_simnet_tvar_20[4][213] , 
	\_zy_simnet_tvar_20[4][212] , \_zy_simnet_tvar_20[4][211] , 
	\_zy_simnet_tvar_20[4][210] , \_zy_simnet_tvar_20[4][209] , 
	\_zy_simnet_tvar_20[4][208] , \_zy_simnet_tvar_20[4][207] , 
	\_zy_simnet_tvar_20[4][206] , \_zy_simnet_tvar_20[4][205] , 
	\_zy_simnet_tvar_20[4][204] , \_zy_simnet_tvar_20[4][203] , 
	\_zy_simnet_tvar_20[4][202] , \_zy_simnet_tvar_20[4][201] , 
	\_zy_simnet_tvar_20[4][200] , \_zy_simnet_tvar_20[4][199] , 
	\_zy_simnet_tvar_20[4][198] , \_zy_simnet_tvar_20[4][197] , 
	\_zy_simnet_tvar_20[4][196] , \_zy_simnet_tvar_20[4][195] , 
	\_zy_simnet_tvar_20[4][194] , \_zy_simnet_tvar_20[4][193] , 
	\_zy_simnet_tvar_20[4][192] , \_zy_simnet_tvar_20[4][191] , 
	\_zy_simnet_tvar_20[4][190] , \_zy_simnet_tvar_20[4][189] , 
	\_zy_simnet_tvar_20[4][188] , \_zy_simnet_tvar_20[4][187] , 
	\_zy_simnet_tvar_20[4][186] , \_zy_simnet_tvar_20[4][185] , 
	\_zy_simnet_tvar_20[4][184] , \_zy_simnet_tvar_20[4][183] , 
	\_zy_simnet_tvar_20[4][182] , \_zy_simnet_tvar_20[4][181] , 
	\_zy_simnet_tvar_20[4][180] , \_zy_simnet_tvar_20[4][179] , 
	\_zy_simnet_tvar_20[4][178] , \_zy_simnet_tvar_20[4][177] , 
	\_zy_simnet_tvar_20[4][176] , \_zy_simnet_tvar_20[4][175] , 
	\_zy_simnet_tvar_20[4][174] , \_zy_simnet_tvar_20[4][173] , 
	\_zy_simnet_tvar_20[4][172] , \_zy_simnet_tvar_20[4][171] , 
	\_zy_simnet_tvar_20[4][170] , \_zy_simnet_tvar_20[4][169] , 
	\_zy_simnet_tvar_20[4][168] , \_zy_simnet_tvar_20[4][167] , 
	\_zy_simnet_tvar_20[4][166] , \_zy_simnet_tvar_20[4][165] , 
	\_zy_simnet_tvar_20[4][164] , \_zy_simnet_tvar_20[4][163] , 
	\_zy_simnet_tvar_20[4][162] , \_zy_simnet_tvar_20[4][161] , 
	\_zy_simnet_tvar_20[4][160] , \_zy_simnet_tvar_20[4][159] , 
	\_zy_simnet_tvar_20[4][158] , \_zy_simnet_tvar_20[4][157] , 
	\_zy_simnet_tvar_20[4][156] , \_zy_simnet_tvar_20[4][155] , 
	\_zy_simnet_tvar_20[4][154] , \_zy_simnet_tvar_20[4][153] , 
	\_zy_simnet_tvar_20[4][152] , \_zy_simnet_tvar_20[4][151] , 
	\_zy_simnet_tvar_20[4][150] , \_zy_simnet_tvar_20[4][149] , 
	\_zy_simnet_tvar_20[4][148] , \_zy_simnet_tvar_20[4][147] , 
	\_zy_simnet_tvar_20[4][146] , \_zy_simnet_tvar_20[4][145] , 
	\_zy_simnet_tvar_20[4][144] , \_zy_simnet_tvar_20[4][143] , 
	\_zy_simnet_tvar_20[4][142] , \_zy_simnet_tvar_20[4][141] , 
	\_zy_simnet_tvar_20[4][140] , \_zy_simnet_tvar_20[4][139] , 
	\_zy_simnet_tvar_20[4][138] , \_zy_simnet_tvar_20[4][137] , 
	\_zy_simnet_tvar_20[4][136] , \_zy_simnet_tvar_20[4][135] , 
	\_zy_simnet_tvar_20[4][134] , \_zy_simnet_tvar_20[4][133] , 
	\_zy_simnet_tvar_20[4][132] , \_zy_simnet_tvar_20[4][131] , 
	\_zy_simnet_tvar_20[4][130] , \_zy_simnet_tvar_20[4][129] , 
	\_zy_simnet_tvar_20[4][128] , \_zy_simnet_tvar_20[4][127] , 
	\_zy_simnet_tvar_20[4][126] , \_zy_simnet_tvar_20[4][125] , 
	\_zy_simnet_tvar_20[4][124] , \_zy_simnet_tvar_20[4][123] , 
	\_zy_simnet_tvar_20[4][122] , \_zy_simnet_tvar_20[4][121] , 
	\_zy_simnet_tvar_20[4][120] , \_zy_simnet_tvar_20[4][119] , 
	\_zy_simnet_tvar_20[4][118] , \_zy_simnet_tvar_20[4][117] , 
	\_zy_simnet_tvar_20[4][116] , \_zy_simnet_tvar_20[4][115] , 
	\_zy_simnet_tvar_20[4][114] , \_zy_simnet_tvar_20[4][113] , 
	\_zy_simnet_tvar_20[4][112] , \_zy_simnet_tvar_20[4][111] , 
	\_zy_simnet_tvar_20[4][110] , \_zy_simnet_tvar_20[4][109] , 
	\_zy_simnet_tvar_20[4][108] , \_zy_simnet_tvar_20[4][107] , 
	\_zy_simnet_tvar_20[4][106] , \_zy_simnet_tvar_20[4][105] , 
	\_zy_simnet_tvar_20[4][104] , \_zy_simnet_tvar_20[4][103] , 
	\_zy_simnet_tvar_20[4][102] , \_zy_simnet_tvar_20[4][101] , 
	\_zy_simnet_tvar_20[4][100] , \_zy_simnet_tvar_20[4][99] , 
	\_zy_simnet_tvar_20[4][98] , \_zy_simnet_tvar_20[4][97] , 
	\_zy_simnet_tvar_20[4][96] , \_zy_simnet_tvar_20[4][95] , 
	\_zy_simnet_tvar_20[4][94] , \_zy_simnet_tvar_20[4][93] , 
	\_zy_simnet_tvar_20[4][92] , \_zy_simnet_tvar_20[4][91] , 
	\_zy_simnet_tvar_20[4][90] , \_zy_simnet_tvar_20[4][89] , 
	\_zy_simnet_tvar_20[4][88] , \_zy_simnet_tvar_20[4][87] , 
	\_zy_simnet_tvar_20[4][86] , \_zy_simnet_tvar_20[4][85] , 
	\_zy_simnet_tvar_20[4][84] , \_zy_simnet_tvar_20[4][83] , 
	\_zy_simnet_tvar_20[4][82] , \_zy_simnet_tvar_20[4][81] , 
	\_zy_simnet_tvar_20[4][80] , \_zy_simnet_tvar_20[4][79] , 
	\_zy_simnet_tvar_20[4][78] , \_zy_simnet_tvar_20[4][77] , 
	\_zy_simnet_tvar_20[4][76] , \_zy_simnet_tvar_20[4][75] , 
	\_zy_simnet_tvar_20[4][74] , \_zy_simnet_tvar_20[4][73] , 
	\_zy_simnet_tvar_20[4][72] , \_zy_simnet_tvar_20[4][71] , 
	\_zy_simnet_tvar_20[4][70] , \_zy_simnet_tvar_20[4][69] , 
	\_zy_simnet_tvar_20[4][68] , \_zy_simnet_tvar_20[4][67] , 
	\_zy_simnet_tvar_20[4][66] , \_zy_simnet_tvar_20[4][65] , 
	\_zy_simnet_tvar_20[4][64] , \_zy_simnet_tvar_20[4][63] , 
	\_zy_simnet_tvar_20[4][62] , \_zy_simnet_tvar_20[4][61] , 
	\_zy_simnet_tvar_20[4][60] , \_zy_simnet_tvar_20[4][59] , 
	\_zy_simnet_tvar_20[4][58] , \_zy_simnet_tvar_20[4][57] , 
	\_zy_simnet_tvar_20[4][56] , \_zy_simnet_tvar_20[4][55] , 
	\_zy_simnet_tvar_20[4][54] , \_zy_simnet_tvar_20[4][53] , 
	\_zy_simnet_tvar_20[4][52] , \_zy_simnet_tvar_20[4][51] , 
	\_zy_simnet_tvar_20[4][50] , \_zy_simnet_tvar_20[4][49] , 
	\_zy_simnet_tvar_20[4][48] , \_zy_simnet_tvar_20[4][47] , 
	\_zy_simnet_tvar_20[4][46] , \_zy_simnet_tvar_20[4][45] , 
	\_zy_simnet_tvar_20[4][44] , \_zy_simnet_tvar_20[4][43] , 
	\_zy_simnet_tvar_20[4][42] , \_zy_simnet_tvar_20[4][41] , 
	\_zy_simnet_tvar_20[4][40] , \_zy_simnet_tvar_20[4][39] , 
	\_zy_simnet_tvar_20[4][38] , \_zy_simnet_tvar_20[4][37] , 
	\_zy_simnet_tvar_20[4][36] , \_zy_simnet_tvar_20[4][35] , 
	\_zy_simnet_tvar_20[4][34] , \_zy_simnet_tvar_20[4][33] , 
	\_zy_simnet_tvar_20[4][32] , \_zy_simnet_tvar_20[4][31] , 
	\_zy_simnet_tvar_20[4][30] , \_zy_simnet_tvar_20[4][29] , 
	\_zy_simnet_tvar_20[4][28] , \_zy_simnet_tvar_20[4][27] , 
	\_zy_simnet_tvar_20[4][26] , \_zy_simnet_tvar_20[4][25] , 
	\_zy_simnet_tvar_20[4][24] , \_zy_simnet_tvar_20[4][23] , 
	\_zy_simnet_tvar_20[4][22] , \_zy_simnet_tvar_20[4][21] , 
	\_zy_simnet_tvar_20[4][20] , \_zy_simnet_tvar_20[4][19] , 
	\_zy_simnet_tvar_20[4][18] , \_zy_simnet_tvar_20[4][17] , 
	\_zy_simnet_tvar_20[4][16] , \_zy_simnet_tvar_20[4][15] , 
	\_zy_simnet_tvar_20[4][14] , \_zy_simnet_tvar_20[4][13] , 
	\_zy_simnet_tvar_20[4][12] , \_zy_simnet_tvar_20[4][11] , 
	\_zy_simnet_tvar_20[4][10] , \_zy_simnet_tvar_20[4][9] , 
	\_zy_simnet_tvar_20[4][8] , \_zy_simnet_tvar_20[4][7] , 
	\_zy_simnet_tvar_20[4][6] , \_zy_simnet_tvar_20[4][5] , 
	\_zy_simnet_tvar_20[4][4] , \_zy_simnet_tvar_20[4][3] , 
	\_zy_simnet_tvar_20[4][2] , \_zy_simnet_tvar_20[4][1] , 
	\_zy_simnet_tvar_20[4][0] , \_zy_simnet_tvar_20[3][271] , 
	\_zy_simnet_tvar_20[3][270] , \_zy_simnet_tvar_20[3][269] , 
	\_zy_simnet_tvar_20[3][268] , \_zy_simnet_tvar_20[3][267] , 
	\_zy_simnet_tvar_20[3][266] , \_zy_simnet_tvar_20[3][265] , 
	\_zy_simnet_tvar_20[3][264] , \_zy_simnet_tvar_20[3][263] , 
	\_zy_simnet_tvar_20[3][262] , \_zy_simnet_tvar_20[3][261] , 
	\_zy_simnet_tvar_20[3][260] , \_zy_simnet_tvar_20[3][259] , 
	\_zy_simnet_tvar_20[3][258] , \_zy_simnet_tvar_20[3][257] , 
	\_zy_simnet_tvar_20[3][256] , \_zy_simnet_tvar_20[3][255] , 
	\_zy_simnet_tvar_20[3][254] , \_zy_simnet_tvar_20[3][253] , 
	\_zy_simnet_tvar_20[3][252] , \_zy_simnet_tvar_20[3][251] , 
	\_zy_simnet_tvar_20[3][250] , \_zy_simnet_tvar_20[3][249] , 
	\_zy_simnet_tvar_20[3][248] , \_zy_simnet_tvar_20[3][247] , 
	\_zy_simnet_tvar_20[3][246] , \_zy_simnet_tvar_20[3][245] , 
	\_zy_simnet_tvar_20[3][244] , \_zy_simnet_tvar_20[3][243] , 
	\_zy_simnet_tvar_20[3][242] , \_zy_simnet_tvar_20[3][241] , 
	\_zy_simnet_tvar_20[3][240] , \_zy_simnet_tvar_20[3][239] , 
	\_zy_simnet_tvar_20[3][238] , \_zy_simnet_tvar_20[3][237] , 
	\_zy_simnet_tvar_20[3][236] , \_zy_simnet_tvar_20[3][235] , 
	\_zy_simnet_tvar_20[3][234] , \_zy_simnet_tvar_20[3][233] , 
	\_zy_simnet_tvar_20[3][232] , \_zy_simnet_tvar_20[3][231] , 
	\_zy_simnet_tvar_20[3][230] , \_zy_simnet_tvar_20[3][229] , 
	\_zy_simnet_tvar_20[3][228] , \_zy_simnet_tvar_20[3][227] , 
	\_zy_simnet_tvar_20[3][226] , \_zy_simnet_tvar_20[3][225] , 
	\_zy_simnet_tvar_20[3][224] , \_zy_simnet_tvar_20[3][223] , 
	\_zy_simnet_tvar_20[3][222] , \_zy_simnet_tvar_20[3][221] , 
	\_zy_simnet_tvar_20[3][220] , \_zy_simnet_tvar_20[3][219] , 
	\_zy_simnet_tvar_20[3][218] , \_zy_simnet_tvar_20[3][217] , 
	\_zy_simnet_tvar_20[3][216] , \_zy_simnet_tvar_20[3][215] , 
	\_zy_simnet_tvar_20[3][214] , \_zy_simnet_tvar_20[3][213] , 
	\_zy_simnet_tvar_20[3][212] , \_zy_simnet_tvar_20[3][211] , 
	\_zy_simnet_tvar_20[3][210] , \_zy_simnet_tvar_20[3][209] , 
	\_zy_simnet_tvar_20[3][208] , \_zy_simnet_tvar_20[3][207] , 
	\_zy_simnet_tvar_20[3][206] , \_zy_simnet_tvar_20[3][205] , 
	\_zy_simnet_tvar_20[3][204] , \_zy_simnet_tvar_20[3][203] , 
	\_zy_simnet_tvar_20[3][202] , \_zy_simnet_tvar_20[3][201] , 
	\_zy_simnet_tvar_20[3][200] , \_zy_simnet_tvar_20[3][199] , 
	\_zy_simnet_tvar_20[3][198] , \_zy_simnet_tvar_20[3][197] , 
	\_zy_simnet_tvar_20[3][196] , \_zy_simnet_tvar_20[3][195] , 
	\_zy_simnet_tvar_20[3][194] , \_zy_simnet_tvar_20[3][193] , 
	\_zy_simnet_tvar_20[3][192] , \_zy_simnet_tvar_20[3][191] , 
	\_zy_simnet_tvar_20[3][190] , \_zy_simnet_tvar_20[3][189] , 
	\_zy_simnet_tvar_20[3][188] , \_zy_simnet_tvar_20[3][187] , 
	\_zy_simnet_tvar_20[3][186] , \_zy_simnet_tvar_20[3][185] , 
	\_zy_simnet_tvar_20[3][184] , \_zy_simnet_tvar_20[3][183] , 
	\_zy_simnet_tvar_20[3][182] , \_zy_simnet_tvar_20[3][181] , 
	\_zy_simnet_tvar_20[3][180] , \_zy_simnet_tvar_20[3][179] , 
	\_zy_simnet_tvar_20[3][178] , \_zy_simnet_tvar_20[3][177] , 
	\_zy_simnet_tvar_20[3][176] , \_zy_simnet_tvar_20[3][175] , 
	\_zy_simnet_tvar_20[3][174] , \_zy_simnet_tvar_20[3][173] , 
	\_zy_simnet_tvar_20[3][172] , \_zy_simnet_tvar_20[3][171] , 
	\_zy_simnet_tvar_20[3][170] , \_zy_simnet_tvar_20[3][169] , 
	\_zy_simnet_tvar_20[3][168] , \_zy_simnet_tvar_20[3][167] , 
	\_zy_simnet_tvar_20[3][166] , \_zy_simnet_tvar_20[3][165] , 
	\_zy_simnet_tvar_20[3][164] , \_zy_simnet_tvar_20[3][163] , 
	\_zy_simnet_tvar_20[3][162] , \_zy_simnet_tvar_20[3][161] , 
	\_zy_simnet_tvar_20[3][160] , \_zy_simnet_tvar_20[3][159] , 
	\_zy_simnet_tvar_20[3][158] , \_zy_simnet_tvar_20[3][157] , 
	\_zy_simnet_tvar_20[3][156] , \_zy_simnet_tvar_20[3][155] , 
	\_zy_simnet_tvar_20[3][154] , \_zy_simnet_tvar_20[3][153] , 
	\_zy_simnet_tvar_20[3][152] , \_zy_simnet_tvar_20[3][151] , 
	\_zy_simnet_tvar_20[3][150] , \_zy_simnet_tvar_20[3][149] , 
	\_zy_simnet_tvar_20[3][148] , \_zy_simnet_tvar_20[3][147] , 
	\_zy_simnet_tvar_20[3][146] , \_zy_simnet_tvar_20[3][145] , 
	\_zy_simnet_tvar_20[3][144] , \_zy_simnet_tvar_20[3][143] , 
	\_zy_simnet_tvar_20[3][142] , \_zy_simnet_tvar_20[3][141] , 
	\_zy_simnet_tvar_20[3][140] , \_zy_simnet_tvar_20[3][139] , 
	\_zy_simnet_tvar_20[3][138] , \_zy_simnet_tvar_20[3][137] , 
	\_zy_simnet_tvar_20[3][136] , \_zy_simnet_tvar_20[3][135] , 
	\_zy_simnet_tvar_20[3][134] , \_zy_simnet_tvar_20[3][133] , 
	\_zy_simnet_tvar_20[3][132] , \_zy_simnet_tvar_20[3][131] , 
	\_zy_simnet_tvar_20[3][130] , \_zy_simnet_tvar_20[3][129] , 
	\_zy_simnet_tvar_20[3][128] , \_zy_simnet_tvar_20[3][127] , 
	\_zy_simnet_tvar_20[3][126] , \_zy_simnet_tvar_20[3][125] , 
	\_zy_simnet_tvar_20[3][124] , \_zy_simnet_tvar_20[3][123] , 
	\_zy_simnet_tvar_20[3][122] , \_zy_simnet_tvar_20[3][121] , 
	\_zy_simnet_tvar_20[3][120] , \_zy_simnet_tvar_20[3][119] , 
	\_zy_simnet_tvar_20[3][118] , \_zy_simnet_tvar_20[3][117] , 
	\_zy_simnet_tvar_20[3][116] , \_zy_simnet_tvar_20[3][115] , 
	\_zy_simnet_tvar_20[3][114] , \_zy_simnet_tvar_20[3][113] , 
	\_zy_simnet_tvar_20[3][112] , \_zy_simnet_tvar_20[3][111] , 
	\_zy_simnet_tvar_20[3][110] , \_zy_simnet_tvar_20[3][109] , 
	\_zy_simnet_tvar_20[3][108] , \_zy_simnet_tvar_20[3][107] , 
	\_zy_simnet_tvar_20[3][106] , \_zy_simnet_tvar_20[3][105] , 
	\_zy_simnet_tvar_20[3][104] , \_zy_simnet_tvar_20[3][103] , 
	\_zy_simnet_tvar_20[3][102] , \_zy_simnet_tvar_20[3][101] , 
	\_zy_simnet_tvar_20[3][100] , \_zy_simnet_tvar_20[3][99] , 
	\_zy_simnet_tvar_20[3][98] , \_zy_simnet_tvar_20[3][97] , 
	\_zy_simnet_tvar_20[3][96] , \_zy_simnet_tvar_20[3][95] , 
	\_zy_simnet_tvar_20[3][94] , \_zy_simnet_tvar_20[3][93] , 
	\_zy_simnet_tvar_20[3][92] , \_zy_simnet_tvar_20[3][91] , 
	\_zy_simnet_tvar_20[3][90] , \_zy_simnet_tvar_20[3][89] , 
	\_zy_simnet_tvar_20[3][88] , \_zy_simnet_tvar_20[3][87] , 
	\_zy_simnet_tvar_20[3][86] , \_zy_simnet_tvar_20[3][85] , 
	\_zy_simnet_tvar_20[3][84] , \_zy_simnet_tvar_20[3][83] , 
	\_zy_simnet_tvar_20[3][82] , \_zy_simnet_tvar_20[3][81] , 
	\_zy_simnet_tvar_20[3][80] , \_zy_simnet_tvar_20[3][79] , 
	\_zy_simnet_tvar_20[3][78] , \_zy_simnet_tvar_20[3][77] , 
	\_zy_simnet_tvar_20[3][76] , \_zy_simnet_tvar_20[3][75] , 
	\_zy_simnet_tvar_20[3][74] , \_zy_simnet_tvar_20[3][73] , 
	\_zy_simnet_tvar_20[3][72] , \_zy_simnet_tvar_20[3][71] , 
	\_zy_simnet_tvar_20[3][70] , \_zy_simnet_tvar_20[3][69] , 
	\_zy_simnet_tvar_20[3][68] , \_zy_simnet_tvar_20[3][67] , 
	\_zy_simnet_tvar_20[3][66] , \_zy_simnet_tvar_20[3][65] , 
	\_zy_simnet_tvar_20[3][64] , \_zy_simnet_tvar_20[3][63] , 
	\_zy_simnet_tvar_20[3][62] , \_zy_simnet_tvar_20[3][61] , 
	\_zy_simnet_tvar_20[3][60] , \_zy_simnet_tvar_20[3][59] , 
	\_zy_simnet_tvar_20[3][58] , \_zy_simnet_tvar_20[3][57] , 
	\_zy_simnet_tvar_20[3][56] , \_zy_simnet_tvar_20[3][55] , 
	\_zy_simnet_tvar_20[3][54] , \_zy_simnet_tvar_20[3][53] , 
	\_zy_simnet_tvar_20[3][52] , \_zy_simnet_tvar_20[3][51] , 
	\_zy_simnet_tvar_20[3][50] , \_zy_simnet_tvar_20[3][49] , 
	\_zy_simnet_tvar_20[3][48] , \_zy_simnet_tvar_20[3][47] , 
	\_zy_simnet_tvar_20[3][46] , \_zy_simnet_tvar_20[3][45] , 
	\_zy_simnet_tvar_20[3][44] , \_zy_simnet_tvar_20[3][43] , 
	\_zy_simnet_tvar_20[3][42] , \_zy_simnet_tvar_20[3][41] , 
	\_zy_simnet_tvar_20[3][40] , \_zy_simnet_tvar_20[3][39] , 
	\_zy_simnet_tvar_20[3][38] , \_zy_simnet_tvar_20[3][37] , 
	\_zy_simnet_tvar_20[3][36] , \_zy_simnet_tvar_20[3][35] , 
	\_zy_simnet_tvar_20[3][34] , \_zy_simnet_tvar_20[3][33] , 
	\_zy_simnet_tvar_20[3][32] , \_zy_simnet_tvar_20[3][31] , 
	\_zy_simnet_tvar_20[3][30] , \_zy_simnet_tvar_20[3][29] , 
	\_zy_simnet_tvar_20[3][28] , \_zy_simnet_tvar_20[3][27] , 
	\_zy_simnet_tvar_20[3][26] , \_zy_simnet_tvar_20[3][25] , 
	\_zy_simnet_tvar_20[3][24] , \_zy_simnet_tvar_20[3][23] , 
	\_zy_simnet_tvar_20[3][22] , \_zy_simnet_tvar_20[3][21] , 
	\_zy_simnet_tvar_20[3][20] , \_zy_simnet_tvar_20[3][19] , 
	\_zy_simnet_tvar_20[3][18] , \_zy_simnet_tvar_20[3][17] , 
	\_zy_simnet_tvar_20[3][16] , \_zy_simnet_tvar_20[3][15] , 
	\_zy_simnet_tvar_20[3][14] , \_zy_simnet_tvar_20[3][13] , 
	\_zy_simnet_tvar_20[3][12] , \_zy_simnet_tvar_20[3][11] , 
	\_zy_simnet_tvar_20[3][10] , \_zy_simnet_tvar_20[3][9] , 
	\_zy_simnet_tvar_20[3][8] , \_zy_simnet_tvar_20[3][7] , 
	\_zy_simnet_tvar_20[3][6] , \_zy_simnet_tvar_20[3][5] , 
	\_zy_simnet_tvar_20[3][4] , \_zy_simnet_tvar_20[3][3] , 
	\_zy_simnet_tvar_20[3][2] , \_zy_simnet_tvar_20[3][1] , 
	\_zy_simnet_tvar_20[3][0] , \_zy_simnet_tvar_20[2][271] , 
	\_zy_simnet_tvar_20[2][270] , \_zy_simnet_tvar_20[2][269] , 
	\_zy_simnet_tvar_20[2][268] , \_zy_simnet_tvar_20[2][267] , 
	\_zy_simnet_tvar_20[2][266] , \_zy_simnet_tvar_20[2][265] , 
	\_zy_simnet_tvar_20[2][264] , \_zy_simnet_tvar_20[2][263] , 
	\_zy_simnet_tvar_20[2][262] , \_zy_simnet_tvar_20[2][261] , 
	\_zy_simnet_tvar_20[2][260] , \_zy_simnet_tvar_20[2][259] , 
	\_zy_simnet_tvar_20[2][258] , \_zy_simnet_tvar_20[2][257] , 
	\_zy_simnet_tvar_20[2][256] , \_zy_simnet_tvar_20[2][255] , 
	\_zy_simnet_tvar_20[2][254] , \_zy_simnet_tvar_20[2][253] , 
	\_zy_simnet_tvar_20[2][252] , \_zy_simnet_tvar_20[2][251] , 
	\_zy_simnet_tvar_20[2][250] , \_zy_simnet_tvar_20[2][249] , 
	\_zy_simnet_tvar_20[2][248] , \_zy_simnet_tvar_20[2][247] , 
	\_zy_simnet_tvar_20[2][246] , \_zy_simnet_tvar_20[2][245] , 
	\_zy_simnet_tvar_20[2][244] , \_zy_simnet_tvar_20[2][243] , 
	\_zy_simnet_tvar_20[2][242] , \_zy_simnet_tvar_20[2][241] , 
	\_zy_simnet_tvar_20[2][240] , \_zy_simnet_tvar_20[2][239] , 
	\_zy_simnet_tvar_20[2][238] , \_zy_simnet_tvar_20[2][237] , 
	\_zy_simnet_tvar_20[2][236] , \_zy_simnet_tvar_20[2][235] , 
	\_zy_simnet_tvar_20[2][234] , \_zy_simnet_tvar_20[2][233] , 
	\_zy_simnet_tvar_20[2][232] , \_zy_simnet_tvar_20[2][231] , 
	\_zy_simnet_tvar_20[2][230] , \_zy_simnet_tvar_20[2][229] , 
	\_zy_simnet_tvar_20[2][228] , \_zy_simnet_tvar_20[2][227] , 
	\_zy_simnet_tvar_20[2][226] , \_zy_simnet_tvar_20[2][225] , 
	\_zy_simnet_tvar_20[2][224] , \_zy_simnet_tvar_20[2][223] , 
	\_zy_simnet_tvar_20[2][222] , \_zy_simnet_tvar_20[2][221] , 
	\_zy_simnet_tvar_20[2][220] , \_zy_simnet_tvar_20[2][219] , 
	\_zy_simnet_tvar_20[2][218] , \_zy_simnet_tvar_20[2][217] , 
	\_zy_simnet_tvar_20[2][216] , \_zy_simnet_tvar_20[2][215] , 
	\_zy_simnet_tvar_20[2][214] , \_zy_simnet_tvar_20[2][213] , 
	\_zy_simnet_tvar_20[2][212] , \_zy_simnet_tvar_20[2][211] , 
	\_zy_simnet_tvar_20[2][210] , \_zy_simnet_tvar_20[2][209] , 
	\_zy_simnet_tvar_20[2][208] , \_zy_simnet_tvar_20[2][207] , 
	\_zy_simnet_tvar_20[2][206] , \_zy_simnet_tvar_20[2][205] , 
	\_zy_simnet_tvar_20[2][204] , \_zy_simnet_tvar_20[2][203] , 
	\_zy_simnet_tvar_20[2][202] , \_zy_simnet_tvar_20[2][201] , 
	\_zy_simnet_tvar_20[2][200] , \_zy_simnet_tvar_20[2][199] , 
	\_zy_simnet_tvar_20[2][198] , \_zy_simnet_tvar_20[2][197] , 
	\_zy_simnet_tvar_20[2][196] , \_zy_simnet_tvar_20[2][195] , 
	\_zy_simnet_tvar_20[2][194] , \_zy_simnet_tvar_20[2][193] , 
	\_zy_simnet_tvar_20[2][192] , \_zy_simnet_tvar_20[2][191] , 
	\_zy_simnet_tvar_20[2][190] , \_zy_simnet_tvar_20[2][189] , 
	\_zy_simnet_tvar_20[2][188] , \_zy_simnet_tvar_20[2][187] , 
	\_zy_simnet_tvar_20[2][186] , \_zy_simnet_tvar_20[2][185] , 
	\_zy_simnet_tvar_20[2][184] , \_zy_simnet_tvar_20[2][183] , 
	\_zy_simnet_tvar_20[2][182] , \_zy_simnet_tvar_20[2][181] , 
	\_zy_simnet_tvar_20[2][180] , \_zy_simnet_tvar_20[2][179] , 
	\_zy_simnet_tvar_20[2][178] , \_zy_simnet_tvar_20[2][177] , 
	\_zy_simnet_tvar_20[2][176] , \_zy_simnet_tvar_20[2][175] , 
	\_zy_simnet_tvar_20[2][174] , \_zy_simnet_tvar_20[2][173] , 
	\_zy_simnet_tvar_20[2][172] , \_zy_simnet_tvar_20[2][171] , 
	\_zy_simnet_tvar_20[2][170] , \_zy_simnet_tvar_20[2][169] , 
	\_zy_simnet_tvar_20[2][168] , \_zy_simnet_tvar_20[2][167] , 
	\_zy_simnet_tvar_20[2][166] , \_zy_simnet_tvar_20[2][165] , 
	\_zy_simnet_tvar_20[2][164] , \_zy_simnet_tvar_20[2][163] , 
	\_zy_simnet_tvar_20[2][162] , \_zy_simnet_tvar_20[2][161] , 
	\_zy_simnet_tvar_20[2][160] , \_zy_simnet_tvar_20[2][159] , 
	\_zy_simnet_tvar_20[2][158] , \_zy_simnet_tvar_20[2][157] , 
	\_zy_simnet_tvar_20[2][156] , \_zy_simnet_tvar_20[2][155] , 
	\_zy_simnet_tvar_20[2][154] , \_zy_simnet_tvar_20[2][153] , 
	\_zy_simnet_tvar_20[2][152] , \_zy_simnet_tvar_20[2][151] , 
	\_zy_simnet_tvar_20[2][150] , \_zy_simnet_tvar_20[2][149] , 
	\_zy_simnet_tvar_20[2][148] , \_zy_simnet_tvar_20[2][147] , 
	\_zy_simnet_tvar_20[2][146] , \_zy_simnet_tvar_20[2][145] , 
	\_zy_simnet_tvar_20[2][144] , \_zy_simnet_tvar_20[2][143] , 
	\_zy_simnet_tvar_20[2][142] , \_zy_simnet_tvar_20[2][141] , 
	\_zy_simnet_tvar_20[2][140] , \_zy_simnet_tvar_20[2][139] , 
	\_zy_simnet_tvar_20[2][138] , \_zy_simnet_tvar_20[2][137] , 
	\_zy_simnet_tvar_20[2][136] , \_zy_simnet_tvar_20[2][135] , 
	\_zy_simnet_tvar_20[2][134] , \_zy_simnet_tvar_20[2][133] , 
	\_zy_simnet_tvar_20[2][132] , \_zy_simnet_tvar_20[2][131] , 
	\_zy_simnet_tvar_20[2][130] , \_zy_simnet_tvar_20[2][129] , 
	\_zy_simnet_tvar_20[2][128] , \_zy_simnet_tvar_20[2][127] , 
	\_zy_simnet_tvar_20[2][126] , \_zy_simnet_tvar_20[2][125] , 
	\_zy_simnet_tvar_20[2][124] , \_zy_simnet_tvar_20[2][123] , 
	\_zy_simnet_tvar_20[2][122] , \_zy_simnet_tvar_20[2][121] , 
	\_zy_simnet_tvar_20[2][120] , \_zy_simnet_tvar_20[2][119] , 
	\_zy_simnet_tvar_20[2][118] , \_zy_simnet_tvar_20[2][117] , 
	\_zy_simnet_tvar_20[2][116] , \_zy_simnet_tvar_20[2][115] , 
	\_zy_simnet_tvar_20[2][114] , \_zy_simnet_tvar_20[2][113] , 
	\_zy_simnet_tvar_20[2][112] , \_zy_simnet_tvar_20[2][111] , 
	\_zy_simnet_tvar_20[2][110] , \_zy_simnet_tvar_20[2][109] , 
	\_zy_simnet_tvar_20[2][108] , \_zy_simnet_tvar_20[2][107] , 
	\_zy_simnet_tvar_20[2][106] , \_zy_simnet_tvar_20[2][105] , 
	\_zy_simnet_tvar_20[2][104] , \_zy_simnet_tvar_20[2][103] , 
	\_zy_simnet_tvar_20[2][102] , \_zy_simnet_tvar_20[2][101] , 
	\_zy_simnet_tvar_20[2][100] , \_zy_simnet_tvar_20[2][99] , 
	\_zy_simnet_tvar_20[2][98] , \_zy_simnet_tvar_20[2][97] , 
	\_zy_simnet_tvar_20[2][96] , \_zy_simnet_tvar_20[2][95] , 
	\_zy_simnet_tvar_20[2][94] , \_zy_simnet_tvar_20[2][93] , 
	\_zy_simnet_tvar_20[2][92] , \_zy_simnet_tvar_20[2][91] , 
	\_zy_simnet_tvar_20[2][90] , \_zy_simnet_tvar_20[2][89] , 
	\_zy_simnet_tvar_20[2][88] , \_zy_simnet_tvar_20[2][87] , 
	\_zy_simnet_tvar_20[2][86] , \_zy_simnet_tvar_20[2][85] , 
	\_zy_simnet_tvar_20[2][84] , \_zy_simnet_tvar_20[2][83] , 
	\_zy_simnet_tvar_20[2][82] , \_zy_simnet_tvar_20[2][81] , 
	\_zy_simnet_tvar_20[2][80] , \_zy_simnet_tvar_20[2][79] , 
	\_zy_simnet_tvar_20[2][78] , \_zy_simnet_tvar_20[2][77] , 
	\_zy_simnet_tvar_20[2][76] , \_zy_simnet_tvar_20[2][75] , 
	\_zy_simnet_tvar_20[2][74] , \_zy_simnet_tvar_20[2][73] , 
	\_zy_simnet_tvar_20[2][72] , \_zy_simnet_tvar_20[2][71] , 
	\_zy_simnet_tvar_20[2][70] , \_zy_simnet_tvar_20[2][69] , 
	\_zy_simnet_tvar_20[2][68] , \_zy_simnet_tvar_20[2][67] , 
	\_zy_simnet_tvar_20[2][66] , \_zy_simnet_tvar_20[2][65] , 
	\_zy_simnet_tvar_20[2][64] , \_zy_simnet_tvar_20[2][63] , 
	\_zy_simnet_tvar_20[2][62] , \_zy_simnet_tvar_20[2][61] , 
	\_zy_simnet_tvar_20[2][60] , \_zy_simnet_tvar_20[2][59] , 
	\_zy_simnet_tvar_20[2][58] , \_zy_simnet_tvar_20[2][57] , 
	\_zy_simnet_tvar_20[2][56] , \_zy_simnet_tvar_20[2][55] , 
	\_zy_simnet_tvar_20[2][54] , \_zy_simnet_tvar_20[2][53] , 
	\_zy_simnet_tvar_20[2][52] , \_zy_simnet_tvar_20[2][51] , 
	\_zy_simnet_tvar_20[2][50] , \_zy_simnet_tvar_20[2][49] , 
	\_zy_simnet_tvar_20[2][48] , \_zy_simnet_tvar_20[2][47] , 
	\_zy_simnet_tvar_20[2][46] , \_zy_simnet_tvar_20[2][45] , 
	\_zy_simnet_tvar_20[2][44] , \_zy_simnet_tvar_20[2][43] , 
	\_zy_simnet_tvar_20[2][42] , \_zy_simnet_tvar_20[2][41] , 
	\_zy_simnet_tvar_20[2][40] , \_zy_simnet_tvar_20[2][39] , 
	\_zy_simnet_tvar_20[2][38] , \_zy_simnet_tvar_20[2][37] , 
	\_zy_simnet_tvar_20[2][36] , \_zy_simnet_tvar_20[2][35] , 
	\_zy_simnet_tvar_20[2][34] , \_zy_simnet_tvar_20[2][33] , 
	\_zy_simnet_tvar_20[2][32] , \_zy_simnet_tvar_20[2][31] , 
	\_zy_simnet_tvar_20[2][30] , \_zy_simnet_tvar_20[2][29] , 
	\_zy_simnet_tvar_20[2][28] , \_zy_simnet_tvar_20[2][27] , 
	\_zy_simnet_tvar_20[2][26] , \_zy_simnet_tvar_20[2][25] , 
	\_zy_simnet_tvar_20[2][24] , \_zy_simnet_tvar_20[2][23] , 
	\_zy_simnet_tvar_20[2][22] , \_zy_simnet_tvar_20[2][21] , 
	\_zy_simnet_tvar_20[2][20] , \_zy_simnet_tvar_20[2][19] , 
	\_zy_simnet_tvar_20[2][18] , \_zy_simnet_tvar_20[2][17] , 
	\_zy_simnet_tvar_20[2][16] , \_zy_simnet_tvar_20[2][15] , 
	\_zy_simnet_tvar_20[2][14] , \_zy_simnet_tvar_20[2][13] , 
	\_zy_simnet_tvar_20[2][12] , \_zy_simnet_tvar_20[2][11] , 
	\_zy_simnet_tvar_20[2][10] , \_zy_simnet_tvar_20[2][9] , 
	\_zy_simnet_tvar_20[2][8] , \_zy_simnet_tvar_20[2][7] , 
	\_zy_simnet_tvar_20[2][6] , \_zy_simnet_tvar_20[2][5] , 
	\_zy_simnet_tvar_20[2][4] , \_zy_simnet_tvar_20[2][3] , 
	\_zy_simnet_tvar_20[2][2] , \_zy_simnet_tvar_20[2][1] , 
	\_zy_simnet_tvar_20[2][0] , \_zy_simnet_tvar_20[1][271] , 
	\_zy_simnet_tvar_20[1][270] , \_zy_simnet_tvar_20[1][269] , 
	\_zy_simnet_tvar_20[1][268] , \_zy_simnet_tvar_20[1][267] , 
	\_zy_simnet_tvar_20[1][266] , \_zy_simnet_tvar_20[1][265] , 
	\_zy_simnet_tvar_20[1][264] , \_zy_simnet_tvar_20[1][263] , 
	\_zy_simnet_tvar_20[1][262] , \_zy_simnet_tvar_20[1][261] , 
	\_zy_simnet_tvar_20[1][260] , \_zy_simnet_tvar_20[1][259] , 
	\_zy_simnet_tvar_20[1][258] , \_zy_simnet_tvar_20[1][257] , 
	\_zy_simnet_tvar_20[1][256] , \_zy_simnet_tvar_20[1][255] , 
	\_zy_simnet_tvar_20[1][254] , \_zy_simnet_tvar_20[1][253] , 
	\_zy_simnet_tvar_20[1][252] , \_zy_simnet_tvar_20[1][251] , 
	\_zy_simnet_tvar_20[1][250] , \_zy_simnet_tvar_20[1][249] , 
	\_zy_simnet_tvar_20[1][248] , \_zy_simnet_tvar_20[1][247] , 
	\_zy_simnet_tvar_20[1][246] , \_zy_simnet_tvar_20[1][245] , 
	\_zy_simnet_tvar_20[1][244] , \_zy_simnet_tvar_20[1][243] , 
	\_zy_simnet_tvar_20[1][242] , \_zy_simnet_tvar_20[1][241] , 
	\_zy_simnet_tvar_20[1][240] , \_zy_simnet_tvar_20[1][239] , 
	\_zy_simnet_tvar_20[1][238] , \_zy_simnet_tvar_20[1][237] , 
	\_zy_simnet_tvar_20[1][236] , \_zy_simnet_tvar_20[1][235] , 
	\_zy_simnet_tvar_20[1][234] , \_zy_simnet_tvar_20[1][233] , 
	\_zy_simnet_tvar_20[1][232] , \_zy_simnet_tvar_20[1][231] , 
	\_zy_simnet_tvar_20[1][230] , \_zy_simnet_tvar_20[1][229] , 
	\_zy_simnet_tvar_20[1][228] , \_zy_simnet_tvar_20[1][227] , 
	\_zy_simnet_tvar_20[1][226] , \_zy_simnet_tvar_20[1][225] , 
	\_zy_simnet_tvar_20[1][224] , \_zy_simnet_tvar_20[1][223] , 
	\_zy_simnet_tvar_20[1][222] , \_zy_simnet_tvar_20[1][221] , 
	\_zy_simnet_tvar_20[1][220] , \_zy_simnet_tvar_20[1][219] , 
	\_zy_simnet_tvar_20[1][218] , \_zy_simnet_tvar_20[1][217] , 
	\_zy_simnet_tvar_20[1][216] , \_zy_simnet_tvar_20[1][215] , 
	\_zy_simnet_tvar_20[1][214] , \_zy_simnet_tvar_20[1][213] , 
	\_zy_simnet_tvar_20[1][212] , \_zy_simnet_tvar_20[1][211] , 
	\_zy_simnet_tvar_20[1][210] , \_zy_simnet_tvar_20[1][209] , 
	\_zy_simnet_tvar_20[1][208] , \_zy_simnet_tvar_20[1][207] , 
	\_zy_simnet_tvar_20[1][206] , \_zy_simnet_tvar_20[1][205] , 
	\_zy_simnet_tvar_20[1][204] , \_zy_simnet_tvar_20[1][203] , 
	\_zy_simnet_tvar_20[1][202] , \_zy_simnet_tvar_20[1][201] , 
	\_zy_simnet_tvar_20[1][200] , \_zy_simnet_tvar_20[1][199] , 
	\_zy_simnet_tvar_20[1][198] , \_zy_simnet_tvar_20[1][197] , 
	\_zy_simnet_tvar_20[1][196] , \_zy_simnet_tvar_20[1][195] , 
	\_zy_simnet_tvar_20[1][194] , \_zy_simnet_tvar_20[1][193] , 
	\_zy_simnet_tvar_20[1][192] , \_zy_simnet_tvar_20[1][191] , 
	\_zy_simnet_tvar_20[1][190] , \_zy_simnet_tvar_20[1][189] , 
	\_zy_simnet_tvar_20[1][188] , \_zy_simnet_tvar_20[1][187] , 
	\_zy_simnet_tvar_20[1][186] , \_zy_simnet_tvar_20[1][185] , 
	\_zy_simnet_tvar_20[1][184] , \_zy_simnet_tvar_20[1][183] , 
	\_zy_simnet_tvar_20[1][182] , \_zy_simnet_tvar_20[1][181] , 
	\_zy_simnet_tvar_20[1][180] , \_zy_simnet_tvar_20[1][179] , 
	\_zy_simnet_tvar_20[1][178] , \_zy_simnet_tvar_20[1][177] , 
	\_zy_simnet_tvar_20[1][176] , \_zy_simnet_tvar_20[1][175] , 
	\_zy_simnet_tvar_20[1][174] , \_zy_simnet_tvar_20[1][173] , 
	\_zy_simnet_tvar_20[1][172] , \_zy_simnet_tvar_20[1][171] , 
	\_zy_simnet_tvar_20[1][170] , \_zy_simnet_tvar_20[1][169] , 
	\_zy_simnet_tvar_20[1][168] , \_zy_simnet_tvar_20[1][167] , 
	\_zy_simnet_tvar_20[1][166] , \_zy_simnet_tvar_20[1][165] , 
	\_zy_simnet_tvar_20[1][164] , \_zy_simnet_tvar_20[1][163] , 
	\_zy_simnet_tvar_20[1][162] , \_zy_simnet_tvar_20[1][161] , 
	\_zy_simnet_tvar_20[1][160] , \_zy_simnet_tvar_20[1][159] , 
	\_zy_simnet_tvar_20[1][158] , \_zy_simnet_tvar_20[1][157] , 
	\_zy_simnet_tvar_20[1][156] , \_zy_simnet_tvar_20[1][155] , 
	\_zy_simnet_tvar_20[1][154] , \_zy_simnet_tvar_20[1][153] , 
	\_zy_simnet_tvar_20[1][152] , \_zy_simnet_tvar_20[1][151] , 
	\_zy_simnet_tvar_20[1][150] , \_zy_simnet_tvar_20[1][149] , 
	\_zy_simnet_tvar_20[1][148] , \_zy_simnet_tvar_20[1][147] , 
	\_zy_simnet_tvar_20[1][146] , \_zy_simnet_tvar_20[1][145] , 
	\_zy_simnet_tvar_20[1][144] , \_zy_simnet_tvar_20[1][143] , 
	\_zy_simnet_tvar_20[1][142] , \_zy_simnet_tvar_20[1][141] , 
	\_zy_simnet_tvar_20[1][140] , \_zy_simnet_tvar_20[1][139] , 
	\_zy_simnet_tvar_20[1][138] , \_zy_simnet_tvar_20[1][137] , 
	\_zy_simnet_tvar_20[1][136] , \_zy_simnet_tvar_20[1][135] , 
	\_zy_simnet_tvar_20[1][134] , \_zy_simnet_tvar_20[1][133] , 
	\_zy_simnet_tvar_20[1][132] , \_zy_simnet_tvar_20[1][131] , 
	\_zy_simnet_tvar_20[1][130] , \_zy_simnet_tvar_20[1][129] , 
	\_zy_simnet_tvar_20[1][128] , \_zy_simnet_tvar_20[1][127] , 
	\_zy_simnet_tvar_20[1][126] , \_zy_simnet_tvar_20[1][125] , 
	\_zy_simnet_tvar_20[1][124] , \_zy_simnet_tvar_20[1][123] , 
	\_zy_simnet_tvar_20[1][122] , \_zy_simnet_tvar_20[1][121] , 
	\_zy_simnet_tvar_20[1][120] , \_zy_simnet_tvar_20[1][119] , 
	\_zy_simnet_tvar_20[1][118] , \_zy_simnet_tvar_20[1][117] , 
	\_zy_simnet_tvar_20[1][116] , \_zy_simnet_tvar_20[1][115] , 
	\_zy_simnet_tvar_20[1][114] , \_zy_simnet_tvar_20[1][113] , 
	\_zy_simnet_tvar_20[1][112] , \_zy_simnet_tvar_20[1][111] , 
	\_zy_simnet_tvar_20[1][110] , \_zy_simnet_tvar_20[1][109] , 
	\_zy_simnet_tvar_20[1][108] , \_zy_simnet_tvar_20[1][107] , 
	\_zy_simnet_tvar_20[1][106] , \_zy_simnet_tvar_20[1][105] , 
	\_zy_simnet_tvar_20[1][104] , \_zy_simnet_tvar_20[1][103] , 
	\_zy_simnet_tvar_20[1][102] , \_zy_simnet_tvar_20[1][101] , 
	\_zy_simnet_tvar_20[1][100] , \_zy_simnet_tvar_20[1][99] , 
	\_zy_simnet_tvar_20[1][98] , \_zy_simnet_tvar_20[1][97] , 
	\_zy_simnet_tvar_20[1][96] , \_zy_simnet_tvar_20[1][95] , 
	\_zy_simnet_tvar_20[1][94] , \_zy_simnet_tvar_20[1][93] , 
	\_zy_simnet_tvar_20[1][92] , \_zy_simnet_tvar_20[1][91] , 
	\_zy_simnet_tvar_20[1][90] , \_zy_simnet_tvar_20[1][89] , 
	\_zy_simnet_tvar_20[1][88] , \_zy_simnet_tvar_20[1][87] , 
	\_zy_simnet_tvar_20[1][86] , \_zy_simnet_tvar_20[1][85] , 
	\_zy_simnet_tvar_20[1][84] , \_zy_simnet_tvar_20[1][83] , 
	\_zy_simnet_tvar_20[1][82] , \_zy_simnet_tvar_20[1][81] , 
	\_zy_simnet_tvar_20[1][80] , \_zy_simnet_tvar_20[1][79] , 
	\_zy_simnet_tvar_20[1][78] , \_zy_simnet_tvar_20[1][77] , 
	\_zy_simnet_tvar_20[1][76] , \_zy_simnet_tvar_20[1][75] , 
	\_zy_simnet_tvar_20[1][74] , \_zy_simnet_tvar_20[1][73] , 
	\_zy_simnet_tvar_20[1][72] , \_zy_simnet_tvar_20[1][71] , 
	\_zy_simnet_tvar_20[1][70] , \_zy_simnet_tvar_20[1][69] , 
	\_zy_simnet_tvar_20[1][68] , \_zy_simnet_tvar_20[1][67] , 
	\_zy_simnet_tvar_20[1][66] , \_zy_simnet_tvar_20[1][65] , 
	\_zy_simnet_tvar_20[1][64] , \_zy_simnet_tvar_20[1][63] , 
	\_zy_simnet_tvar_20[1][62] , \_zy_simnet_tvar_20[1][61] , 
	\_zy_simnet_tvar_20[1][60] , \_zy_simnet_tvar_20[1][59] , 
	\_zy_simnet_tvar_20[1][58] , \_zy_simnet_tvar_20[1][57] , 
	\_zy_simnet_tvar_20[1][56] , \_zy_simnet_tvar_20[1][55] , 
	\_zy_simnet_tvar_20[1][54] , \_zy_simnet_tvar_20[1][53] , 
	\_zy_simnet_tvar_20[1][52] , \_zy_simnet_tvar_20[1][51] , 
	\_zy_simnet_tvar_20[1][50] , \_zy_simnet_tvar_20[1][49] , 
	\_zy_simnet_tvar_20[1][48] , \_zy_simnet_tvar_20[1][47] , 
	\_zy_simnet_tvar_20[1][46] , \_zy_simnet_tvar_20[1][45] , 
	\_zy_simnet_tvar_20[1][44] , \_zy_simnet_tvar_20[1][43] , 
	\_zy_simnet_tvar_20[1][42] , \_zy_simnet_tvar_20[1][41] , 
	\_zy_simnet_tvar_20[1][40] , \_zy_simnet_tvar_20[1][39] , 
	\_zy_simnet_tvar_20[1][38] , \_zy_simnet_tvar_20[1][37] , 
	\_zy_simnet_tvar_20[1][36] , \_zy_simnet_tvar_20[1][35] , 
	\_zy_simnet_tvar_20[1][34] , \_zy_simnet_tvar_20[1][33] , 
	\_zy_simnet_tvar_20[1][32] , \_zy_simnet_tvar_20[1][31] , 
	\_zy_simnet_tvar_20[1][30] , \_zy_simnet_tvar_20[1][29] , 
	\_zy_simnet_tvar_20[1][28] , \_zy_simnet_tvar_20[1][27] , 
	\_zy_simnet_tvar_20[1][26] , \_zy_simnet_tvar_20[1][25] , 
	\_zy_simnet_tvar_20[1][24] , \_zy_simnet_tvar_20[1][23] , 
	\_zy_simnet_tvar_20[1][22] , \_zy_simnet_tvar_20[1][21] , 
	\_zy_simnet_tvar_20[1][20] , \_zy_simnet_tvar_20[1][19] , 
	\_zy_simnet_tvar_20[1][18] , \_zy_simnet_tvar_20[1][17] , 
	\_zy_simnet_tvar_20[1][16] , \_zy_simnet_tvar_20[1][15] , 
	\_zy_simnet_tvar_20[1][14] , \_zy_simnet_tvar_20[1][13] , 
	\_zy_simnet_tvar_20[1][12] , \_zy_simnet_tvar_20[1][11] , 
	\_zy_simnet_tvar_20[1][10] , \_zy_simnet_tvar_20[1][9] , 
	\_zy_simnet_tvar_20[1][8] , \_zy_simnet_tvar_20[1][7] , 
	\_zy_simnet_tvar_20[1][6] , \_zy_simnet_tvar_20[1][5] , 
	\_zy_simnet_tvar_20[1][4] , \_zy_simnet_tvar_20[1][3] , 
	\_zy_simnet_tvar_20[1][2] , \_zy_simnet_tvar_20[1][1] , 
	\_zy_simnet_tvar_20[1][0] , \_zy_simnet_tvar_20[0][271] , 
	\_zy_simnet_tvar_20[0][270] , \_zy_simnet_tvar_20[0][269] , 
	\_zy_simnet_tvar_20[0][268] , \_zy_simnet_tvar_20[0][267] , 
	\_zy_simnet_tvar_20[0][266] , \_zy_simnet_tvar_20[0][265] , 
	\_zy_simnet_tvar_20[0][264] , \_zy_simnet_tvar_20[0][263] , 
	\_zy_simnet_tvar_20[0][262] , \_zy_simnet_tvar_20[0][261] , 
	\_zy_simnet_tvar_20[0][260] , \_zy_simnet_tvar_20[0][259] , 
	\_zy_simnet_tvar_20[0][258] , \_zy_simnet_tvar_20[0][257] , 
	\_zy_simnet_tvar_20[0][256] , \_zy_simnet_tvar_20[0][255] , 
	\_zy_simnet_tvar_20[0][254] , \_zy_simnet_tvar_20[0][253] , 
	\_zy_simnet_tvar_20[0][252] , \_zy_simnet_tvar_20[0][251] , 
	\_zy_simnet_tvar_20[0][250] , \_zy_simnet_tvar_20[0][249] , 
	\_zy_simnet_tvar_20[0][248] , \_zy_simnet_tvar_20[0][247] , 
	\_zy_simnet_tvar_20[0][246] , \_zy_simnet_tvar_20[0][245] , 
	\_zy_simnet_tvar_20[0][244] , \_zy_simnet_tvar_20[0][243] , 
	\_zy_simnet_tvar_20[0][242] , \_zy_simnet_tvar_20[0][241] , 
	\_zy_simnet_tvar_20[0][240] , \_zy_simnet_tvar_20[0][239] , 
	\_zy_simnet_tvar_20[0][238] , \_zy_simnet_tvar_20[0][237] , 
	\_zy_simnet_tvar_20[0][236] , \_zy_simnet_tvar_20[0][235] , 
	\_zy_simnet_tvar_20[0][234] , \_zy_simnet_tvar_20[0][233] , 
	\_zy_simnet_tvar_20[0][232] , \_zy_simnet_tvar_20[0][231] , 
	\_zy_simnet_tvar_20[0][230] , \_zy_simnet_tvar_20[0][229] , 
	\_zy_simnet_tvar_20[0][228] , \_zy_simnet_tvar_20[0][227] , 
	\_zy_simnet_tvar_20[0][226] , \_zy_simnet_tvar_20[0][225] , 
	\_zy_simnet_tvar_20[0][224] , \_zy_simnet_tvar_20[0][223] , 
	\_zy_simnet_tvar_20[0][222] , \_zy_simnet_tvar_20[0][221] , 
	\_zy_simnet_tvar_20[0][220] , \_zy_simnet_tvar_20[0][219] , 
	\_zy_simnet_tvar_20[0][218] , \_zy_simnet_tvar_20[0][217] , 
	\_zy_simnet_tvar_20[0][216] , \_zy_simnet_tvar_20[0][215] , 
	\_zy_simnet_tvar_20[0][214] , \_zy_simnet_tvar_20[0][213] , 
	\_zy_simnet_tvar_20[0][212] , \_zy_simnet_tvar_20[0][211] , 
	\_zy_simnet_tvar_20[0][210] , \_zy_simnet_tvar_20[0][209] , 
	\_zy_simnet_tvar_20[0][208] , \_zy_simnet_tvar_20[0][207] , 
	\_zy_simnet_tvar_20[0][206] , \_zy_simnet_tvar_20[0][205] , 
	\_zy_simnet_tvar_20[0][204] , \_zy_simnet_tvar_20[0][203] , 
	\_zy_simnet_tvar_20[0][202] , \_zy_simnet_tvar_20[0][201] , 
	\_zy_simnet_tvar_20[0][200] , \_zy_simnet_tvar_20[0][199] , 
	\_zy_simnet_tvar_20[0][198] , \_zy_simnet_tvar_20[0][197] , 
	\_zy_simnet_tvar_20[0][196] , \_zy_simnet_tvar_20[0][195] , 
	\_zy_simnet_tvar_20[0][194] , \_zy_simnet_tvar_20[0][193] , 
	\_zy_simnet_tvar_20[0][192] , \_zy_simnet_tvar_20[0][191] , 
	\_zy_simnet_tvar_20[0][190] , \_zy_simnet_tvar_20[0][189] , 
	\_zy_simnet_tvar_20[0][188] , \_zy_simnet_tvar_20[0][187] , 
	\_zy_simnet_tvar_20[0][186] , \_zy_simnet_tvar_20[0][185] , 
	\_zy_simnet_tvar_20[0][184] , \_zy_simnet_tvar_20[0][183] , 
	\_zy_simnet_tvar_20[0][182] , \_zy_simnet_tvar_20[0][181] , 
	\_zy_simnet_tvar_20[0][180] , \_zy_simnet_tvar_20[0][179] , 
	\_zy_simnet_tvar_20[0][178] , \_zy_simnet_tvar_20[0][177] , 
	\_zy_simnet_tvar_20[0][176] , \_zy_simnet_tvar_20[0][175] , 
	\_zy_simnet_tvar_20[0][174] , \_zy_simnet_tvar_20[0][173] , 
	\_zy_simnet_tvar_20[0][172] , \_zy_simnet_tvar_20[0][171] , 
	\_zy_simnet_tvar_20[0][170] , \_zy_simnet_tvar_20[0][169] , 
	\_zy_simnet_tvar_20[0][168] , \_zy_simnet_tvar_20[0][167] , 
	\_zy_simnet_tvar_20[0][166] , \_zy_simnet_tvar_20[0][165] , 
	\_zy_simnet_tvar_20[0][164] , \_zy_simnet_tvar_20[0][163] , 
	\_zy_simnet_tvar_20[0][162] , \_zy_simnet_tvar_20[0][161] , 
	\_zy_simnet_tvar_20[0][160] , \_zy_simnet_tvar_20[0][159] , 
	\_zy_simnet_tvar_20[0][158] , \_zy_simnet_tvar_20[0][157] , 
	\_zy_simnet_tvar_20[0][156] , \_zy_simnet_tvar_20[0][155] , 
	\_zy_simnet_tvar_20[0][154] , \_zy_simnet_tvar_20[0][153] , 
	\_zy_simnet_tvar_20[0][152] , \_zy_simnet_tvar_20[0][151] , 
	\_zy_simnet_tvar_20[0][150] , \_zy_simnet_tvar_20[0][149] , 
	\_zy_simnet_tvar_20[0][148] , \_zy_simnet_tvar_20[0][147] , 
	\_zy_simnet_tvar_20[0][146] , \_zy_simnet_tvar_20[0][145] , 
	\_zy_simnet_tvar_20[0][144] , \_zy_simnet_tvar_20[0][143] , 
	\_zy_simnet_tvar_20[0][142] , \_zy_simnet_tvar_20[0][141] , 
	\_zy_simnet_tvar_20[0][140] , \_zy_simnet_tvar_20[0][139] , 
	\_zy_simnet_tvar_20[0][138] , \_zy_simnet_tvar_20[0][137] , 
	\_zy_simnet_tvar_20[0][136] , \_zy_simnet_tvar_20[0][135] , 
	\_zy_simnet_tvar_20[0][134] , \_zy_simnet_tvar_20[0][133] , 
	\_zy_simnet_tvar_20[0][132] , \_zy_simnet_tvar_20[0][131] , 
	\_zy_simnet_tvar_20[0][130] , \_zy_simnet_tvar_20[0][129] , 
	\_zy_simnet_tvar_20[0][128] , \_zy_simnet_tvar_20[0][127] , 
	\_zy_simnet_tvar_20[0][126] , \_zy_simnet_tvar_20[0][125] , 
	\_zy_simnet_tvar_20[0][124] , \_zy_simnet_tvar_20[0][123] , 
	\_zy_simnet_tvar_20[0][122] , \_zy_simnet_tvar_20[0][121] , 
	\_zy_simnet_tvar_20[0][120] , \_zy_simnet_tvar_20[0][119] , 
	\_zy_simnet_tvar_20[0][118] , \_zy_simnet_tvar_20[0][117] , 
	\_zy_simnet_tvar_20[0][116] , \_zy_simnet_tvar_20[0][115] , 
	\_zy_simnet_tvar_20[0][114] , \_zy_simnet_tvar_20[0][113] , 
	\_zy_simnet_tvar_20[0][112] , \_zy_simnet_tvar_20[0][111] , 
	\_zy_simnet_tvar_20[0][110] , \_zy_simnet_tvar_20[0][109] , 
	\_zy_simnet_tvar_20[0][108] , \_zy_simnet_tvar_20[0][107] , 
	\_zy_simnet_tvar_20[0][106] , \_zy_simnet_tvar_20[0][105] , 
	\_zy_simnet_tvar_20[0][104] , \_zy_simnet_tvar_20[0][103] , 
	\_zy_simnet_tvar_20[0][102] , \_zy_simnet_tvar_20[0][101] , 
	\_zy_simnet_tvar_20[0][100] , \_zy_simnet_tvar_20[0][99] , 
	\_zy_simnet_tvar_20[0][98] , \_zy_simnet_tvar_20[0][97] , 
	\_zy_simnet_tvar_20[0][96] , \_zy_simnet_tvar_20[0][95] , 
	\_zy_simnet_tvar_20[0][94] , \_zy_simnet_tvar_20[0][93] , 
	\_zy_simnet_tvar_20[0][92] , \_zy_simnet_tvar_20[0][91] , 
	\_zy_simnet_tvar_20[0][90] , \_zy_simnet_tvar_20[0][89] , 
	\_zy_simnet_tvar_20[0][88] , \_zy_simnet_tvar_20[0][87] , 
	\_zy_simnet_tvar_20[0][86] , \_zy_simnet_tvar_20[0][85] , 
	\_zy_simnet_tvar_20[0][84] , \_zy_simnet_tvar_20[0][83] , 
	\_zy_simnet_tvar_20[0][82] , \_zy_simnet_tvar_20[0][81] , 
	\_zy_simnet_tvar_20[0][80] , \_zy_simnet_tvar_20[0][79] , 
	\_zy_simnet_tvar_20[0][78] , \_zy_simnet_tvar_20[0][77] , 
	\_zy_simnet_tvar_20[0][76] , \_zy_simnet_tvar_20[0][75] , 
	\_zy_simnet_tvar_20[0][74] , \_zy_simnet_tvar_20[0][73] , 
	\_zy_simnet_tvar_20[0][72] , \_zy_simnet_tvar_20[0][71] , 
	\_zy_simnet_tvar_20[0][70] , \_zy_simnet_tvar_20[0][69] , 
	\_zy_simnet_tvar_20[0][68] , \_zy_simnet_tvar_20[0][67] , 
	\_zy_simnet_tvar_20[0][66] , \_zy_simnet_tvar_20[0][65] , 
	\_zy_simnet_tvar_20[0][64] , \_zy_simnet_tvar_20[0][63] , 
	\_zy_simnet_tvar_20[0][62] , \_zy_simnet_tvar_20[0][61] , 
	\_zy_simnet_tvar_20[0][60] , \_zy_simnet_tvar_20[0][59] , 
	\_zy_simnet_tvar_20[0][58] , \_zy_simnet_tvar_20[0][57] , 
	\_zy_simnet_tvar_20[0][56] , \_zy_simnet_tvar_20[0][55] , 
	\_zy_simnet_tvar_20[0][54] , \_zy_simnet_tvar_20[0][53] , 
	\_zy_simnet_tvar_20[0][52] , \_zy_simnet_tvar_20[0][51] , 
	\_zy_simnet_tvar_20[0][50] , \_zy_simnet_tvar_20[0][49] , 
	\_zy_simnet_tvar_20[0][48] , \_zy_simnet_tvar_20[0][47] , 
	\_zy_simnet_tvar_20[0][46] , \_zy_simnet_tvar_20[0][45] , 
	\_zy_simnet_tvar_20[0][44] , \_zy_simnet_tvar_20[0][43] , 
	\_zy_simnet_tvar_20[0][42] , \_zy_simnet_tvar_20[0][41] , 
	\_zy_simnet_tvar_20[0][40] , \_zy_simnet_tvar_20[0][39] , 
	\_zy_simnet_tvar_20[0][38] , \_zy_simnet_tvar_20[0][37] , 
	\_zy_simnet_tvar_20[0][36] , \_zy_simnet_tvar_20[0][35] , 
	\_zy_simnet_tvar_20[0][34] , \_zy_simnet_tvar_20[0][33] , 
	\_zy_simnet_tvar_20[0][32] , \_zy_simnet_tvar_20[0][31] , 
	\_zy_simnet_tvar_20[0][30] , \_zy_simnet_tvar_20[0][29] , 
	\_zy_simnet_tvar_20[0][28] , \_zy_simnet_tvar_20[0][27] , 
	\_zy_simnet_tvar_20[0][26] , \_zy_simnet_tvar_20[0][25] , 
	\_zy_simnet_tvar_20[0][24] , \_zy_simnet_tvar_20[0][23] , 
	\_zy_simnet_tvar_20[0][22] , \_zy_simnet_tvar_20[0][21] , 
	\_zy_simnet_tvar_20[0][20] , \_zy_simnet_tvar_20[0][19] , 
	\_zy_simnet_tvar_20[0][18] , \_zy_simnet_tvar_20[0][17] , 
	\_zy_simnet_tvar_20[0][16] , \_zy_simnet_tvar_20[0][15] , 
	\_zy_simnet_tvar_20[0][14] , \_zy_simnet_tvar_20[0][13] , 
	\_zy_simnet_tvar_20[0][12] , \_zy_simnet_tvar_20[0][11] , 
	\_zy_simnet_tvar_20[0][10] , \_zy_simnet_tvar_20[0][9] , 
	\_zy_simnet_tvar_20[0][8] , \_zy_simnet_tvar_20[0][7] , 
	\_zy_simnet_tvar_20[0][6] , \_zy_simnet_tvar_20[0][5] , 
	\_zy_simnet_tvar_20[0][4] , \_zy_simnet_tvar_20[0][3] , 
	\_zy_simnet_tvar_20[0][2] , \_zy_simnet_tvar_20[0][1] , 
	\_zy_simnet_tvar_20[0][0] }), .seed0_valid( seed0_valid), 
	.seed0_internal_state_key( seed0_internal_state_key[255:0]), 
	.seed0_internal_state_value( seed0_internal_state_value[127:0]), 
	.seed0_reseed_interval( seed0_reseed_interval[47:0]), 
	.seed1_valid( seed1_valid), .seed1_internal_state_key( 
	seed1_internal_state_key[255:0]), .seed1_internal_state_value( 
	seed1_internal_state_value[127:0]), .seed1_reseed_interval( 
	seed1_reseed_interval[47:0]), .tready_override( 
	_zy_simnet_tready_override_21_w$[0:8]), 
	.cceip_encrypt_kop_fifo_override( 
	_zy_simnet_cceip_encrypt_kop_fifo_override_22_w$[0:6]), 
	.cceip_validate_kop_fifo_override( 
	_zy_simnet_cceip_validate_kop_fifo_override_23_w$[0:6]), 
	.cddip_decrypt_kop_fifo_override( 
	_zy_simnet_cddip_decrypt_kop_fifo_override_24_w$[0:6]), 
	.kdf_test_key_size( kdf_test_key_size[31:0]), .kdf_test_mode_en( 
	kdf_test_mode_en), .sa_global_ctrl( 
	_zy_simnet_sa_global_ctrl_25_w$[0:31]), .sa_ctrl( { \sa_ctrl[31][31] , 
	\sa_ctrl[31][30] , \sa_ctrl[31][29] , \sa_ctrl[31][28] , 
	\sa_ctrl[31][27] , \sa_ctrl[31][26] , \sa_ctrl[31][25] , 
	\sa_ctrl[31][24] , \sa_ctrl[31][23] , \sa_ctrl[31][22] , 
	\sa_ctrl[31][21] , \sa_ctrl[31][20] , \sa_ctrl[31][19] , 
	\sa_ctrl[31][18] , \sa_ctrl[31][17] , \sa_ctrl[31][16] , 
	\sa_ctrl[31][15] , \sa_ctrl[31][14] , \sa_ctrl[31][13] , 
	\sa_ctrl[31][12] , \sa_ctrl[31][11] , \sa_ctrl[31][10] , 
	\sa_ctrl[31][9] , \sa_ctrl[31][8] , \sa_ctrl[31][7] , 
	\sa_ctrl[31][6] , \sa_ctrl[31][5] , \sa_ctrl[31][4] , 
	\sa_ctrl[31][3] , \sa_ctrl[31][2] , \sa_ctrl[31][1] , 
	\sa_ctrl[31][0] , \sa_ctrl[30][31] , \sa_ctrl[30][30] , 
	\sa_ctrl[30][29] , \sa_ctrl[30][28] , \sa_ctrl[30][27] , 
	\sa_ctrl[30][26] , \sa_ctrl[30][25] , \sa_ctrl[30][24] , 
	\sa_ctrl[30][23] , \sa_ctrl[30][22] , \sa_ctrl[30][21] , 
	\sa_ctrl[30][20] , \sa_ctrl[30][19] , \sa_ctrl[30][18] , 
	\sa_ctrl[30][17] , \sa_ctrl[30][16] , \sa_ctrl[30][15] , 
	\sa_ctrl[30][14] , \sa_ctrl[30][13] , \sa_ctrl[30][12] , 
	\sa_ctrl[30][11] , \sa_ctrl[30][10] , \sa_ctrl[30][9] , 
	\sa_ctrl[30][8] , \sa_ctrl[30][7] , \sa_ctrl[30][6] , 
	\sa_ctrl[30][5] , \sa_ctrl[30][4] , \sa_ctrl[30][3] , 
	\sa_ctrl[30][2] , \sa_ctrl[30][1] , \sa_ctrl[30][0] , 
	\sa_ctrl[29][31] , \sa_ctrl[29][30] , \sa_ctrl[29][29] , 
	\sa_ctrl[29][28] , \sa_ctrl[29][27] , \sa_ctrl[29][26] , 
	\sa_ctrl[29][25] , \sa_ctrl[29][24] , \sa_ctrl[29][23] , 
	\sa_ctrl[29][22] , \sa_ctrl[29][21] , \sa_ctrl[29][20] , 
	\sa_ctrl[29][19] , \sa_ctrl[29][18] , \sa_ctrl[29][17] , 
	\sa_ctrl[29][16] , \sa_ctrl[29][15] , \sa_ctrl[29][14] , 
	\sa_ctrl[29][13] , \sa_ctrl[29][12] , \sa_ctrl[29][11] , 
	\sa_ctrl[29][10] , \sa_ctrl[29][9] , \sa_ctrl[29][8] , 
	\sa_ctrl[29][7] , \sa_ctrl[29][6] , \sa_ctrl[29][5] , 
	\sa_ctrl[29][4] , \sa_ctrl[29][3] , \sa_ctrl[29][2] , 
	\sa_ctrl[29][1] , \sa_ctrl[29][0] , \sa_ctrl[28][31] , 
	\sa_ctrl[28][30] , \sa_ctrl[28][29] , \sa_ctrl[28][28] , 
	\sa_ctrl[28][27] , \sa_ctrl[28][26] , \sa_ctrl[28][25] , 
	\sa_ctrl[28][24] , \sa_ctrl[28][23] , \sa_ctrl[28][22] , 
	\sa_ctrl[28][21] , \sa_ctrl[28][20] , \sa_ctrl[28][19] , 
	\sa_ctrl[28][18] , \sa_ctrl[28][17] , \sa_ctrl[28][16] , 
	\sa_ctrl[28][15] , \sa_ctrl[28][14] , \sa_ctrl[28][13] , 
	\sa_ctrl[28][12] , \sa_ctrl[28][11] , \sa_ctrl[28][10] , 
	\sa_ctrl[28][9] , \sa_ctrl[28][8] , \sa_ctrl[28][7] , 
	\sa_ctrl[28][6] , \sa_ctrl[28][5] , \sa_ctrl[28][4] , 
	\sa_ctrl[28][3] , \sa_ctrl[28][2] , \sa_ctrl[28][1] , 
	\sa_ctrl[28][0] , \sa_ctrl[27][31] , \sa_ctrl[27][30] , 
	\sa_ctrl[27][29] , \sa_ctrl[27][28] , \sa_ctrl[27][27] , 
	\sa_ctrl[27][26] , \sa_ctrl[27][25] , \sa_ctrl[27][24] , 
	\sa_ctrl[27][23] , \sa_ctrl[27][22] , \sa_ctrl[27][21] , 
	\sa_ctrl[27][20] , \sa_ctrl[27][19] , \sa_ctrl[27][18] , 
	\sa_ctrl[27][17] , \sa_ctrl[27][16] , \sa_ctrl[27][15] , 
	\sa_ctrl[27][14] , \sa_ctrl[27][13] , \sa_ctrl[27][12] , 
	\sa_ctrl[27][11] , \sa_ctrl[27][10] , \sa_ctrl[27][9] , 
	\sa_ctrl[27][8] , \sa_ctrl[27][7] , \sa_ctrl[27][6] , 
	\sa_ctrl[27][5] , \sa_ctrl[27][4] , \sa_ctrl[27][3] , 
	\sa_ctrl[27][2] , \sa_ctrl[27][1] , \sa_ctrl[27][0] , 
	\sa_ctrl[26][31] , \sa_ctrl[26][30] , \sa_ctrl[26][29] , 
	\sa_ctrl[26][28] , \sa_ctrl[26][27] , \sa_ctrl[26][26] , 
	\sa_ctrl[26][25] , \sa_ctrl[26][24] , \sa_ctrl[26][23] , 
	\sa_ctrl[26][22] , \sa_ctrl[26][21] , \sa_ctrl[26][20] , 
	\sa_ctrl[26][19] , \sa_ctrl[26][18] , \sa_ctrl[26][17] , 
	\sa_ctrl[26][16] , \sa_ctrl[26][15] , \sa_ctrl[26][14] , 
	\sa_ctrl[26][13] , \sa_ctrl[26][12] , \sa_ctrl[26][11] , 
	\sa_ctrl[26][10] , \sa_ctrl[26][9] , \sa_ctrl[26][8] , 
	\sa_ctrl[26][7] , \sa_ctrl[26][6] , \sa_ctrl[26][5] , 
	\sa_ctrl[26][4] , \sa_ctrl[26][3] , \sa_ctrl[26][2] , 
	\sa_ctrl[26][1] , \sa_ctrl[26][0] , \sa_ctrl[25][31] , 
	\sa_ctrl[25][30] , \sa_ctrl[25][29] , \sa_ctrl[25][28] , 
	\sa_ctrl[25][27] , \sa_ctrl[25][26] , \sa_ctrl[25][25] , 
	\sa_ctrl[25][24] , \sa_ctrl[25][23] , \sa_ctrl[25][22] , 
	\sa_ctrl[25][21] , \sa_ctrl[25][20] , \sa_ctrl[25][19] , 
	\sa_ctrl[25][18] , \sa_ctrl[25][17] , \sa_ctrl[25][16] , 
	\sa_ctrl[25][15] , \sa_ctrl[25][14] , \sa_ctrl[25][13] , 
	\sa_ctrl[25][12] , \sa_ctrl[25][11] , \sa_ctrl[25][10] , 
	\sa_ctrl[25][9] , \sa_ctrl[25][8] , \sa_ctrl[25][7] , 
	\sa_ctrl[25][6] , \sa_ctrl[25][5] , \sa_ctrl[25][4] , 
	\sa_ctrl[25][3] , \sa_ctrl[25][2] , \sa_ctrl[25][1] , 
	\sa_ctrl[25][0] , \sa_ctrl[24][31] , \sa_ctrl[24][30] , 
	\sa_ctrl[24][29] , \sa_ctrl[24][28] , \sa_ctrl[24][27] , 
	\sa_ctrl[24][26] , \sa_ctrl[24][25] , \sa_ctrl[24][24] , 
	\sa_ctrl[24][23] , \sa_ctrl[24][22] , \sa_ctrl[24][21] , 
	\sa_ctrl[24][20] , \sa_ctrl[24][19] , \sa_ctrl[24][18] , 
	\sa_ctrl[24][17] , \sa_ctrl[24][16] , \sa_ctrl[24][15] , 
	\sa_ctrl[24][14] , \sa_ctrl[24][13] , \sa_ctrl[24][12] , 
	\sa_ctrl[24][11] , \sa_ctrl[24][10] , \sa_ctrl[24][9] , 
	\sa_ctrl[24][8] , \sa_ctrl[24][7] , \sa_ctrl[24][6] , 
	\sa_ctrl[24][5] , \sa_ctrl[24][4] , \sa_ctrl[24][3] , 
	\sa_ctrl[24][2] , \sa_ctrl[24][1] , \sa_ctrl[24][0] , 
	\sa_ctrl[23][31] , \sa_ctrl[23][30] , \sa_ctrl[23][29] , 
	\sa_ctrl[23][28] , \sa_ctrl[23][27] , \sa_ctrl[23][26] , 
	\sa_ctrl[23][25] , \sa_ctrl[23][24] , \sa_ctrl[23][23] , 
	\sa_ctrl[23][22] , \sa_ctrl[23][21] , \sa_ctrl[23][20] , 
	\sa_ctrl[23][19] , \sa_ctrl[23][18] , \sa_ctrl[23][17] , 
	\sa_ctrl[23][16] , \sa_ctrl[23][15] , \sa_ctrl[23][14] , 
	\sa_ctrl[23][13] , \sa_ctrl[23][12] , \sa_ctrl[23][11] , 
	\sa_ctrl[23][10] , \sa_ctrl[23][9] , \sa_ctrl[23][8] , 
	\sa_ctrl[23][7] , \sa_ctrl[23][6] , \sa_ctrl[23][5] , 
	\sa_ctrl[23][4] , \sa_ctrl[23][3] , \sa_ctrl[23][2] , 
	\sa_ctrl[23][1] , \sa_ctrl[23][0] , \sa_ctrl[22][31] , 
	\sa_ctrl[22][30] , \sa_ctrl[22][29] , \sa_ctrl[22][28] , 
	\sa_ctrl[22][27] , \sa_ctrl[22][26] , \sa_ctrl[22][25] , 
	\sa_ctrl[22][24] , \sa_ctrl[22][23] , \sa_ctrl[22][22] , 
	\sa_ctrl[22][21] , \sa_ctrl[22][20] , \sa_ctrl[22][19] , 
	\sa_ctrl[22][18] , \sa_ctrl[22][17] , \sa_ctrl[22][16] , 
	\sa_ctrl[22][15] , \sa_ctrl[22][14] , \sa_ctrl[22][13] , 
	\sa_ctrl[22][12] , \sa_ctrl[22][11] , \sa_ctrl[22][10] , 
	\sa_ctrl[22][9] , \sa_ctrl[22][8] , \sa_ctrl[22][7] , 
	\sa_ctrl[22][6] , \sa_ctrl[22][5] , \sa_ctrl[22][4] , 
	\sa_ctrl[22][3] , \sa_ctrl[22][2] , \sa_ctrl[22][1] , 
	\sa_ctrl[22][0] , \sa_ctrl[21][31] , \sa_ctrl[21][30] , 
	\sa_ctrl[21][29] , \sa_ctrl[21][28] , \sa_ctrl[21][27] , 
	\sa_ctrl[21][26] , \sa_ctrl[21][25] , \sa_ctrl[21][24] , 
	\sa_ctrl[21][23] , \sa_ctrl[21][22] , \sa_ctrl[21][21] , 
	\sa_ctrl[21][20] , \sa_ctrl[21][19] , \sa_ctrl[21][18] , 
	\sa_ctrl[21][17] , \sa_ctrl[21][16] , \sa_ctrl[21][15] , 
	\sa_ctrl[21][14] , \sa_ctrl[21][13] , \sa_ctrl[21][12] , 
	\sa_ctrl[21][11] , \sa_ctrl[21][10] , \sa_ctrl[21][9] , 
	\sa_ctrl[21][8] , \sa_ctrl[21][7] , \sa_ctrl[21][6] , 
	\sa_ctrl[21][5] , \sa_ctrl[21][4] , \sa_ctrl[21][3] , 
	\sa_ctrl[21][2] , \sa_ctrl[21][1] , \sa_ctrl[21][0] , 
	\sa_ctrl[20][31] , \sa_ctrl[20][30] , \sa_ctrl[20][29] , 
	\sa_ctrl[20][28] , \sa_ctrl[20][27] , \sa_ctrl[20][26] , 
	\sa_ctrl[20][25] , \sa_ctrl[20][24] , \sa_ctrl[20][23] , 
	\sa_ctrl[20][22] , \sa_ctrl[20][21] , \sa_ctrl[20][20] , 
	\sa_ctrl[20][19] , \sa_ctrl[20][18] , \sa_ctrl[20][17] , 
	\sa_ctrl[20][16] , \sa_ctrl[20][15] , \sa_ctrl[20][14] , 
	\sa_ctrl[20][13] , \sa_ctrl[20][12] , \sa_ctrl[20][11] , 
	\sa_ctrl[20][10] , \sa_ctrl[20][9] , \sa_ctrl[20][8] , 
	\sa_ctrl[20][7] , \sa_ctrl[20][6] , \sa_ctrl[20][5] , 
	\sa_ctrl[20][4] , \sa_ctrl[20][3] , \sa_ctrl[20][2] , 
	\sa_ctrl[20][1] , \sa_ctrl[20][0] , \sa_ctrl[19][31] , 
	\sa_ctrl[19][30] , \sa_ctrl[19][29] , \sa_ctrl[19][28] , 
	\sa_ctrl[19][27] , \sa_ctrl[19][26] , \sa_ctrl[19][25] , 
	\sa_ctrl[19][24] , \sa_ctrl[19][23] , \sa_ctrl[19][22] , 
	\sa_ctrl[19][21] , \sa_ctrl[19][20] , \sa_ctrl[19][19] , 
	\sa_ctrl[19][18] , \sa_ctrl[19][17] , \sa_ctrl[19][16] , 
	\sa_ctrl[19][15] , \sa_ctrl[19][14] , \sa_ctrl[19][13] , 
	\sa_ctrl[19][12] , \sa_ctrl[19][11] , \sa_ctrl[19][10] , 
	\sa_ctrl[19][9] , \sa_ctrl[19][8] , \sa_ctrl[19][7] , 
	\sa_ctrl[19][6] , \sa_ctrl[19][5] , \sa_ctrl[19][4] , 
	\sa_ctrl[19][3] , \sa_ctrl[19][2] , \sa_ctrl[19][1] , 
	\sa_ctrl[19][0] , \sa_ctrl[18][31] , \sa_ctrl[18][30] , 
	\sa_ctrl[18][29] , \sa_ctrl[18][28] , \sa_ctrl[18][27] , 
	\sa_ctrl[18][26] , \sa_ctrl[18][25] , \sa_ctrl[18][24] , 
	\sa_ctrl[18][23] , \sa_ctrl[18][22] , \sa_ctrl[18][21] , 
	\sa_ctrl[18][20] , \sa_ctrl[18][19] , \sa_ctrl[18][18] , 
	\sa_ctrl[18][17] , \sa_ctrl[18][16] , \sa_ctrl[18][15] , 
	\sa_ctrl[18][14] , \sa_ctrl[18][13] , \sa_ctrl[18][12] , 
	\sa_ctrl[18][11] , \sa_ctrl[18][10] , \sa_ctrl[18][9] , 
	\sa_ctrl[18][8] , \sa_ctrl[18][7] , \sa_ctrl[18][6] , 
	\sa_ctrl[18][5] , \sa_ctrl[18][4] , \sa_ctrl[18][3] , 
	\sa_ctrl[18][2] , \sa_ctrl[18][1] , \sa_ctrl[18][0] , 
	\sa_ctrl[17][31] , \sa_ctrl[17][30] , \sa_ctrl[17][29] , 
	\sa_ctrl[17][28] , \sa_ctrl[17][27] , \sa_ctrl[17][26] , 
	\sa_ctrl[17][25] , \sa_ctrl[17][24] , \sa_ctrl[17][23] , 
	\sa_ctrl[17][22] , \sa_ctrl[17][21] , \sa_ctrl[17][20] , 
	\sa_ctrl[17][19] , \sa_ctrl[17][18] , \sa_ctrl[17][17] , 
	\sa_ctrl[17][16] , \sa_ctrl[17][15] , \sa_ctrl[17][14] , 
	\sa_ctrl[17][13] , \sa_ctrl[17][12] , \sa_ctrl[17][11] , 
	\sa_ctrl[17][10] , \sa_ctrl[17][9] , \sa_ctrl[17][8] , 
	\sa_ctrl[17][7] , \sa_ctrl[17][6] , \sa_ctrl[17][5] , 
	\sa_ctrl[17][4] , \sa_ctrl[17][3] , \sa_ctrl[17][2] , 
	\sa_ctrl[17][1] , \sa_ctrl[17][0] , \sa_ctrl[16][31] , 
	\sa_ctrl[16][30] , \sa_ctrl[16][29] , \sa_ctrl[16][28] , 
	\sa_ctrl[16][27] , \sa_ctrl[16][26] , \sa_ctrl[16][25] , 
	\sa_ctrl[16][24] , \sa_ctrl[16][23] , \sa_ctrl[16][22] , 
	\sa_ctrl[16][21] , \sa_ctrl[16][20] , \sa_ctrl[16][19] , 
	\sa_ctrl[16][18] , \sa_ctrl[16][17] , \sa_ctrl[16][16] , 
	\sa_ctrl[16][15] , \sa_ctrl[16][14] , \sa_ctrl[16][13] , 
	\sa_ctrl[16][12] , \sa_ctrl[16][11] , \sa_ctrl[16][10] , 
	\sa_ctrl[16][9] , \sa_ctrl[16][8] , \sa_ctrl[16][7] , 
	\sa_ctrl[16][6] , \sa_ctrl[16][5] , \sa_ctrl[16][4] , 
	\sa_ctrl[16][3] , \sa_ctrl[16][2] , \sa_ctrl[16][1] , 
	\sa_ctrl[16][0] , \sa_ctrl[15][31] , \sa_ctrl[15][30] , 
	\sa_ctrl[15][29] , \sa_ctrl[15][28] , \sa_ctrl[15][27] , 
	\sa_ctrl[15][26] , \sa_ctrl[15][25] , \sa_ctrl[15][24] , 
	\sa_ctrl[15][23] , \sa_ctrl[15][22] , \sa_ctrl[15][21] , 
	\sa_ctrl[15][20] , \sa_ctrl[15][19] , \sa_ctrl[15][18] , 
	\sa_ctrl[15][17] , \sa_ctrl[15][16] , \sa_ctrl[15][15] , 
	\sa_ctrl[15][14] , \sa_ctrl[15][13] , \sa_ctrl[15][12] , 
	\sa_ctrl[15][11] , \sa_ctrl[15][10] , \sa_ctrl[15][9] , 
	\sa_ctrl[15][8] , \sa_ctrl[15][7] , \sa_ctrl[15][6] , 
	\sa_ctrl[15][5] , \sa_ctrl[15][4] , \sa_ctrl[15][3] , 
	\sa_ctrl[15][2] , \sa_ctrl[15][1] , \sa_ctrl[15][0] , 
	\sa_ctrl[14][31] , \sa_ctrl[14][30] , \sa_ctrl[14][29] , 
	\sa_ctrl[14][28] , \sa_ctrl[14][27] , \sa_ctrl[14][26] , 
	\sa_ctrl[14][25] , \sa_ctrl[14][24] , \sa_ctrl[14][23] , 
	\sa_ctrl[14][22] , \sa_ctrl[14][21] , \sa_ctrl[14][20] , 
	\sa_ctrl[14][19] , \sa_ctrl[14][18] , \sa_ctrl[14][17] , 
	\sa_ctrl[14][16] , \sa_ctrl[14][15] , \sa_ctrl[14][14] , 
	\sa_ctrl[14][13] , \sa_ctrl[14][12] , \sa_ctrl[14][11] , 
	\sa_ctrl[14][10] , \sa_ctrl[14][9] , \sa_ctrl[14][8] , 
	\sa_ctrl[14][7] , \sa_ctrl[14][6] , \sa_ctrl[14][5] , 
	\sa_ctrl[14][4] , \sa_ctrl[14][3] , \sa_ctrl[14][2] , 
	\sa_ctrl[14][1] , \sa_ctrl[14][0] , \sa_ctrl[13][31] , 
	\sa_ctrl[13][30] , \sa_ctrl[13][29] , \sa_ctrl[13][28] , 
	\sa_ctrl[13][27] , \sa_ctrl[13][26] , \sa_ctrl[13][25] , 
	\sa_ctrl[13][24] , \sa_ctrl[13][23] , \sa_ctrl[13][22] , 
	\sa_ctrl[13][21] , \sa_ctrl[13][20] , \sa_ctrl[13][19] , 
	\sa_ctrl[13][18] , \sa_ctrl[13][17] , \sa_ctrl[13][16] , 
	\sa_ctrl[13][15] , \sa_ctrl[13][14] , \sa_ctrl[13][13] , 
	\sa_ctrl[13][12] , \sa_ctrl[13][11] , \sa_ctrl[13][10] , 
	\sa_ctrl[13][9] , \sa_ctrl[13][8] , \sa_ctrl[13][7] , 
	\sa_ctrl[13][6] , \sa_ctrl[13][5] , \sa_ctrl[13][4] , 
	\sa_ctrl[13][3] , \sa_ctrl[13][2] , \sa_ctrl[13][1] , 
	\sa_ctrl[13][0] , \sa_ctrl[12][31] , \sa_ctrl[12][30] , 
	\sa_ctrl[12][29] , \sa_ctrl[12][28] , \sa_ctrl[12][27] , 
	\sa_ctrl[12][26] , \sa_ctrl[12][25] , \sa_ctrl[12][24] , 
	\sa_ctrl[12][23] , \sa_ctrl[12][22] , \sa_ctrl[12][21] , 
	\sa_ctrl[12][20] , \sa_ctrl[12][19] , \sa_ctrl[12][18] , 
	\sa_ctrl[12][17] , \sa_ctrl[12][16] , \sa_ctrl[12][15] , 
	\sa_ctrl[12][14] , \sa_ctrl[12][13] , \sa_ctrl[12][12] , 
	\sa_ctrl[12][11] , \sa_ctrl[12][10] , \sa_ctrl[12][9] , 
	\sa_ctrl[12][8] , \sa_ctrl[12][7] , \sa_ctrl[12][6] , 
	\sa_ctrl[12][5] , \sa_ctrl[12][4] , \sa_ctrl[12][3] , 
	\sa_ctrl[12][2] , \sa_ctrl[12][1] , \sa_ctrl[12][0] , 
	\sa_ctrl[11][31] , \sa_ctrl[11][30] , \sa_ctrl[11][29] , 
	\sa_ctrl[11][28] , \sa_ctrl[11][27] , \sa_ctrl[11][26] , 
	\sa_ctrl[11][25] , \sa_ctrl[11][24] , \sa_ctrl[11][23] , 
	\sa_ctrl[11][22] , \sa_ctrl[11][21] , \sa_ctrl[11][20] , 
	\sa_ctrl[11][19] , \sa_ctrl[11][18] , \sa_ctrl[11][17] , 
	\sa_ctrl[11][16] , \sa_ctrl[11][15] , \sa_ctrl[11][14] , 
	\sa_ctrl[11][13] , \sa_ctrl[11][12] , \sa_ctrl[11][11] , 
	\sa_ctrl[11][10] , \sa_ctrl[11][9] , \sa_ctrl[11][8] , 
	\sa_ctrl[11][7] , \sa_ctrl[11][6] , \sa_ctrl[11][5] , 
	\sa_ctrl[11][4] , \sa_ctrl[11][3] , \sa_ctrl[11][2] , 
	\sa_ctrl[11][1] , \sa_ctrl[11][0] , \sa_ctrl[10][31] , 
	\sa_ctrl[10][30] , \sa_ctrl[10][29] , \sa_ctrl[10][28] , 
	\sa_ctrl[10][27] , \sa_ctrl[10][26] , \sa_ctrl[10][25] , 
	\sa_ctrl[10][24] , \sa_ctrl[10][23] , \sa_ctrl[10][22] , 
	\sa_ctrl[10][21] , \sa_ctrl[10][20] , \sa_ctrl[10][19] , 
	\sa_ctrl[10][18] , \sa_ctrl[10][17] , \sa_ctrl[10][16] , 
	\sa_ctrl[10][15] , \sa_ctrl[10][14] , \sa_ctrl[10][13] , 
	\sa_ctrl[10][12] , \sa_ctrl[10][11] , \sa_ctrl[10][10] , 
	\sa_ctrl[10][9] , \sa_ctrl[10][8] , \sa_ctrl[10][7] , 
	\sa_ctrl[10][6] , \sa_ctrl[10][5] , \sa_ctrl[10][4] , 
	\sa_ctrl[10][3] , \sa_ctrl[10][2] , \sa_ctrl[10][1] , 
	\sa_ctrl[10][0] , \sa_ctrl[9][31] , \sa_ctrl[9][30] , 
	\sa_ctrl[9][29] , \sa_ctrl[9][28] , \sa_ctrl[9][27] , 
	\sa_ctrl[9][26] , \sa_ctrl[9][25] , \sa_ctrl[9][24] , 
	\sa_ctrl[9][23] , \sa_ctrl[9][22] , \sa_ctrl[9][21] , 
	\sa_ctrl[9][20] , \sa_ctrl[9][19] , \sa_ctrl[9][18] , 
	\sa_ctrl[9][17] , \sa_ctrl[9][16] , \sa_ctrl[9][15] , 
	\sa_ctrl[9][14] , \sa_ctrl[9][13] , \sa_ctrl[9][12] , 
	\sa_ctrl[9][11] , \sa_ctrl[9][10] , \sa_ctrl[9][9] , \sa_ctrl[9][8] , 
	\sa_ctrl[9][7] , \sa_ctrl[9][6] , \sa_ctrl[9][5] , \sa_ctrl[9][4] , 
	\sa_ctrl[9][3] , \sa_ctrl[9][2] , \sa_ctrl[9][1] , \sa_ctrl[9][0] , 
	\sa_ctrl[8][31] , \sa_ctrl[8][30] , \sa_ctrl[8][29] , 
	\sa_ctrl[8][28] , \sa_ctrl[8][27] , \sa_ctrl[8][26] , 
	\sa_ctrl[8][25] , \sa_ctrl[8][24] , \sa_ctrl[8][23] , 
	\sa_ctrl[8][22] , \sa_ctrl[8][21] , \sa_ctrl[8][20] , 
	\sa_ctrl[8][19] , \sa_ctrl[8][18] , \sa_ctrl[8][17] , 
	\sa_ctrl[8][16] , \sa_ctrl[8][15] , \sa_ctrl[8][14] , 
	\sa_ctrl[8][13] , \sa_ctrl[8][12] , \sa_ctrl[8][11] , 
	\sa_ctrl[8][10] , \sa_ctrl[8][9] , \sa_ctrl[8][8] , \sa_ctrl[8][7] , 
	\sa_ctrl[8][6] , \sa_ctrl[8][5] , \sa_ctrl[8][4] , \sa_ctrl[8][3] , 
	\sa_ctrl[8][2] , \sa_ctrl[8][1] , \sa_ctrl[8][0] , \sa_ctrl[7][31] , 
	\sa_ctrl[7][30] , \sa_ctrl[7][29] , \sa_ctrl[7][28] , 
	\sa_ctrl[7][27] , \sa_ctrl[7][26] , \sa_ctrl[7][25] , 
	\sa_ctrl[7][24] , \sa_ctrl[7][23] , \sa_ctrl[7][22] , 
	\sa_ctrl[7][21] , \sa_ctrl[7][20] , \sa_ctrl[7][19] , 
	\sa_ctrl[7][18] , \sa_ctrl[7][17] , \sa_ctrl[7][16] , 
	\sa_ctrl[7][15] , \sa_ctrl[7][14] , \sa_ctrl[7][13] , 
	\sa_ctrl[7][12] , \sa_ctrl[7][11] , \sa_ctrl[7][10] , 
	\sa_ctrl[7][9] , \sa_ctrl[7][8] , \sa_ctrl[7][7] , \sa_ctrl[7][6] , 
	\sa_ctrl[7][5] , \sa_ctrl[7][4] , \sa_ctrl[7][3] , \sa_ctrl[7][2] , 
	\sa_ctrl[7][1] , \sa_ctrl[7][0] , \sa_ctrl[6][31] , \sa_ctrl[6][30] , 
	\sa_ctrl[6][29] , \sa_ctrl[6][28] , \sa_ctrl[6][27] , 
	\sa_ctrl[6][26] , \sa_ctrl[6][25] , \sa_ctrl[6][24] , 
	\sa_ctrl[6][23] , \sa_ctrl[6][22] , \sa_ctrl[6][21] , 
	\sa_ctrl[6][20] , \sa_ctrl[6][19] , \sa_ctrl[6][18] , 
	\sa_ctrl[6][17] , \sa_ctrl[6][16] , \sa_ctrl[6][15] , 
	\sa_ctrl[6][14] , \sa_ctrl[6][13] , \sa_ctrl[6][12] , 
	\sa_ctrl[6][11] , \sa_ctrl[6][10] , \sa_ctrl[6][9] , \sa_ctrl[6][8] , 
	\sa_ctrl[6][7] , \sa_ctrl[6][6] , \sa_ctrl[6][5] , \sa_ctrl[6][4] , 
	\sa_ctrl[6][3] , \sa_ctrl[6][2] , \sa_ctrl[6][1] , \sa_ctrl[6][0] , 
	\sa_ctrl[5][31] , \sa_ctrl[5][30] , \sa_ctrl[5][29] , 
	\sa_ctrl[5][28] , \sa_ctrl[5][27] , \sa_ctrl[5][26] , 
	\sa_ctrl[5][25] , \sa_ctrl[5][24] , \sa_ctrl[5][23] , 
	\sa_ctrl[5][22] , \sa_ctrl[5][21] , \sa_ctrl[5][20] , 
	\sa_ctrl[5][19] , \sa_ctrl[5][18] , \sa_ctrl[5][17] , 
	\sa_ctrl[5][16] , \sa_ctrl[5][15] , \sa_ctrl[5][14] , 
	\sa_ctrl[5][13] , \sa_ctrl[5][12] , \sa_ctrl[5][11] , 
	\sa_ctrl[5][10] , \sa_ctrl[5][9] , \sa_ctrl[5][8] , \sa_ctrl[5][7] , 
	\sa_ctrl[5][6] , \sa_ctrl[5][5] , \sa_ctrl[5][4] , \sa_ctrl[5][3] , 
	\sa_ctrl[5][2] , \sa_ctrl[5][1] , \sa_ctrl[5][0] , \sa_ctrl[4][31] , 
	\sa_ctrl[4][30] , \sa_ctrl[4][29] , \sa_ctrl[4][28] , 
	\sa_ctrl[4][27] , \sa_ctrl[4][26] , \sa_ctrl[4][25] , 
	\sa_ctrl[4][24] , \sa_ctrl[4][23] , \sa_ctrl[4][22] , 
	\sa_ctrl[4][21] , \sa_ctrl[4][20] , \sa_ctrl[4][19] , 
	\sa_ctrl[4][18] , \sa_ctrl[4][17] , \sa_ctrl[4][16] , 
	\sa_ctrl[4][15] , \sa_ctrl[4][14] , \sa_ctrl[4][13] , 
	\sa_ctrl[4][12] , \sa_ctrl[4][11] , \sa_ctrl[4][10] , 
	\sa_ctrl[4][9] , \sa_ctrl[4][8] , \sa_ctrl[4][7] , \sa_ctrl[4][6] , 
	\sa_ctrl[4][5] , \sa_ctrl[4][4] , \sa_ctrl[4][3] , \sa_ctrl[4][2] , 
	\sa_ctrl[4][1] , \sa_ctrl[4][0] , \sa_ctrl[3][31] , \sa_ctrl[3][30] , 
	\sa_ctrl[3][29] , \sa_ctrl[3][28] , \sa_ctrl[3][27] , 
	\sa_ctrl[3][26] , \sa_ctrl[3][25] , \sa_ctrl[3][24] , 
	\sa_ctrl[3][23] , \sa_ctrl[3][22] , \sa_ctrl[3][21] , 
	\sa_ctrl[3][20] , \sa_ctrl[3][19] , \sa_ctrl[3][18] , 
	\sa_ctrl[3][17] , \sa_ctrl[3][16] , \sa_ctrl[3][15] , 
	\sa_ctrl[3][14] , \sa_ctrl[3][13] , \sa_ctrl[3][12] , 
	\sa_ctrl[3][11] , \sa_ctrl[3][10] , \sa_ctrl[3][9] , \sa_ctrl[3][8] , 
	\sa_ctrl[3][7] , \sa_ctrl[3][6] , \sa_ctrl[3][5] , \sa_ctrl[3][4] , 
	\sa_ctrl[3][3] , \sa_ctrl[3][2] , \sa_ctrl[3][1] , \sa_ctrl[3][0] , 
	\sa_ctrl[2][31] , \sa_ctrl[2][30] , \sa_ctrl[2][29] , 
	\sa_ctrl[2][28] , \sa_ctrl[2][27] , \sa_ctrl[2][26] , 
	\sa_ctrl[2][25] , \sa_ctrl[2][24] , \sa_ctrl[2][23] , 
	\sa_ctrl[2][22] , \sa_ctrl[2][21] , \sa_ctrl[2][20] , 
	\sa_ctrl[2][19] , \sa_ctrl[2][18] , \sa_ctrl[2][17] , 
	\sa_ctrl[2][16] , \sa_ctrl[2][15] , \sa_ctrl[2][14] , 
	\sa_ctrl[2][13] , \sa_ctrl[2][12] , \sa_ctrl[2][11] , 
	\sa_ctrl[2][10] , \sa_ctrl[2][9] , \sa_ctrl[2][8] , \sa_ctrl[2][7] , 
	\sa_ctrl[2][6] , \sa_ctrl[2][5] , \sa_ctrl[2][4] , \sa_ctrl[2][3] , 
	\sa_ctrl[2][2] , \sa_ctrl[2][1] , \sa_ctrl[2][0] , \sa_ctrl[1][31] , 
	\sa_ctrl[1][30] , \sa_ctrl[1][29] , \sa_ctrl[1][28] , 
	\sa_ctrl[1][27] , \sa_ctrl[1][26] , \sa_ctrl[1][25] , 
	\sa_ctrl[1][24] , \sa_ctrl[1][23] , \sa_ctrl[1][22] , 
	\sa_ctrl[1][21] , \sa_ctrl[1][20] , \sa_ctrl[1][19] , 
	\sa_ctrl[1][18] , \sa_ctrl[1][17] , \sa_ctrl[1][16] , 
	\sa_ctrl[1][15] , \sa_ctrl[1][14] , \sa_ctrl[1][13] , 
	\sa_ctrl[1][12] , \sa_ctrl[1][11] , \sa_ctrl[1][10] , 
	\sa_ctrl[1][9] , \sa_ctrl[1][8] , \sa_ctrl[1][7] , \sa_ctrl[1][6] , 
	\sa_ctrl[1][5] , \sa_ctrl[1][4] , \sa_ctrl[1][3] , \sa_ctrl[1][2] , 
	\sa_ctrl[1][1] , \sa_ctrl[1][0] , \sa_ctrl[0][31] , \sa_ctrl[0][30] , 
	\sa_ctrl[0][29] , \sa_ctrl[0][28] , \sa_ctrl[0][27] , 
	\sa_ctrl[0][26] , \sa_ctrl[0][25] , \sa_ctrl[0][24] , 
	\sa_ctrl[0][23] , \sa_ctrl[0][22] , \sa_ctrl[0][21] , 
	\sa_ctrl[0][20] , \sa_ctrl[0][19] , \sa_ctrl[0][18] , 
	\sa_ctrl[0][17] , \sa_ctrl[0][16] , \sa_ctrl[0][15] , 
	\sa_ctrl[0][14] , \sa_ctrl[0][13] , \sa_ctrl[0][12] , 
	\sa_ctrl[0][11] , \sa_ctrl[0][10] , \sa_ctrl[0][9] , \sa_ctrl[0][8] , 
	\sa_ctrl[0][7] , \sa_ctrl[0][6] , \sa_ctrl[0][5] , \sa_ctrl[0][4] , 
	\sa_ctrl[0][3] , \sa_ctrl[0][2] , \sa_ctrl[0][1] , \sa_ctrl[0][0] }));
cr_rst_sync cr_rst_sync ( .clk( clk), .async_rst_n( rst_n), .bypass_reset( 
	scan_mode), .test_rst_n( scan_rst_n), .rst_n( rst_sync_n));
ixc_expEv _zyclock_1_x$tbcp ( _zyclock_1_x$tbc, clock_1);
ixc_assign_32 _zz_strnp_85 ( _zy_simnet_idle_components_78_w$[0:31], 
	idle_components[31:0]);
ixc_assign _zz_strnp_84 ( _zy_simnet_kme_cddip3_ob_in_77_w$, 
	kme_cddip3_ob_in[0]);
ixc_assign_83 _zz_strnp_83 ( _zy_simnet_kme_cddip3_ob_out_pre_76_w$[0:82], 
	kme_cddip3_ob_out_pre[82:0]);
ixc_assign _zz_strnp_82 ( _zy_simnet_kme_cddip2_ob_in_75_w$, 
	kme_cddip2_ob_in[0]);
ixc_assign_83 _zz_strnp_81 ( _zy_simnet_kme_cddip2_ob_out_pre_74_w$[0:82], 
	kme_cddip2_ob_out_pre[82:0]);
ixc_assign _zz_strnp_80 ( _zy_simnet_kme_cddip1_ob_in_73_w$, 
	kme_cddip1_ob_in[0]);
ixc_assign_83 _zz_strnp_79 ( _zy_simnet_kme_cddip1_ob_out_pre_72_w$[0:82], 
	kme_cddip1_ob_out_pre[82:0]);
ixc_assign _zz_strnp_78 ( _zy_simnet_kme_cddip0_ob_in_71_w$, 
	kme_cddip0_ob_in[0]);
ixc_assign_83 _zz_strnp_77 ( _zy_simnet_kme_cddip0_ob_out_pre_70_w$[0:82], 
	kme_cddip0_ob_out_pre[82:0]);
ixc_assign _zz_strnp_76 ( _zy_simnet_kme_cceip3_ob_in_69_w$, 
	kme_cceip3_ob_in[0]);
ixc_assign_83 _zz_strnp_75 ( _zy_simnet_kme_cceip3_ob_out_pre_68_w$[0:82], 
	kme_cceip3_ob_out_pre[82:0]);
ixc_assign _zz_strnp_74 ( _zy_simnet_kme_cceip2_ob_in_67_w$, 
	kme_cceip2_ob_in[0]);
ixc_assign_83 _zz_strnp_73 ( _zy_simnet_kme_cceip2_ob_out_pre_66_w$[0:82], 
	kme_cceip2_ob_out_pre[82:0]);
ixc_assign _zz_strnp_72 ( _zy_simnet_kme_cceip1_ob_in_65_w$, 
	kme_cceip1_ob_in[0]);
ixc_assign_83 _zz_strnp_71 ( _zy_simnet_kme_cceip1_ob_out_pre_64_w$[0:82], 
	kme_cceip1_ob_out_pre[82:0]);
ixc_assign _zz_strnp_70 ( _zy_simnet_kme_cceip0_ob_in_63_w$, 
	kme_cceip0_ob_in[0]);
ixc_assign_83 _zz_strnp_69 ( _zy_simnet_kme_cceip0_ob_out_pre_62_w$[0:82], 
	kme_cceip0_ob_out_pre[82:0]);
ixc_assign_84 _zz_strnp_68 ( _zy_simnet_rbus_ring_i_59_w$[0:83], 
	rbus_ring_i[83:0]);
ixc_assign_32 _zz_strnp_67 ( sa_global_ctrl[31:0], 
	_zy_simnet_sa_global_ctrl_58_w$[0:31]);
ixc_assign_7 _zz_strnp_66 ( cddip_decrypt_kop_fifo_override[6:0], 
	_zy_simnet_cddip_decrypt_kop_fifo_override_57_w$[0:6]);
ixc_assign_7 _zz_strnp_65 ( cceip_validate_kop_fifo_override[6:0], 
	_zy_simnet_cceip_validate_kop_fifo_override_56_w$[0:6]);
ixc_assign_7 _zz_strnp_64 ( cceip_encrypt_kop_fifo_override[6:0], 
	_zy_simnet_cceip_encrypt_kop_fifo_override_55_w$[0:6]);
ixc_assign_9 _zz_strnp_63 ( tready_override[8:0], 
	_zy_simnet_tready_override_54_w$[0:8]);
ixc_assign_38 _zz_strnp_61 ( kim_dout[37:0], _zy_simnet_kim_dout_52_w$[0:37]);
ixc_assign _zz_strnp_60 ( kme_cddip3_ob_in_mod[0], 
	_zy_simnet_kme_cddip3_ob_in_mod_51_w$);
ixc_assign_83 _zz_strnp_59 ( kme_cddip3_ob_out[82:0], 
	_zy_simnet_kme_cddip3_ob_out_50_w$[0:82]);
ixc_assign _zz_strnp_58 ( kme_cddip2_ob_in_mod[0], 
	_zy_simnet_kme_cddip2_ob_in_mod_49_w$);
ixc_assign_83 _zz_strnp_57 ( kme_cddip2_ob_out[82:0], 
	_zy_simnet_kme_cddip2_ob_out_48_w$[0:82]);
ixc_assign _zz_strnp_56 ( kme_cddip1_ob_in_mod[0], 
	_zy_simnet_kme_cddip1_ob_in_mod_47_w$);
ixc_assign_83 _zz_strnp_55 ( kme_cddip1_ob_out[82:0], 
	_zy_simnet_kme_cddip1_ob_out_46_w$[0:82]);
ixc_assign _zz_strnp_54 ( kme_cddip0_ob_in_mod[0], 
	_zy_simnet_kme_cddip0_ob_in_mod_45_w$);
ixc_assign_83 _zz_strnp_53 ( kme_cddip0_ob_out[82:0], 
	_zy_simnet_kme_cddip0_ob_out_44_w$[0:82]);
ixc_assign _zz_strnp_52 ( kme_cceip3_ob_in_mod[0], 
	_zy_simnet_kme_cceip3_ob_in_mod_43_w$);
ixc_assign_83 _zz_strnp_51 ( kme_cceip3_ob_out[82:0], 
	_zy_simnet_kme_cceip3_ob_out_42_w$[0:82]);
ixc_assign _zz_strnp_50 ( kme_cceip2_ob_in_mod[0], 
	_zy_simnet_kme_cceip2_ob_in_mod_41_w$);
ixc_assign_83 _zz_strnp_49 ( kme_cceip2_ob_out[82:0], 
	_zy_simnet_kme_cceip2_ob_out_40_w$[0:82]);
ixc_assign _zz_strnp_48 ( kme_cceip1_ob_in_mod[0], 
	_zy_simnet_kme_cceip1_ob_in_mod_39_w$);
ixc_assign_83 _zz_strnp_47 ( kme_cceip1_ob_out[82:0], 
	_zy_simnet_kme_cceip1_ob_out_38_w$[0:82]);
ixc_assign _zz_strnp_46 ( kme_cceip0_ob_in_mod[0], 
	_zy_simnet_kme_cceip0_ob_in_mod_37_w$);
ixc_assign_83 _zz_strnp_45 ( kme_cceip0_ob_out[82:0], 
	_zy_simnet_kme_cceip0_ob_out_36_w$[0:82]);
ixc_assign_84 _zz_strnp_44 ( rbus_ring_o[83:0], 
	_zy_simnet_rbus_ring_o_35_w$[0:83]);
ixc_assign _zz_strnp_43 ( _zy_simnet_rbus_ring_o_34_w$, rbus_ring_o[34]);
ixc_assign _zz_strnp_42 ( _zy_simnet_rbus_ring_o_33_w$, rbus_ring_o[67]);
ixc_assign _zz_strnp_41 ( _zy_simnet_rbus_ring_o_32_w$, rbus_ring_o[0]);
ixc_assign _zz_strnp_40 ( _zy_simnet_rbus_ring_o_31_w$, rbus_ring_o[1]);
ixc_assign_32 _zz_strnp_39 ( _zy_simnet_rbus_ring_o_30_w$[0:31], 
	rbus_ring_o[33:2]);
ixc_assign _zz_strnp_38 ( rbus_ring_i[34], _zy_simnet_rbus_ring_i_29_w$);
ixc_assign_32 _zz_strnp_37 ( rbus_ring_i[66:35], 
	_zy_simnet_rbus_ring_i_28_w$[0:31]);
ixc_assign _zz_strnp_36 ( rbus_ring_i[67], _zy_simnet_rbus_ring_i_27_w$);
ixc_assign_16 _zz_strnp_35 ( rbus_ring_i[83:68], 
	_zy_simnet_rbus_ring_i_26_w$[0:15]);
ixc_assign_32 _zz_strnp_34 ( _zy_simnet_sa_global_ctrl_25_w$[0:31], 
	sa_global_ctrl[31:0]);
ixc_assign_7 _zz_strnp_33 ( 
	_zy_simnet_cddip_decrypt_kop_fifo_override_24_w$[0:6], 
	cddip_decrypt_kop_fifo_override[6:0]);
ixc_assign_7 _zz_strnp_32 ( 
	_zy_simnet_cceip_validate_kop_fifo_override_23_w$[0:6], 
	cceip_validate_kop_fifo_override[6:0]);
ixc_assign_7 _zz_strnp_31 ( 
	_zy_simnet_cceip_encrypt_kop_fifo_override_22_w$[0:6], 
	cceip_encrypt_kop_fifo_override[6:0]);
ixc_assign_9 _zz_strnp_30 ( _zy_simnet_tready_override_21_w$[0:8], 
	tready_override[8:0]);
ixc_assign_38 _zz_strnp_28 ( _zy_simnet_kim_dout_19_w$[0:37], kim_dout[37:0]);
ixc_assign _zz_strnp_27 ( _zy_simnet_kme_cddip3_ob_in_mod_18_w$, 
	kme_cddip3_ob_in_mod[0]);
ixc_assign _zz_strnp_26 ( _zy_simnet_kme_cddip2_ob_in_mod_17_w$, 
	kme_cddip2_ob_in_mod[0]);
ixc_assign _zz_strnp_25 ( _zy_simnet_kme_cddip1_ob_in_mod_16_w$, 
	kme_cddip1_ob_in_mod[0]);
ixc_assign _zz_strnp_24 ( _zy_simnet_kme_cddip0_ob_in_mod_15_w$, 
	kme_cddip0_ob_in_mod[0]);
ixc_assign _zz_strnp_23 ( _zy_simnet_kme_cceip3_ob_in_mod_14_w$, 
	kme_cceip3_ob_in_mod[0]);
ixc_assign _zz_strnp_22 ( _zy_simnet_kme_cceip2_ob_in_mod_13_w$, 
	kme_cceip2_ob_in_mod[0]);
ixc_assign _zz_strnp_21 ( _zy_simnet_kme_cceip1_ob_in_mod_12_w$, 
	kme_cceip1_ob_in_mod[0]);
ixc_assign _zz_strnp_20 ( _zy_simnet_kme_cceip0_ob_in_mod_11_w$, 
	kme_cceip0_ob_in_mod[0]);
ixc_assign_83 _zz_strnp_19 ( _zy_simnet_kme_ib_in_10_w$[0:82], 
	kme_ib_in[82:0]);
ixc_assign_32 _zz_strnp_18 ( idle_components[31:0], 
	_zy_simnet_idle_components_9_w$[0:31]);
ixc_assign_83 _zz_strnp_17 ( kme_cddip3_ob_out_pre[82:0], 
	_zy_simnet_kme_cddip3_ob_out_pre_8_w$[0:82]);
ixc_assign_83 _zz_strnp_16 ( kme_cddip2_ob_out_pre[82:0], 
	_zy_simnet_kme_cddip2_ob_out_pre_7_w$[0:82]);
ixc_assign_83 _zz_strnp_15 ( kme_cddip1_ob_out_pre[82:0], 
	_zy_simnet_kme_cddip1_ob_out_pre_6_w$[0:82]);
ixc_assign_83 _zz_strnp_14 ( kme_cddip0_ob_out_pre[82:0], 
	_zy_simnet_kme_cddip0_ob_out_pre_5_w$[0:82]);
ixc_assign_83 _zz_strnp_13 ( kme_cceip3_ob_out_pre[82:0], 
	_zy_simnet_kme_cceip3_ob_out_pre_4_w$[0:82]);
ixc_assign_83 _zz_strnp_12 ( kme_cceip2_ob_out_pre[82:0], 
	_zy_simnet_kme_cceip2_ob_out_pre_3_w$[0:82]);
ixc_assign_83 _zz_strnp_11 ( kme_cceip1_ob_out_pre[82:0], 
	_zy_simnet_kme_cceip1_ob_out_pre_2_w$[0:82]);
ixc_assign_83 _zz_strnp_10 ( kme_cceip0_ob_out_pre[82:0], 
	_zy_simnet_kme_cceip0_ob_out_pre_1_w$[0:82]);
ixc_assign _zz_strnp_9 ( kme_ib_out[0], _zy_simnet_kme_ib_out_0_w$);
ixc_assign _zz_strnp_8 ( kme_cceip0_ob_in[0], kme_cceip0_ob_tready);
ixc_assign_64 _zz_strnp_7 ( kme_cceip0_ob_tdata[63:0], 
	kme_cceip0_ob_out[63:0]);
ixc_assign_8 _zz_strnp_6 ( kme_cceip0_ob_tuser[7:0], kme_cceip0_ob_out[71:64]);
ixc_assign_8 _zz_strnp_5 ( kme_cceip0_ob_tstrb[7:0], kme_cceip0_ob_out[79:72]);
ixc_assign _zz_strnp_4 ( kme_cceip0_ob_tid[0], kme_cceip0_ob_out[80]);
ixc_assign _zz_strnp_3 ( kme_cceip0_ob_tlast, kme_cceip0_ob_out[81]);
ixc_assign _zz_strnp_2 ( kme_cceip0_ob_tvalid, kme_cceip0_ob_out[82]);
ixc_assign _zz_strnp_1 ( clock_1, clock);
ixc_assign _zz_strnp_0 ( clk, clock);
Q_MX02 U164 ( .S(manual_txc), .A0(kme_ib_tvalid), .A1(debug_kme_ib_tvalid), .Z(kme_ib_in[82]));
Q_MX02 U165 ( .S(manual_txc), .A0(kme_ib_tlast), .A1(debug_kme_ib_tlast), .Z(kme_ib_in[81]));
Q_MX02 U166 ( .S(manual_txc), .A0(kme_ib_tid[0]), .A1(debug_kme_ib_tid[0]), .Z(kme_ib_in[80]));
Q_MX02 U167 ( .S(manual_txc), .A0(kme_ib_tstrb[0]), .A1(debug_kme_ib_tstrb[0]), .Z(kme_ib_in[72]));
Q_MX02 U168 ( .S(manual_txc), .A0(kme_ib_tstrb[1]), .A1(debug_kme_ib_tstrb[1]), .Z(kme_ib_in[73]));
Q_MX02 U169 ( .S(manual_txc), .A0(kme_ib_tstrb[2]), .A1(debug_kme_ib_tstrb[2]), .Z(kme_ib_in[74]));
Q_MX02 U170 ( .S(manual_txc), .A0(kme_ib_tstrb[3]), .A1(debug_kme_ib_tstrb[3]), .Z(kme_ib_in[75]));
Q_MX02 U171 ( .S(manual_txc), .A0(kme_ib_tstrb[4]), .A1(debug_kme_ib_tstrb[4]), .Z(kme_ib_in[76]));
Q_MX02 U172 ( .S(manual_txc), .A0(kme_ib_tstrb[5]), .A1(debug_kme_ib_tstrb[5]), .Z(kme_ib_in[77]));
Q_MX02 U173 ( .S(manual_txc), .A0(kme_ib_tstrb[6]), .A1(debug_kme_ib_tstrb[6]), .Z(kme_ib_in[78]));
Q_MX02 U174 ( .S(manual_txc), .A0(kme_ib_tstrb[7]), .A1(debug_kme_ib_tstrb[7]), .Z(kme_ib_in[79]));
Q_MX02 U175 ( .S(manual_txc), .A0(kme_ib_tuser[0]), .A1(debug_kme_ib_tuser[0]), .Z(kme_ib_in[64]));
Q_MX02 U176 ( .S(manual_txc), .A0(kme_ib_tuser[1]), .A1(debug_kme_ib_tuser[1]), .Z(kme_ib_in[65]));
Q_MX02 U177 ( .S(manual_txc), .A0(kme_ib_tuser[2]), .A1(debug_kme_ib_tuser[2]), .Z(kme_ib_in[66]));
Q_MX02 U178 ( .S(manual_txc), .A0(kme_ib_tuser[3]), .A1(debug_kme_ib_tuser[3]), .Z(kme_ib_in[67]));
Q_MX02 U179 ( .S(manual_txc), .A0(kme_ib_tuser[4]), .A1(debug_kme_ib_tuser[4]), .Z(kme_ib_in[68]));
Q_MX02 U180 ( .S(manual_txc), .A0(kme_ib_tuser[5]), .A1(debug_kme_ib_tuser[5]), .Z(kme_ib_in[69]));
Q_MX02 U181 ( .S(manual_txc), .A0(kme_ib_tuser[6]), .A1(debug_kme_ib_tuser[6]), .Z(kme_ib_in[70]));
Q_MX02 U182 ( .S(manual_txc), .A0(kme_ib_tuser[7]), .A1(debug_kme_ib_tuser[7]), .Z(kme_ib_in[71]));
Q_MX02 U183 ( .S(manual_txc), .A0(kme_ib_tdata[0]), .A1(debug_kme_ib_tdata[0]), .Z(kme_ib_in[0]));
Q_MX02 U184 ( .S(manual_txc), .A0(kme_ib_tdata[1]), .A1(debug_kme_ib_tdata[1]), .Z(kme_ib_in[1]));
Q_MX02 U185 ( .S(manual_txc), .A0(kme_ib_tdata[2]), .A1(debug_kme_ib_tdata[2]), .Z(kme_ib_in[2]));
Q_MX02 U186 ( .S(manual_txc), .A0(kme_ib_tdata[3]), .A1(debug_kme_ib_tdata[3]), .Z(kme_ib_in[3]));
Q_MX02 U187 ( .S(manual_txc), .A0(kme_ib_tdata[4]), .A1(debug_kme_ib_tdata[4]), .Z(kme_ib_in[4]));
Q_MX02 U188 ( .S(manual_txc), .A0(kme_ib_tdata[5]), .A1(debug_kme_ib_tdata[5]), .Z(kme_ib_in[5]));
Q_MX02 U189 ( .S(manual_txc), .A0(kme_ib_tdata[6]), .A1(debug_kme_ib_tdata[6]), .Z(kme_ib_in[6]));
Q_MX02 U190 ( .S(manual_txc), .A0(kme_ib_tdata[7]), .A1(debug_kme_ib_tdata[7]), .Z(kme_ib_in[7]));
Q_MX02 U191 ( .S(manual_txc), .A0(kme_ib_tdata[8]), .A1(debug_kme_ib_tdata[8]), .Z(kme_ib_in[8]));
Q_MX02 U192 ( .S(manual_txc), .A0(kme_ib_tdata[9]), .A1(debug_kme_ib_tdata[9]), .Z(kme_ib_in[9]));
Q_MX02 U193 ( .S(manual_txc), .A0(kme_ib_tdata[10]), .A1(debug_kme_ib_tdata[10]), .Z(kme_ib_in[10]));
Q_MX02 U194 ( .S(manual_txc), .A0(kme_ib_tdata[11]), .A1(debug_kme_ib_tdata[11]), .Z(kme_ib_in[11]));
Q_MX02 U195 ( .S(manual_txc), .A0(kme_ib_tdata[12]), .A1(debug_kme_ib_tdata[12]), .Z(kme_ib_in[12]));
Q_MX02 U196 ( .S(manual_txc), .A0(kme_ib_tdata[13]), .A1(debug_kme_ib_tdata[13]), .Z(kme_ib_in[13]));
Q_MX02 U197 ( .S(manual_txc), .A0(kme_ib_tdata[14]), .A1(debug_kme_ib_tdata[14]), .Z(kme_ib_in[14]));
Q_MX02 U198 ( .S(manual_txc), .A0(kme_ib_tdata[15]), .A1(debug_kme_ib_tdata[15]), .Z(kme_ib_in[15]));
Q_MX02 U199 ( .S(manual_txc), .A0(kme_ib_tdata[16]), .A1(debug_kme_ib_tdata[16]), .Z(kme_ib_in[16]));
Q_MX02 U200 ( .S(manual_txc), .A0(kme_ib_tdata[17]), .A1(debug_kme_ib_tdata[17]), .Z(kme_ib_in[17]));
Q_MX02 U201 ( .S(manual_txc), .A0(kme_ib_tdata[18]), .A1(debug_kme_ib_tdata[18]), .Z(kme_ib_in[18]));
Q_MX02 U202 ( .S(manual_txc), .A0(kme_ib_tdata[19]), .A1(debug_kme_ib_tdata[19]), .Z(kme_ib_in[19]));
Q_MX02 U203 ( .S(manual_txc), .A0(kme_ib_tdata[20]), .A1(debug_kme_ib_tdata[20]), .Z(kme_ib_in[20]));
Q_MX02 U204 ( .S(manual_txc), .A0(kme_ib_tdata[21]), .A1(debug_kme_ib_tdata[21]), .Z(kme_ib_in[21]));
Q_MX02 U205 ( .S(manual_txc), .A0(kme_ib_tdata[22]), .A1(debug_kme_ib_tdata[22]), .Z(kme_ib_in[22]));
Q_MX02 U206 ( .S(manual_txc), .A0(kme_ib_tdata[23]), .A1(debug_kme_ib_tdata[23]), .Z(kme_ib_in[23]));
Q_MX02 U207 ( .S(manual_txc), .A0(kme_ib_tdata[24]), .A1(debug_kme_ib_tdata[24]), .Z(kme_ib_in[24]));
Q_MX02 U208 ( .S(manual_txc), .A0(kme_ib_tdata[25]), .A1(debug_kme_ib_tdata[25]), .Z(kme_ib_in[25]));
Q_MX02 U209 ( .S(manual_txc), .A0(kme_ib_tdata[26]), .A1(debug_kme_ib_tdata[26]), .Z(kme_ib_in[26]));
Q_MX02 U210 ( .S(manual_txc), .A0(kme_ib_tdata[27]), .A1(debug_kme_ib_tdata[27]), .Z(kme_ib_in[27]));
Q_MX02 U211 ( .S(manual_txc), .A0(kme_ib_tdata[28]), .A1(debug_kme_ib_tdata[28]), .Z(kme_ib_in[28]));
Q_MX02 U212 ( .S(manual_txc), .A0(kme_ib_tdata[29]), .A1(debug_kme_ib_tdata[29]), .Z(kme_ib_in[29]));
Q_MX02 U213 ( .S(manual_txc), .A0(kme_ib_tdata[30]), .A1(debug_kme_ib_tdata[30]), .Z(kme_ib_in[30]));
Q_MX02 U214 ( .S(manual_txc), .A0(kme_ib_tdata[31]), .A1(debug_kme_ib_tdata[31]), .Z(kme_ib_in[31]));
Q_MX02 U215 ( .S(manual_txc), .A0(kme_ib_tdata[32]), .A1(debug_kme_ib_tdata[32]), .Z(kme_ib_in[32]));
Q_MX02 U216 ( .S(manual_txc), .A0(kme_ib_tdata[33]), .A1(debug_kme_ib_tdata[33]), .Z(kme_ib_in[33]));
Q_MX02 U217 ( .S(manual_txc), .A0(kme_ib_tdata[34]), .A1(debug_kme_ib_tdata[34]), .Z(kme_ib_in[34]));
Q_MX02 U218 ( .S(manual_txc), .A0(kme_ib_tdata[35]), .A1(debug_kme_ib_tdata[35]), .Z(kme_ib_in[35]));
Q_MX02 U219 ( .S(manual_txc), .A0(kme_ib_tdata[36]), .A1(debug_kme_ib_tdata[36]), .Z(kme_ib_in[36]));
Q_MX02 U220 ( .S(manual_txc), .A0(kme_ib_tdata[37]), .A1(debug_kme_ib_tdata[37]), .Z(kme_ib_in[37]));
Q_MX02 U221 ( .S(manual_txc), .A0(kme_ib_tdata[38]), .A1(debug_kme_ib_tdata[38]), .Z(kme_ib_in[38]));
Q_MX02 U222 ( .S(manual_txc), .A0(kme_ib_tdata[39]), .A1(debug_kme_ib_tdata[39]), .Z(kme_ib_in[39]));
Q_MX02 U223 ( .S(manual_txc), .A0(kme_ib_tdata[40]), .A1(debug_kme_ib_tdata[40]), .Z(kme_ib_in[40]));
Q_MX02 U224 ( .S(manual_txc), .A0(kme_ib_tdata[41]), .A1(debug_kme_ib_tdata[41]), .Z(kme_ib_in[41]));
Q_MX02 U225 ( .S(manual_txc), .A0(kme_ib_tdata[42]), .A1(debug_kme_ib_tdata[42]), .Z(kme_ib_in[42]));
Q_MX02 U226 ( .S(manual_txc), .A0(kme_ib_tdata[43]), .A1(debug_kme_ib_tdata[43]), .Z(kme_ib_in[43]));
Q_MX02 U227 ( .S(manual_txc), .A0(kme_ib_tdata[44]), .A1(debug_kme_ib_tdata[44]), .Z(kme_ib_in[44]));
Q_MX02 U228 ( .S(manual_txc), .A0(kme_ib_tdata[45]), .A1(debug_kme_ib_tdata[45]), .Z(kme_ib_in[45]));
Q_MX02 U229 ( .S(manual_txc), .A0(kme_ib_tdata[46]), .A1(debug_kme_ib_tdata[46]), .Z(kme_ib_in[46]));
Q_MX02 U230 ( .S(manual_txc), .A0(kme_ib_tdata[47]), .A1(debug_kme_ib_tdata[47]), .Z(kme_ib_in[47]));
Q_MX02 U231 ( .S(manual_txc), .A0(kme_ib_tdata[48]), .A1(debug_kme_ib_tdata[48]), .Z(kme_ib_in[48]));
Q_MX02 U232 ( .S(manual_txc), .A0(kme_ib_tdata[49]), .A1(debug_kme_ib_tdata[49]), .Z(kme_ib_in[49]));
Q_MX02 U233 ( .S(manual_txc), .A0(kme_ib_tdata[50]), .A1(debug_kme_ib_tdata[50]), .Z(kme_ib_in[50]));
Q_MX02 U234 ( .S(manual_txc), .A0(kme_ib_tdata[51]), .A1(debug_kme_ib_tdata[51]), .Z(kme_ib_in[51]));
Q_MX02 U235 ( .S(manual_txc), .A0(kme_ib_tdata[52]), .A1(debug_kme_ib_tdata[52]), .Z(kme_ib_in[52]));
Q_MX02 U236 ( .S(manual_txc), .A0(kme_ib_tdata[53]), .A1(debug_kme_ib_tdata[53]), .Z(kme_ib_in[53]));
Q_MX02 U237 ( .S(manual_txc), .A0(kme_ib_tdata[54]), .A1(debug_kme_ib_tdata[54]), .Z(kme_ib_in[54]));
Q_MX02 U238 ( .S(manual_txc), .A0(kme_ib_tdata[55]), .A1(debug_kme_ib_tdata[55]), .Z(kme_ib_in[55]));
Q_MX02 U239 ( .S(manual_txc), .A0(kme_ib_tdata[56]), .A1(debug_kme_ib_tdata[56]), .Z(kme_ib_in[56]));
Q_MX02 U240 ( .S(manual_txc), .A0(kme_ib_tdata[57]), .A1(debug_kme_ib_tdata[57]), .Z(kme_ib_in[57]));
Q_MX02 U241 ( .S(manual_txc), .A0(kme_ib_tdata[58]), .A1(debug_kme_ib_tdata[58]), .Z(kme_ib_in[58]));
Q_MX02 U242 ( .S(manual_txc), .A0(kme_ib_tdata[59]), .A1(debug_kme_ib_tdata[59]), .Z(kme_ib_in[59]));
Q_MX02 U243 ( .S(manual_txc), .A0(kme_ib_tdata[60]), .A1(debug_kme_ib_tdata[60]), .Z(kme_ib_in[60]));
Q_MX02 U244 ( .S(manual_txc), .A0(kme_ib_tdata[61]), .A1(debug_kme_ib_tdata[61]), .Z(kme_ib_in[61]));
Q_MX02 U245 ( .S(manual_txc), .A0(kme_ib_tdata[62]), .A1(debug_kme_ib_tdata[62]), .Z(kme_ib_in[62]));
Q_MX02 U246 ( .S(manual_txc), .A0(kme_ib_tdata[63]), .A1(debug_kme_ib_tdata[63]), .Z(kme_ib_in[63]));
Q_OR02 U247 ( .A0(manual_txc), .A1(kme_ib_out[0]), .Z(kme_ib_tready));
Q_INV U248 ( .A(manual_txc), .Z(n3));
Q_OR02 U249 ( .A0(n3), .A1(kme_ib_out[0]), .Z(debug_kme_ib_tready));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "_zy_simnet_tvar_20 (2,0) 1 271 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m2 "_zy_simnet_tvar_53 (2,0) 1 271 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m3 "labels (2,0) 1 271 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m4 "sa_count 1 63 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m5 "sa_ctrl 1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m6 "sa_snapshot 1 63 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "6"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\_zy_simnet_tvar_20%s.guid_size  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\_zy_simnet_tvar_20%s.label_size  1 5 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\_zy_simnet_tvar_20%s.label  1 255 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\_zy_simnet_tvar_20%s.delimiter_valid  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\_zy_simnet_tvar_20%s.delimiter  1 7 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\_zy_simnet_tvar_53%s.guid_size  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\_zy_simnet_tvar_53%s.label_size  1 5 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\_zy_simnet_tvar_53%s.label  1 255 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\_zy_simnet_tvar_53%s.delimiter_valid  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\_zy_simnet_tvar_53%s.delimiter  1 7 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\rbus_ring_i.addr  (1,0) 1 15 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\rbus_ring_i.wr_data  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\rbus_ring_i.rd_data  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\rbus_ring_o.addr  (1,0) 1 15 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\rbus_ring_o.wr_data  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\rbus_ring_o.rd_data  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\kme_ib_in.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\kme_ib_in.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\kme_ib_in.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\kme_ib_in.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\kme_cceip0_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\kme_cceip0_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\kme_cceip0_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\kme_cceip0_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\kme_cceip1_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\kme_cceip1_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\kme_cceip1_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\kme_cceip1_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\kme_cceip2_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\kme_cceip2_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\kme_cceip2_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\kme_cceip2_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\kme_cceip3_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\kme_cceip3_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\kme_cceip3_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\kme_cceip3_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\kme_cddip0_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\kme_cddip0_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m39 "\kme_cddip0_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m40 "\kme_cddip0_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m41 "\kme_cddip1_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m42 "\kme_cddip1_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m43 "\kme_cddip1_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m44 "\kme_cddip1_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m45 "\kme_cddip2_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m46 "\kme_cddip2_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m47 "\kme_cddip2_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m48 "\kme_cddip2_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m49 "\kme_cddip3_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m50 "\kme_cddip3_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m51 "\kme_cddip3_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m52 "\kme_cddip3_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m53 "\cceip_encrypt_kop_fifo_override.r.part0  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m54 "\cceip_validate_kop_fifo_override.r.part0  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m55 "\cddip_decrypt_kop_fifo_override.r.part0  (1,0) 1 6 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m56 "\idle_components.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m57 "\idle_components.f.num_key_tlvs_in_flight  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m58 "\kim_dout.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m59 "\kim_dout.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m60 "\kim_dout.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m61 "\kim_dout.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m62 "\kim_dout.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m63 "\kim_dout.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m64 "\kim_dout.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m65 "\kme_cceip0_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m66 "\kme_cceip0_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m67 "\kme_cceip0_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m68 "\kme_cceip0_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m69 "\kme_cceip1_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m70 "\kme_cceip1_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m71 "\kme_cceip1_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m72 "\kme_cceip1_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m73 "\kme_cceip2_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m74 "\kme_cceip2_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m75 "\kme_cceip2_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m76 "\kme_cceip2_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m77 "\kme_cceip3_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m78 "\kme_cceip3_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m79 "\kme_cceip3_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m80 "\kme_cceip3_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m81 "\kme_cddip0_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m82 "\kme_cddip0_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m83 "\kme_cddip0_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m84 "\kme_cddip0_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m85 "\kme_cddip1_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m86 "\kme_cddip1_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m87 "\kme_cddip1_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m88 "\kme_cddip1_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m89 "\kme_cddip2_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m90 "\kme_cddip2_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m91 "\kme_cddip2_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m92 "\kme_cddip2_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m93 "\kme_cddip3_ob_out_pre.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m94 "\kme_cddip3_ob_out_pre.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m95 "\kme_cddip3_ob_out_pre.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m96 "\kme_cddip3_ob_out_pre.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m97 "\labels%s.guid_size  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m98 "\labels%s.label_size  1 5 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m99 "\labels%s.label  1 255 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m100 "\labels%s.delimiter_valid  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m101 "\labels%s.delimiter  1 7 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m102 "\sa_count%s.r.part1  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m103 "\sa_count%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m104 "\sa_count%s.f.unused  1 13 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m105 "\sa_count%s.f.upper  1 17 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m106 "\sa_count%s.f.lower  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m107 "\sa_ctrl%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m108 "\sa_ctrl%s.f.spare  1 26 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m109 "\sa_ctrl%s.f.sa_event_sel  1 4 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m110 "\sa_global_ctrl.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m111 "\sa_global_ctrl.f.spare  (1,0) 1 29 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m112 "\sa_snapshot%s.r.part1  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m113 "\sa_snapshot%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m114 "\sa_snapshot%s.f.unused  1 13 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m115 "\sa_snapshot%s.f.upper  1 17 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m116 "\sa_snapshot%s.f.lower  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m117 "\tready_override.r.part0  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "117"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "_zy_simnet_tvar_20%s 5 \_zy_simnet_tvar_20%s.guid_size  \_zy_simnet_tvar_20%s.label_size  \_zy_simnet_tvar_20%s.label  \_zy_simnet_tvar_20%s.delimiter_valid  \_zy_simnet_tvar_20%s.delimiter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "_zy_simnet_tvar_53%s 5 \_zy_simnet_tvar_53%s.guid_size  \_zy_simnet_tvar_53%s.label_size  \_zy_simnet_tvar_53%s.label  \_zy_simnet_tvar_53%s.delimiter_valid  \_zy_simnet_tvar_53%s.delimiter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "rbus_ring_i 7 \rbus_ring_i.addr  \rbus_ring_i.wr_strb  \rbus_ring_i.wr_data  \rbus_ring_i.rd_strb  \rbus_ring_i.rd_data  \rbus_ring_i.ack  \rbus_ring_i.err_ack "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "rbus_ring_o 7 \rbus_ring_o.addr  \rbus_ring_o.wr_strb  \rbus_ring_o.wr_data  \rbus_ring_o.rd_strb  \rbus_ring_o.rd_data  \rbus_ring_o.ack  \rbus_ring_o.err_ack "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "kme_ib_in 6 \kme_ib_in.tvalid  \kme_ib_in.tlast  \kme_ib_in.tid  \kme_ib_in.tstrb  \kme_ib_in.tuser  \kme_ib_in.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "kme_ib_out 1 \kme_ib_out.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "kme_cceip0_ob_out 6 \kme_cceip0_ob_out.tvalid  \kme_cceip0_ob_out.tlast  \kme_cceip0_ob_out.tid  \kme_cceip0_ob_out.tstrb  \kme_cceip0_ob_out.tuser  \kme_cceip0_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r8 "kme_cceip1_ob_out 6 \kme_cceip1_ob_out.tvalid  \kme_cceip1_ob_out.tlast  \kme_cceip1_ob_out.tid  \kme_cceip1_ob_out.tstrb  \kme_cceip1_ob_out.tuser  \kme_cceip1_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r9 "kme_cceip2_ob_out 6 \kme_cceip2_ob_out.tvalid  \kme_cceip2_ob_out.tlast  \kme_cceip2_ob_out.tid  \kme_cceip2_ob_out.tstrb  \kme_cceip2_ob_out.tuser  \kme_cceip2_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r10 "kme_cceip3_ob_out 6 \kme_cceip3_ob_out.tvalid  \kme_cceip3_ob_out.tlast  \kme_cceip3_ob_out.tid  \kme_cceip3_ob_out.tstrb  \kme_cceip3_ob_out.tuser  \kme_cceip3_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r11 "kme_cceip0_ob_in 1 \kme_cceip0_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r12 "kme_cceip1_ob_in 1 \kme_cceip1_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r13 "kme_cceip2_ob_in 1 \kme_cceip2_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r14 "kme_cceip3_ob_in 1 \kme_cceip3_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r15 "kme_cddip0_ob_out 6 \kme_cddip0_ob_out.tvalid  \kme_cddip0_ob_out.tlast  \kme_cddip0_ob_out.tid  \kme_cddip0_ob_out.tstrb  \kme_cddip0_ob_out.tuser  \kme_cddip0_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r16 "kme_cddip1_ob_out 6 \kme_cddip1_ob_out.tvalid  \kme_cddip1_ob_out.tlast  \kme_cddip1_ob_out.tid  \kme_cddip1_ob_out.tstrb  \kme_cddip1_ob_out.tuser  \kme_cddip1_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r17 "kme_cddip2_ob_out 6 \kme_cddip2_ob_out.tvalid  \kme_cddip2_ob_out.tlast  \kme_cddip2_ob_out.tid  \kme_cddip2_ob_out.tstrb  \kme_cddip2_ob_out.tuser  \kme_cddip2_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r18 "kme_cddip3_ob_out 6 \kme_cddip3_ob_out.tvalid  \kme_cddip3_ob_out.tlast  \kme_cddip3_ob_out.tid  \kme_cddip3_ob_out.tstrb  \kme_cddip3_ob_out.tuser  \kme_cddip3_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r19 "kme_cddip0_ob_in 1 \kme_cddip0_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r20 "kme_cddip1_ob_in 1 \kme_cddip1_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r21 "kme_cddip2_ob_in 1 \kme_cddip2_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r22 "kme_cddip3_ob_in 1 \kme_cddip3_ob_in.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r1 "cceip_encrypt_kop_fifo_override 2 \cceip_encrypt_kop_fifo_override.r  { \cceip_encrypt_kop_fifo_override.r.part0  } \cceip_encrypt_kop_fifo_override.f  { \cceip_encrypt_kop_fifo_override.f.gcm_status_data_fifo  \cceip_encrypt_kop_fifo_override.f.tlv_sb_data_fifo  \cceip_encrypt_kop_fifo_override.f.kdf_cmd_fifo  \cceip_encrypt_kop_fifo_override.f.kdfstream_cmd_fifo  \cceip_encrypt_kop_fifo_override.f.keyfilter_cmd_fifo  \cceip_encrypt_kop_fifo_override.f.gcm_tag_data_fifo  \cceip_encrypt_kop_fifo_override.f.gcm_cmd_fifo  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r2 "cceip_validate_kop_fifo_override 2 \cceip_validate_kop_fifo_override.r  { \cceip_validate_kop_fifo_override.r.part0  } \cceip_validate_kop_fifo_override.f  { \cceip_validate_kop_fifo_override.f.gcm_status_data_fifo  \cceip_validate_kop_fifo_override.f.tlv_sb_data_fifo  \cceip_validate_kop_fifo_override.f.kdf_cmd_fifo  \cceip_validate_kop_fifo_override.f.kdfstream_cmd_fifo  \cceip_validate_kop_fifo_override.f.keyfilter_cmd_fifo  \cceip_validate_kop_fifo_override.f.gcm_tag_data_fifo  \cceip_validate_kop_fifo_override.f.gcm_cmd_fifo  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r3 "cddip_decrypt_kop_fifo_override 2 \cddip_decrypt_kop_fifo_override.r  { \cddip_decrypt_kop_fifo_override.r.part0  } \cddip_decrypt_kop_fifo_override.f  { \cddip_decrypt_kop_fifo_override.f.gcm_status_data_fifo  \cddip_decrypt_kop_fifo_override.f.tlv_sb_data_fifo  \cddip_decrypt_kop_fifo_override.f.kdf_cmd_fifo  \cddip_decrypt_kop_fifo_override.f.kdfstream_cmd_fifo  \cddip_decrypt_kop_fifo_override.f.keyfilter_cmd_fifo  \cddip_decrypt_kop_fifo_override.f.gcm_tag_data_fifo  \cddip_decrypt_kop_fifo_override.f.gcm_cmd_fifo  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r4 "idle_components 2 \idle_components.r  { \idle_components.r.part0  } \idle_components.f  { \idle_components.f.num_key_tlvs_in_flight  \idle_components.f.cddip0_key_tlv_rsm_idle  \idle_components.f.cddip1_key_tlv_rsm_idle  \idle_components.f.cddip2_key_tlv_rsm_idle  \idle_components.f.cddip3_key_tlv_rsm_idle  \idle_components.f.cceip0_key_tlv_rsm_idle  \idle_components.f.cceip1_key_tlv_rsm_idle  \idle_components.f.cceip2_key_tlv_rsm_idle  \idle_components.f.cceip3_key_tlv_rsm_idle  \idle_components.f.no_key_tlv_in_flight  \idle_components.f.tlv_parser_idle  \idle_components.f.drng_idle  \idle_components.f.kme_slv_empty  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r23 "kim_dout 7 \kim_dout.valid  \kim_dout.label_index  \kim_dout.ckv_length  \kim_dout.ckv_pointer  \kim_dout.pf_num  \kim_dout.vf_num  \kim_dout.vf_valid "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r24 "kme_cceip0_ob_in_mod 1 \kme_cceip0_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r25 "kme_cceip0_ob_out_pre 6 \kme_cceip0_ob_out_pre.tvalid  \kme_cceip0_ob_out_pre.tlast  \kme_cceip0_ob_out_pre.tid  \kme_cceip0_ob_out_pre.tstrb  \kme_cceip0_ob_out_pre.tuser  \kme_cceip0_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r26 "kme_cceip1_ob_in_mod 1 \kme_cceip1_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r27 "kme_cceip1_ob_out_pre 6 \kme_cceip1_ob_out_pre.tvalid  \kme_cceip1_ob_out_pre.tlast  \kme_cceip1_ob_out_pre.tid  \kme_cceip1_ob_out_pre.tstrb  \kme_cceip1_ob_out_pre.tuser  \kme_cceip1_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r28 "kme_cceip2_ob_in_mod 1 \kme_cceip2_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r29 "kme_cceip2_ob_out_pre 6 \kme_cceip2_ob_out_pre.tvalid  \kme_cceip2_ob_out_pre.tlast  \kme_cceip2_ob_out_pre.tid  \kme_cceip2_ob_out_pre.tstrb  \kme_cceip2_ob_out_pre.tuser  \kme_cceip2_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r30 "kme_cceip3_ob_in_mod 1 \kme_cceip3_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r31 "kme_cceip3_ob_out_pre 6 \kme_cceip3_ob_out_pre.tvalid  \kme_cceip3_ob_out_pre.tlast  \kme_cceip3_ob_out_pre.tid  \kme_cceip3_ob_out_pre.tstrb  \kme_cceip3_ob_out_pre.tuser  \kme_cceip3_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r32 "kme_cddip0_ob_in_mod 1 \kme_cddip0_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r33 "kme_cddip0_ob_out_pre 6 \kme_cddip0_ob_out_pre.tvalid  \kme_cddip0_ob_out_pre.tlast  \kme_cddip0_ob_out_pre.tid  \kme_cddip0_ob_out_pre.tstrb  \kme_cddip0_ob_out_pre.tuser  \kme_cddip0_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r34 "kme_cddip1_ob_in_mod 1 \kme_cddip1_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r35 "kme_cddip1_ob_out_pre 6 \kme_cddip1_ob_out_pre.tvalid  \kme_cddip1_ob_out_pre.tlast  \kme_cddip1_ob_out_pre.tid  \kme_cddip1_ob_out_pre.tstrb  \kme_cddip1_ob_out_pre.tuser  \kme_cddip1_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r36 "kme_cddip2_ob_in_mod 1 \kme_cddip2_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r37 "kme_cddip2_ob_out_pre 6 \kme_cddip2_ob_out_pre.tvalid  \kme_cddip2_ob_out_pre.tlast  \kme_cddip2_ob_out_pre.tid  \kme_cddip2_ob_out_pre.tstrb  \kme_cddip2_ob_out_pre.tuser  \kme_cddip2_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r38 "kme_cddip3_ob_in_mod 1 \kme_cddip3_ob_in_mod.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r39 "kme_cddip3_ob_out_pre 6 \kme_cddip3_ob_out_pre.tvalid  \kme_cddip3_ob_out_pre.tlast  \kme_cddip3_ob_out_pre.tid  \kme_cddip3_ob_out_pre.tstrb  \kme_cddip3_ob_out_pre.tuser  \kme_cddip3_ob_out_pre.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r40 "labels%s 5 \labels%s.guid_size  \labels%s.label_size  \labels%s.label  \labels%s.delimiter_valid  \labels%s.delimiter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r5 "sa_count%s 2 \sa_count%s.r  { \sa_count%s.r.part1  \sa_count%s.r.part0  } \sa_count%s.f  { \sa_count%s.f.unused  \sa_count%s.f.upper  \sa_count%s.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r6 "sa_ctrl%s 2 \sa_ctrl%s.r  { \sa_ctrl%s.r.part0  } \sa_ctrl%s.f  { \sa_ctrl%s.f.spare  \sa_ctrl%s.f.sa_event_sel  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r7 "sa_global_ctrl 2 \sa_global_ctrl.r  { \sa_global_ctrl.r.part0  } \sa_global_ctrl.f  { \sa_global_ctrl.f.spare  \sa_global_ctrl.f.sa_snap  \sa_global_ctrl.f.sa_clear_live  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r8 "sa_snapshot%s 2 \sa_snapshot%s.r  { \sa_snapshot%s.r.part1  \sa_snapshot%s.r.part0  } \sa_snapshot%s.f  { \sa_snapshot%s.f.unused  \sa_snapshot%s.f.upper  \sa_snapshot%s.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r9 "tready_override 2 \tready_override.r  { \tready_override.r.part0  } \tready_override.f  { \tready_override.f.txc_tready_override  \tready_override.f.engine_7_tready_override  \tready_override.f.engine_6_tready_override  \tready_override.f.engine_5_tready_override  \tready_override.f.engine_4_tready_override  \tready_override.f.engine_3_tready_override  \tready_override.f.engine_2_tready_override  \tready_override.f.engine_1_tready_override  \tready_override.f.engine_0_tready_override  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "40"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_NUM "9"
endmodule
