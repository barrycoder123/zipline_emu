
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_sa_counter ( sa_count, sa_snapshot, clk, rst_n, sa_event_sel, 
	.sa_events( {\sa_events[15][63] , \sa_events[15][62] , 
	\sa_events[15][61] , \sa_events[15][60] , \sa_events[15][59] , 
	\sa_events[15][58] , \sa_events[15][57] , \sa_events[15][56] , 
	\sa_events[15][55] , \sa_events[15][54] , \sa_events[15][53] , 
	\sa_events[15][52] , \sa_events[15][51] , \sa_events[15][50] , 
	\sa_events[15][49] , \sa_events[15][48] , \sa_events[15][47] , 
	\sa_events[15][46] , \sa_events[15][45] , \sa_events[15][44] , 
	\sa_events[15][43] , \sa_events[15][42] , \sa_events[15][41] , 
	\sa_events[15][40] , \sa_events[15][39] , \sa_events[15][38] , 
	\sa_events[15][37] , \sa_events[15][36] , \sa_events[15][35] , 
	\sa_events[15][34] , \sa_events[15][33] , \sa_events[15][32] , 
	\sa_events[15][31] , \sa_events[15][30] , \sa_events[15][29] , 
	\sa_events[15][28] , \sa_events[15][27] , \sa_events[15][26] , 
	\sa_events[15][25] , \sa_events[15][24] , \sa_events[15][23] , 
	\sa_events[15][22] , \sa_events[15][21] , \sa_events[15][20] , 
	\sa_events[15][19] , \sa_events[15][18] , \sa_events[15][17] , 
	\sa_events[15][16] , \sa_events[15][15] , \sa_events[15][14] , 
	\sa_events[15][13] , \sa_events[15][12] , \sa_events[15][11] , 
	\sa_events[15][10] , \sa_events[15][9] , \sa_events[15][8] , 
	\sa_events[15][7] , \sa_events[15][6] , \sa_events[15][5] , 
	\sa_events[15][4] , \sa_events[15][3] , \sa_events[15][2] , 
	\sa_events[15][1] , \sa_events[15][0] , \sa_events[14][63] , 
	\sa_events[14][62] , \sa_events[14][61] , \sa_events[14][60] , 
	\sa_events[14][59] , \sa_events[14][58] , \sa_events[14][57] , 
	\sa_events[14][56] , \sa_events[14][55] , \sa_events[14][54] , 
	\sa_events[14][53] , \sa_events[14][52] , \sa_events[14][51] , 
	\sa_events[14][50] , \sa_events[14][49] , \sa_events[14][48] , 
	\sa_events[14][47] , \sa_events[14][46] , \sa_events[14][45] , 
	\sa_events[14][44] , \sa_events[14][43] , \sa_events[14][42] , 
	\sa_events[14][41] , \sa_events[14][40] , \sa_events[14][39] , 
	\sa_events[14][38] , \sa_events[14][37] , \sa_events[14][36] , 
	\sa_events[14][35] , \sa_events[14][34] , \sa_events[14][33] , 
	\sa_events[14][32] , \sa_events[14][31] , \sa_events[14][30] , 
	\sa_events[14][29] , \sa_events[14][28] , \sa_events[14][27] , 
	\sa_events[14][26] , \sa_events[14][25] , \sa_events[14][24] , 
	\sa_events[14][23] , \sa_events[14][22] , \sa_events[14][21] , 
	\sa_events[14][20] , \sa_events[14][19] , \sa_events[14][18] , 
	\sa_events[14][17] , \sa_events[14][16] , \sa_events[14][15] , 
	\sa_events[14][14] , \sa_events[14][13] , \sa_events[14][12] , 
	\sa_events[14][11] , \sa_events[14][10] , \sa_events[14][9] , 
	\sa_events[14][8] , \sa_events[14][7] , \sa_events[14][6] , 
	\sa_events[14][5] , \sa_events[14][4] , \sa_events[14][3] , 
	\sa_events[14][2] , \sa_events[14][1] , \sa_events[14][0] , 
	\sa_events[13][63] , \sa_events[13][62] , \sa_events[13][61] , 
	\sa_events[13][60] , \sa_events[13][59] , \sa_events[13][58] , 
	\sa_events[13][57] , \sa_events[13][56] , \sa_events[13][55] , 
	\sa_events[13][54] , \sa_events[13][53] , \sa_events[13][52] , 
	\sa_events[13][51] , \sa_events[13][50] , \sa_events[13][49] , 
	\sa_events[13][48] , \sa_events[13][47] , \sa_events[13][46] , 
	\sa_events[13][45] , \sa_events[13][44] , \sa_events[13][43] , 
	\sa_events[13][42] , \sa_events[13][41] , \sa_events[13][40] , 
	\sa_events[13][39] , \sa_events[13][38] , \sa_events[13][37] , 
	\sa_events[13][36] , \sa_events[13][35] , \sa_events[13][34] , 
	\sa_events[13][33] , \sa_events[13][32] , \sa_events[13][31] , 
	\sa_events[13][30] , \sa_events[13][29] , \sa_events[13][28] , 
	\sa_events[13][27] , \sa_events[13][26] , \sa_events[13][25] , 
	\sa_events[13][24] , \sa_events[13][23] , \sa_events[13][22] , 
	\sa_events[13][21] , \sa_events[13][20] , \sa_events[13][19] , 
	\sa_events[13][18] , \sa_events[13][17] , \sa_events[13][16] , 
	\sa_events[13][15] , \sa_events[13][14] , \sa_events[13][13] , 
	\sa_events[13][12] , \sa_events[13][11] , \sa_events[13][10] , 
	\sa_events[13][9] , \sa_events[13][8] , \sa_events[13][7] , 
	\sa_events[13][6] , \sa_events[13][5] , \sa_events[13][4] , 
	\sa_events[13][3] , \sa_events[13][2] , \sa_events[13][1] , 
	\sa_events[13][0] , \sa_events[12][63] , \sa_events[12][62] , 
	\sa_events[12][61] , \sa_events[12][60] , \sa_events[12][59] , 
	\sa_events[12][58] , \sa_events[12][57] , \sa_events[12][56] , 
	\sa_events[12][55] , \sa_events[12][54] , \sa_events[12][53] , 
	\sa_events[12][52] , \sa_events[12][51] , \sa_events[12][50] , 
	\sa_events[12][49] , \sa_events[12][48] , \sa_events[12][47] , 
	\sa_events[12][46] , \sa_events[12][45] , \sa_events[12][44] , 
	\sa_events[12][43] , \sa_events[12][42] , \sa_events[12][41] , 
	\sa_events[12][40] , \sa_events[12][39] , \sa_events[12][38] , 
	\sa_events[12][37] , \sa_events[12][36] , \sa_events[12][35] , 
	\sa_events[12][34] , \sa_events[12][33] , \sa_events[12][32] , 
	\sa_events[12][31] , \sa_events[12][30] , \sa_events[12][29] , 
	\sa_events[12][28] , \sa_events[12][27] , \sa_events[12][26] , 
	\sa_events[12][25] , \sa_events[12][24] , \sa_events[12][23] , 
	\sa_events[12][22] , \sa_events[12][21] , \sa_events[12][20] , 
	\sa_events[12][19] , \sa_events[12][18] , \sa_events[12][17] , 
	\sa_events[12][16] , \sa_events[12][15] , \sa_events[12][14] , 
	\sa_events[12][13] , \sa_events[12][12] , \sa_events[12][11] , 
	\sa_events[12][10] , \sa_events[12][9] , \sa_events[12][8] , 
	\sa_events[12][7] , \sa_events[12][6] , \sa_events[12][5] , 
	\sa_events[12][4] , \sa_events[12][3] , \sa_events[12][2] , 
	\sa_events[12][1] , \sa_events[12][0] , \sa_events[11][63] , 
	\sa_events[11][62] , \sa_events[11][61] , \sa_events[11][60] , 
	\sa_events[11][59] , \sa_events[11][58] , \sa_events[11][57] , 
	\sa_events[11][56] , \sa_events[11][55] , \sa_events[11][54] , 
	\sa_events[11][53] , \sa_events[11][52] , \sa_events[11][51] , 
	\sa_events[11][50] , \sa_events[11][49] , \sa_events[11][48] , 
	\sa_events[11][47] , \sa_events[11][46] , \sa_events[11][45] , 
	\sa_events[11][44] , \sa_events[11][43] , \sa_events[11][42] , 
	\sa_events[11][41] , \sa_events[11][40] , \sa_events[11][39] , 
	\sa_events[11][38] , \sa_events[11][37] , \sa_events[11][36] , 
	\sa_events[11][35] , \sa_events[11][34] , \sa_events[11][33] , 
	\sa_events[11][32] , \sa_events[11][31] , \sa_events[11][30] , 
	\sa_events[11][29] , \sa_events[11][28] , \sa_events[11][27] , 
	\sa_events[11][26] , \sa_events[11][25] , \sa_events[11][24] , 
	\sa_events[11][23] , \sa_events[11][22] , \sa_events[11][21] , 
	\sa_events[11][20] , \sa_events[11][19] , \sa_events[11][18] , 
	\sa_events[11][17] , \sa_events[11][16] , \sa_events[11][15] , 
	\sa_events[11][14] , \sa_events[11][13] , \sa_events[11][12] , 
	\sa_events[11][11] , \sa_events[11][10] , \sa_events[11][9] , 
	\sa_events[11][8] , \sa_events[11][7] , \sa_events[11][6] , 
	\sa_events[11][5] , \sa_events[11][4] , \sa_events[11][3] , 
	\sa_events[11][2] , \sa_events[11][1] , \sa_events[11][0] , 
	\sa_events[10][63] , \sa_events[10][62] , \sa_events[10][61] , 
	\sa_events[10][60] , \sa_events[10][59] , \sa_events[10][58] , 
	\sa_events[10][57] , \sa_events[10][56] , \sa_events[10][55] , 
	\sa_events[10][54] , \sa_events[10][53] , \sa_events[10][52] , 
	\sa_events[10][51] , \sa_events[10][50] , \sa_events[10][49] , 
	\sa_events[10][48] , \sa_events[10][47] , \sa_events[10][46] , 
	\sa_events[10][45] , \sa_events[10][44] , \sa_events[10][43] , 
	\sa_events[10][42] , \sa_events[10][41] , \sa_events[10][40] , 
	\sa_events[10][39] , \sa_events[10][38] , \sa_events[10][37] , 
	\sa_events[10][36] , \sa_events[10][35] , \sa_events[10][34] , 
	\sa_events[10][33] , \sa_events[10][32] , \sa_events[10][31] , 
	\sa_events[10][30] , \sa_events[10][29] , \sa_events[10][28] , 
	\sa_events[10][27] , \sa_events[10][26] , \sa_events[10][25] , 
	\sa_events[10][24] , \sa_events[10][23] , \sa_events[10][22] , 
	\sa_events[10][21] , \sa_events[10][20] , \sa_events[10][19] , 
	\sa_events[10][18] , \sa_events[10][17] , \sa_events[10][16] , 
	\sa_events[10][15] , \sa_events[10][14] , \sa_events[10][13] , 
	\sa_events[10][12] , \sa_events[10][11] , \sa_events[10][10] , 
	\sa_events[10][9] , \sa_events[10][8] , \sa_events[10][7] , 
	\sa_events[10][6] , \sa_events[10][5] , \sa_events[10][4] , 
	\sa_events[10][3] , \sa_events[10][2] , \sa_events[10][1] , 
	\sa_events[10][0] , \sa_events[9][63] , \sa_events[9][62] , 
	\sa_events[9][61] , \sa_events[9][60] , \sa_events[9][59] , 
	\sa_events[9][58] , \sa_events[9][57] , \sa_events[9][56] , 
	\sa_events[9][55] , \sa_events[9][54] , \sa_events[9][53] , 
	\sa_events[9][52] , \sa_events[9][51] , \sa_events[9][50] , 
	\sa_events[9][49] , \sa_events[9][48] , \sa_events[9][47] , 
	\sa_events[9][46] , \sa_events[9][45] , \sa_events[9][44] , 
	\sa_events[9][43] , \sa_events[9][42] , \sa_events[9][41] , 
	\sa_events[9][40] , \sa_events[9][39] , \sa_events[9][38] , 
	\sa_events[9][37] , \sa_events[9][36] , \sa_events[9][35] , 
	\sa_events[9][34] , \sa_events[9][33] , \sa_events[9][32] , 
	\sa_events[9][31] , \sa_events[9][30] , \sa_events[9][29] , 
	\sa_events[9][28] , \sa_events[9][27] , \sa_events[9][26] , 
	\sa_events[9][25] , \sa_events[9][24] , \sa_events[9][23] , 
	\sa_events[9][22] , \sa_events[9][21] , \sa_events[9][20] , 
	\sa_events[9][19] , \sa_events[9][18] , \sa_events[9][17] , 
	\sa_events[9][16] , \sa_events[9][15] , \sa_events[9][14] , 
	\sa_events[9][13] , \sa_events[9][12] , \sa_events[9][11] , 
	\sa_events[9][10] , \sa_events[9][9] , \sa_events[9][8] , 
	\sa_events[9][7] , \sa_events[9][6] , \sa_events[9][5] , 
	\sa_events[9][4] , \sa_events[9][3] , \sa_events[9][2] , 
	\sa_events[9][1] , \sa_events[9][0] , \sa_events[8][63] , 
	\sa_events[8][62] , \sa_events[8][61] , \sa_events[8][60] , 
	\sa_events[8][59] , \sa_events[8][58] , \sa_events[8][57] , 
	\sa_events[8][56] , \sa_events[8][55] , \sa_events[8][54] , 
	\sa_events[8][53] , \sa_events[8][52] , \sa_events[8][51] , 
	\sa_events[8][50] , \sa_events[8][49] , \sa_events[8][48] , 
	\sa_events[8][47] , \sa_events[8][46] , \sa_events[8][45] , 
	\sa_events[8][44] , \sa_events[8][43] , \sa_events[8][42] , 
	\sa_events[8][41] , \sa_events[8][40] , \sa_events[8][39] , 
	\sa_events[8][38] , \sa_events[8][37] , \sa_events[8][36] , 
	\sa_events[8][35] , \sa_events[8][34] , \sa_events[8][33] , 
	\sa_events[8][32] , \sa_events[8][31] , \sa_events[8][30] , 
	\sa_events[8][29] , \sa_events[8][28] , \sa_events[8][27] , 
	\sa_events[8][26] , \sa_events[8][25] , \sa_events[8][24] , 
	\sa_events[8][23] , \sa_events[8][22] , \sa_events[8][21] , 
	\sa_events[8][20] , \sa_events[8][19] , \sa_events[8][18] , 
	\sa_events[8][17] , \sa_events[8][16] , \sa_events[8][15] , 
	\sa_events[8][14] , \sa_events[8][13] , \sa_events[8][12] , 
	\sa_events[8][11] , \sa_events[8][10] , \sa_events[8][9] , 
	\sa_events[8][8] , \sa_events[8][7] , \sa_events[8][6] , 
	\sa_events[8][5] , \sa_events[8][4] , \sa_events[8][3] , 
	\sa_events[8][2] , \sa_events[8][1] , \sa_events[8][0] , 
	\sa_events[7][63] , \sa_events[7][62] , \sa_events[7][61] , 
	\sa_events[7][60] , \sa_events[7][59] , \sa_events[7][58] , 
	\sa_events[7][57] , \sa_events[7][56] , \sa_events[7][55] , 
	\sa_events[7][54] , \sa_events[7][53] , \sa_events[7][52] , 
	\sa_events[7][51] , \sa_events[7][50] , \sa_events[7][49] , 
	\sa_events[7][48] , \sa_events[7][47] , \sa_events[7][46] , 
	\sa_events[7][45] , \sa_events[7][44] , \sa_events[7][43] , 
	\sa_events[7][42] , \sa_events[7][41] , \sa_events[7][40] , 
	\sa_events[7][39] , \sa_events[7][38] , \sa_events[7][37] , 
	\sa_events[7][36] , \sa_events[7][35] , \sa_events[7][34] , 
	\sa_events[7][33] , \sa_events[7][32] , \sa_events[7][31] , 
	\sa_events[7][30] , \sa_events[7][29] , \sa_events[7][28] , 
	\sa_events[7][27] , \sa_events[7][26] , \sa_events[7][25] , 
	\sa_events[7][24] , \sa_events[7][23] , \sa_events[7][22] , 
	\sa_events[7][21] , \sa_events[7][20] , \sa_events[7][19] , 
	\sa_events[7][18] , \sa_events[7][17] , \sa_events[7][16] , 
	\sa_events[7][15] , \sa_events[7][14] , \sa_events[7][13] , 
	\sa_events[7][12] , \sa_events[7][11] , \sa_events[7][10] , 
	\sa_events[7][9] , \sa_events[7][8] , \sa_events[7][7] , 
	\sa_events[7][6] , \sa_events[7][5] , \sa_events[7][4] , 
	\sa_events[7][3] , \sa_events[7][2] , \sa_events[7][1] , 
	\sa_events[7][0] , \sa_events[6][63] , \sa_events[6][62] , 
	\sa_events[6][61] , \sa_events[6][60] , \sa_events[6][59] , 
	\sa_events[6][58] , \sa_events[6][57] , \sa_events[6][56] , 
	\sa_events[6][55] , \sa_events[6][54] , \sa_events[6][53] , 
	\sa_events[6][52] , \sa_events[6][51] , \sa_events[6][50] , 
	\sa_events[6][49] , \sa_events[6][48] , \sa_events[6][47] , 
	\sa_events[6][46] , \sa_events[6][45] , \sa_events[6][44] , 
	\sa_events[6][43] , \sa_events[6][42] , \sa_events[6][41] , 
	\sa_events[6][40] , \sa_events[6][39] , \sa_events[6][38] , 
	\sa_events[6][37] , \sa_events[6][36] , \sa_events[6][35] , 
	\sa_events[6][34] , \sa_events[6][33] , \sa_events[6][32] , 
	\sa_events[6][31] , \sa_events[6][30] , \sa_events[6][29] , 
	\sa_events[6][28] , \sa_events[6][27] , \sa_events[6][26] , 
	\sa_events[6][25] , \sa_events[6][24] , \sa_events[6][23] , 
	\sa_events[6][22] , \sa_events[6][21] , \sa_events[6][20] , 
	\sa_events[6][19] , \sa_events[6][18] , \sa_events[6][17] , 
	\sa_events[6][16] , \sa_events[6][15] , \sa_events[6][14] , 
	\sa_events[6][13] , \sa_events[6][12] , \sa_events[6][11] , 
	\sa_events[6][10] , \sa_events[6][9] , \sa_events[6][8] , 
	\sa_events[6][7] , \sa_events[6][6] , \sa_events[6][5] , 
	\sa_events[6][4] , \sa_events[6][3] , \sa_events[6][2] , 
	\sa_events[6][1] , \sa_events[6][0] , \sa_events[5][63] , 
	\sa_events[5][62] , \sa_events[5][61] , \sa_events[5][60] , 
	\sa_events[5][59] , \sa_events[5][58] , \sa_events[5][57] , 
	\sa_events[5][56] , \sa_events[5][55] , \sa_events[5][54] , 
	\sa_events[5][53] , \sa_events[5][52] , \sa_events[5][51] , 
	\sa_events[5][50] , \sa_events[5][49] , \sa_events[5][48] , 
	\sa_events[5][47] , \sa_events[5][46] , \sa_events[5][45] , 
	\sa_events[5][44] , \sa_events[5][43] , \sa_events[5][42] , 
	\sa_events[5][41] , \sa_events[5][40] , \sa_events[5][39] , 
	\sa_events[5][38] , \sa_events[5][37] , \sa_events[5][36] , 
	\sa_events[5][35] , \sa_events[5][34] , \sa_events[5][33] , 
	\sa_events[5][32] , \sa_events[5][31] , \sa_events[5][30] , 
	\sa_events[5][29] , \sa_events[5][28] , \sa_events[5][27] , 
	\sa_events[5][26] , \sa_events[5][25] , \sa_events[5][24] , 
	\sa_events[5][23] , \sa_events[5][22] , \sa_events[5][21] , 
	\sa_events[5][20] , \sa_events[5][19] , \sa_events[5][18] , 
	\sa_events[5][17] , \sa_events[5][16] , \sa_events[5][15] , 
	\sa_events[5][14] , \sa_events[5][13] , \sa_events[5][12] , 
	\sa_events[5][11] , \sa_events[5][10] , \sa_events[5][9] , 
	\sa_events[5][8] , \sa_events[5][7] , \sa_events[5][6] , 
	\sa_events[5][5] , \sa_events[5][4] , \sa_events[5][3] , 
	\sa_events[5][2] , \sa_events[5][1] , \sa_events[5][0] , 
	\sa_events[4][63] , \sa_events[4][62] , \sa_events[4][61] , 
	\sa_events[4][60] , \sa_events[4][59] , \sa_events[4][58] , 
	\sa_events[4][57] , \sa_events[4][56] , \sa_events[4][55] , 
	\sa_events[4][54] , \sa_events[4][53] , \sa_events[4][52] , 
	\sa_events[4][51] , \sa_events[4][50] , \sa_events[4][49] , 
	\sa_events[4][48] , \sa_events[4][47] , \sa_events[4][46] , 
	\sa_events[4][45] , \sa_events[4][44] , \sa_events[4][43] , 
	\sa_events[4][42] , \sa_events[4][41] , \sa_events[4][40] , 
	\sa_events[4][39] , \sa_events[4][38] , \sa_events[4][37] , 
	\sa_events[4][36] , \sa_events[4][35] , \sa_events[4][34] , 
	\sa_events[4][33] , \sa_events[4][32] , \sa_events[4][31] , 
	\sa_events[4][30] , \sa_events[4][29] , \sa_events[4][28] , 
	\sa_events[4][27] , \sa_events[4][26] , \sa_events[4][25] , 
	\sa_events[4][24] , \sa_events[4][23] , \sa_events[4][22] , 
	\sa_events[4][21] , \sa_events[4][20] , \sa_events[4][19] , 
	\sa_events[4][18] , \sa_events[4][17] , \sa_events[4][16] , 
	\sa_events[4][15] , \sa_events[4][14] , \sa_events[4][13] , 
	\sa_events[4][12] , \sa_events[4][11] , \sa_events[4][10] , 
	\sa_events[4][9] , \sa_events[4][8] , \sa_events[4][7] , 
	\sa_events[4][6] , \sa_events[4][5] , \sa_events[4][4] , 
	\sa_events[4][3] , \sa_events[4][2] , \sa_events[4][1] , 
	\sa_events[4][0] , \sa_events[3][63] , \sa_events[3][62] , 
	\sa_events[3][61] , \sa_events[3][60] , \sa_events[3][59] , 
	\sa_events[3][58] , \sa_events[3][57] , \sa_events[3][56] , 
	\sa_events[3][55] , \sa_events[3][54] , \sa_events[3][53] , 
	\sa_events[3][52] , \sa_events[3][51] , \sa_events[3][50] , 
	\sa_events[3][49] , \sa_events[3][48] , \sa_events[3][47] , 
	\sa_events[3][46] , \sa_events[3][45] , \sa_events[3][44] , 
	\sa_events[3][43] , \sa_events[3][42] , \sa_events[3][41] , 
	\sa_events[3][40] , \sa_events[3][39] , \sa_events[3][38] , 
	\sa_events[3][37] , \sa_events[3][36] , \sa_events[3][35] , 
	\sa_events[3][34] , \sa_events[3][33] , \sa_events[3][32] , 
	\sa_events[3][31] , \sa_events[3][30] , \sa_events[3][29] , 
	\sa_events[3][28] , \sa_events[3][27] , \sa_events[3][26] , 
	\sa_events[3][25] , \sa_events[3][24] , \sa_events[3][23] , 
	\sa_events[3][22] , \sa_events[3][21] , \sa_events[3][20] , 
	\sa_events[3][19] , \sa_events[3][18] , \sa_events[3][17] , 
	\sa_events[3][16] , \sa_events[3][15] , \sa_events[3][14] , 
	\sa_events[3][13] , \sa_events[3][12] , \sa_events[3][11] , 
	\sa_events[3][10] , \sa_events[3][9] , \sa_events[3][8] , 
	\sa_events[3][7] , \sa_events[3][6] , \sa_events[3][5] , 
	\sa_events[3][4] , \sa_events[3][3] , \sa_events[3][2] , 
	\sa_events[3][1] , \sa_events[3][0] , \sa_events[2][63] , 
	\sa_events[2][62] , \sa_events[2][61] , \sa_events[2][60] , 
	\sa_events[2][59] , \sa_events[2][58] , \sa_events[2][57] , 
	\sa_events[2][56] , \sa_events[2][55] , \sa_events[2][54] , 
	\sa_events[2][53] , \sa_events[2][52] , \sa_events[2][51] , 
	\sa_events[2][50] , \sa_events[2][49] , \sa_events[2][48] , 
	\sa_events[2][47] , \sa_events[2][46] , \sa_events[2][45] , 
	\sa_events[2][44] , \sa_events[2][43] , \sa_events[2][42] , 
	\sa_events[2][41] , \sa_events[2][40] , \sa_events[2][39] , 
	\sa_events[2][38] , \sa_events[2][37] , \sa_events[2][36] , 
	\sa_events[2][35] , \sa_events[2][34] , \sa_events[2][33] , 
	\sa_events[2][32] , \sa_events[2][31] , \sa_events[2][30] , 
	\sa_events[2][29] , \sa_events[2][28] , \sa_events[2][27] , 
	\sa_events[2][26] , \sa_events[2][25] , \sa_events[2][24] , 
	\sa_events[2][23] , \sa_events[2][22] , \sa_events[2][21] , 
	\sa_events[2][20] , \sa_events[2][19] , \sa_events[2][18] , 
	\sa_events[2][17] , \sa_events[2][16] , \sa_events[2][15] , 
	\sa_events[2][14] , \sa_events[2][13] , \sa_events[2][12] , 
	\sa_events[2][11] , \sa_events[2][10] , \sa_events[2][9] , 
	\sa_events[2][8] , \sa_events[2][7] , \sa_events[2][6] , 
	\sa_events[2][5] , \sa_events[2][4] , \sa_events[2][3] , 
	\sa_events[2][2] , \sa_events[2][1] , \sa_events[2][0] , 
	\sa_events[1][63] , \sa_events[1][62] , \sa_events[1][61] , 
	\sa_events[1][60] , \sa_events[1][59] , \sa_events[1][58] , 
	\sa_events[1][57] , \sa_events[1][56] , \sa_events[1][55] , 
	\sa_events[1][54] , \sa_events[1][53] , \sa_events[1][52] , 
	\sa_events[1][51] , \sa_events[1][50] , \sa_events[1][49] , 
	\sa_events[1][48] , \sa_events[1][47] , \sa_events[1][46] , 
	\sa_events[1][45] , \sa_events[1][44] , \sa_events[1][43] , 
	\sa_events[1][42] , \sa_events[1][41] , \sa_events[1][40] , 
	\sa_events[1][39] , \sa_events[1][38] , \sa_events[1][37] , 
	\sa_events[1][36] , \sa_events[1][35] , \sa_events[1][34] , 
	\sa_events[1][33] , \sa_events[1][32] , \sa_events[1][31] , 
	\sa_events[1][30] , \sa_events[1][29] , \sa_events[1][28] , 
	\sa_events[1][27] , \sa_events[1][26] , \sa_events[1][25] , 
	\sa_events[1][24] , \sa_events[1][23] , \sa_events[1][22] , 
	\sa_events[1][21] , \sa_events[1][20] , \sa_events[1][19] , 
	\sa_events[1][18] , \sa_events[1][17] , \sa_events[1][16] , 
	\sa_events[1][15] , \sa_events[1][14] , \sa_events[1][13] , 
	\sa_events[1][12] , \sa_events[1][11] , \sa_events[1][10] , 
	\sa_events[1][9] , \sa_events[1][8] , \sa_events[1][7] , 
	\sa_events[1][6] , \sa_events[1][5] , \sa_events[1][4] , 
	\sa_events[1][3] , \sa_events[1][2] , \sa_events[1][1] , 
	\sa_events[1][0] , \sa_events[0][63] , \sa_events[0][62] , 
	\sa_events[0][61] , \sa_events[0][60] , \sa_events[0][59] , 
	\sa_events[0][58] , \sa_events[0][57] , \sa_events[0][56] , 
	\sa_events[0][55] , \sa_events[0][54] , \sa_events[0][53] , 
	\sa_events[0][52] , \sa_events[0][51] , \sa_events[0][50] , 
	\sa_events[0][49] , \sa_events[0][48] , \sa_events[0][47] , 
	\sa_events[0][46] , \sa_events[0][45] , \sa_events[0][44] , 
	\sa_events[0][43] , \sa_events[0][42] , \sa_events[0][41] , 
	\sa_events[0][40] , \sa_events[0][39] , \sa_events[0][38] , 
	\sa_events[0][37] , \sa_events[0][36] , \sa_events[0][35] , 
	\sa_events[0][34] , \sa_events[0][33] , \sa_events[0][32] , 
	\sa_events[0][31] , \sa_events[0][30] , \sa_events[0][29] , 
	\sa_events[0][28] , \sa_events[0][27] , \sa_events[0][26] , 
	\sa_events[0][25] , \sa_events[0][24] , \sa_events[0][23] , 
	\sa_events[0][22] , \sa_events[0][21] , \sa_events[0][20] , 
	\sa_events[0][19] , \sa_events[0][18] , \sa_events[0][17] , 
	\sa_events[0][16] , \sa_events[0][15] , \sa_events[0][14] , 
	\sa_events[0][13] , \sa_events[0][12] , \sa_events[0][11] , 
	\sa_events[0][10] , \sa_events[0][9] , \sa_events[0][8] , 
	\sa_events[0][7] , \sa_events[0][6] , \sa_events[0][5] , 
	\sa_events[0][4] , \sa_events[0][3] , \sa_events[0][2] , 
	\sa_events[0][1] , \sa_events[0][0] } ), sa_clear, sa_snap);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [49:0] sa_count;
output [49:0] sa_snapshot;
input clk;
input rst_n;
input [9:0] sa_event_sel;
input \sa_events[15][63] ;
input \sa_events[15][62] ;
input \sa_events[15][61] ;
input \sa_events[15][60] ;
input \sa_events[15][59] ;
input \sa_events[15][58] ;
input \sa_events[15][57] ;
input \sa_events[15][56] ;
input \sa_events[15][55] ;
input \sa_events[15][54] ;
input \sa_events[15][53] ;
input \sa_events[15][52] ;
input \sa_events[15][51] ;
input \sa_events[15][50] ;
input \sa_events[15][49] ;
input \sa_events[15][48] ;
input \sa_events[15][47] ;
input \sa_events[15][46] ;
input \sa_events[15][45] ;
input \sa_events[15][44] ;
input \sa_events[15][43] ;
input \sa_events[15][42] ;
input \sa_events[15][41] ;
input \sa_events[15][40] ;
input \sa_events[15][39] ;
input \sa_events[15][38] ;
input \sa_events[15][37] ;
input \sa_events[15][36] ;
input \sa_events[15][35] ;
input \sa_events[15][34] ;
input \sa_events[15][33] ;
input \sa_events[15][32] ;
input \sa_events[15][31] ;
input \sa_events[15][30] ;
input \sa_events[15][29] ;
input \sa_events[15][28] ;
input \sa_events[15][27] ;
input \sa_events[15][26] ;
input \sa_events[15][25] ;
input \sa_events[15][24] ;
input \sa_events[15][23] ;
input \sa_events[15][22] ;
input \sa_events[15][21] ;
input \sa_events[15][20] ;
input \sa_events[15][19] ;
input \sa_events[15][18] ;
input \sa_events[15][17] ;
input \sa_events[15][16] ;
input \sa_events[15][15] ;
input \sa_events[15][14] ;
input \sa_events[15][13] ;
input \sa_events[15][12] ;
input \sa_events[15][11] ;
input \sa_events[15][10] ;
input \sa_events[15][9] ;
input \sa_events[15][8] ;
input \sa_events[15][7] ;
input \sa_events[15][6] ;
input \sa_events[15][5] ;
input \sa_events[15][4] ;
input \sa_events[15][3] ;
input \sa_events[15][2] ;
input \sa_events[15][1] ;
input \sa_events[15][0] ;
input \sa_events[14][63] ;
input \sa_events[14][62] ;
input \sa_events[14][61] ;
input \sa_events[14][60] ;
input \sa_events[14][59] ;
input \sa_events[14][58] ;
input \sa_events[14][57] ;
input \sa_events[14][56] ;
input \sa_events[14][55] ;
input \sa_events[14][54] ;
input \sa_events[14][53] ;
input \sa_events[14][52] ;
input \sa_events[14][51] ;
input \sa_events[14][50] ;
input \sa_events[14][49] ;
input \sa_events[14][48] ;
input \sa_events[14][47] ;
input \sa_events[14][46] ;
input \sa_events[14][45] ;
input \sa_events[14][44] ;
input \sa_events[14][43] ;
input \sa_events[14][42] ;
input \sa_events[14][41] ;
input \sa_events[14][40] ;
input \sa_events[14][39] ;
input \sa_events[14][38] ;
input \sa_events[14][37] ;
input \sa_events[14][36] ;
input \sa_events[14][35] ;
input \sa_events[14][34] ;
input \sa_events[14][33] ;
input \sa_events[14][32] ;
input \sa_events[14][31] ;
input \sa_events[14][30] ;
input \sa_events[14][29] ;
input \sa_events[14][28] ;
input \sa_events[14][27] ;
input \sa_events[14][26] ;
input \sa_events[14][25] ;
input \sa_events[14][24] ;
input \sa_events[14][23] ;
input \sa_events[14][22] ;
input \sa_events[14][21] ;
input \sa_events[14][20] ;
input \sa_events[14][19] ;
input \sa_events[14][18] ;
input \sa_events[14][17] ;
input \sa_events[14][16] ;
input \sa_events[14][15] ;
input \sa_events[14][14] ;
input \sa_events[14][13] ;
input \sa_events[14][12] ;
input \sa_events[14][11] ;
input \sa_events[14][10] ;
input \sa_events[14][9] ;
input \sa_events[14][8] ;
input \sa_events[14][7] ;
input \sa_events[14][6] ;
input \sa_events[14][5] ;
input \sa_events[14][4] ;
input \sa_events[14][3] ;
input \sa_events[14][2] ;
input \sa_events[14][1] ;
input \sa_events[14][0] ;
input \sa_events[13][63] ;
input \sa_events[13][62] ;
input \sa_events[13][61] ;
input \sa_events[13][60] ;
input \sa_events[13][59] ;
input \sa_events[13][58] ;
input \sa_events[13][57] ;
input \sa_events[13][56] ;
input \sa_events[13][55] ;
input \sa_events[13][54] ;
input \sa_events[13][53] ;
input \sa_events[13][52] ;
input \sa_events[13][51] ;
input \sa_events[13][50] ;
input \sa_events[13][49] ;
input \sa_events[13][48] ;
input \sa_events[13][47] ;
input \sa_events[13][46] ;
input \sa_events[13][45] ;
input \sa_events[13][44] ;
input \sa_events[13][43] ;
input \sa_events[13][42] ;
input \sa_events[13][41] ;
input \sa_events[13][40] ;
input \sa_events[13][39] ;
input \sa_events[13][38] ;
input \sa_events[13][37] ;
input \sa_events[13][36] ;
input \sa_events[13][35] ;
input \sa_events[13][34] ;
input \sa_events[13][33] ;
input \sa_events[13][32] ;
input \sa_events[13][31] ;
input \sa_events[13][30] ;
input \sa_events[13][29] ;
input \sa_events[13][28] ;
input \sa_events[13][27] ;
input \sa_events[13][26] ;
input \sa_events[13][25] ;
input \sa_events[13][24] ;
input \sa_events[13][23] ;
input \sa_events[13][22] ;
input \sa_events[13][21] ;
input \sa_events[13][20] ;
input \sa_events[13][19] ;
input \sa_events[13][18] ;
input \sa_events[13][17] ;
input \sa_events[13][16] ;
input \sa_events[13][15] ;
input \sa_events[13][14] ;
input \sa_events[13][13] ;
input \sa_events[13][12] ;
input \sa_events[13][11] ;
input \sa_events[13][10] ;
input \sa_events[13][9] ;
input \sa_events[13][8] ;
input \sa_events[13][7] ;
input \sa_events[13][6] ;
input \sa_events[13][5] ;
input \sa_events[13][4] ;
input \sa_events[13][3] ;
input \sa_events[13][2] ;
input \sa_events[13][1] ;
input \sa_events[13][0] ;
input \sa_events[12][63] ;
input \sa_events[12][62] ;
input \sa_events[12][61] ;
input \sa_events[12][60] ;
input \sa_events[12][59] ;
input \sa_events[12][58] ;
input \sa_events[12][57] ;
input \sa_events[12][56] ;
input \sa_events[12][55] ;
input \sa_events[12][54] ;
input \sa_events[12][53] ;
input \sa_events[12][52] ;
input \sa_events[12][51] ;
input \sa_events[12][50] ;
input \sa_events[12][49] ;
input \sa_events[12][48] ;
input \sa_events[12][47] ;
input \sa_events[12][46] ;
input \sa_events[12][45] ;
input \sa_events[12][44] ;
input \sa_events[12][43] ;
input \sa_events[12][42] ;
input \sa_events[12][41] ;
input \sa_events[12][40] ;
input \sa_events[12][39] ;
input \sa_events[12][38] ;
input \sa_events[12][37] ;
input \sa_events[12][36] ;
input \sa_events[12][35] ;
input \sa_events[12][34] ;
input \sa_events[12][33] ;
input \sa_events[12][32] ;
input \sa_events[12][31] ;
input \sa_events[12][30] ;
input \sa_events[12][29] ;
input \sa_events[12][28] ;
input \sa_events[12][27] ;
input \sa_events[12][26] ;
input \sa_events[12][25] ;
input \sa_events[12][24] ;
input \sa_events[12][23] ;
input \sa_events[12][22] ;
input \sa_events[12][21] ;
input \sa_events[12][20] ;
input \sa_events[12][19] ;
input \sa_events[12][18] ;
input \sa_events[12][17] ;
input \sa_events[12][16] ;
input \sa_events[12][15] ;
input \sa_events[12][14] ;
input \sa_events[12][13] ;
input \sa_events[12][12] ;
input \sa_events[12][11] ;
input \sa_events[12][10] ;
input \sa_events[12][9] ;
input \sa_events[12][8] ;
input \sa_events[12][7] ;
input \sa_events[12][6] ;
input \sa_events[12][5] ;
input \sa_events[12][4] ;
input \sa_events[12][3] ;
input \sa_events[12][2] ;
input \sa_events[12][1] ;
input \sa_events[12][0] ;
input \sa_events[11][63] ;
input \sa_events[11][62] ;
input \sa_events[11][61] ;
input \sa_events[11][60] ;
input \sa_events[11][59] ;
input \sa_events[11][58] ;
input \sa_events[11][57] ;
input \sa_events[11][56] ;
input \sa_events[11][55] ;
input \sa_events[11][54] ;
input \sa_events[11][53] ;
input \sa_events[11][52] ;
input \sa_events[11][51] ;
input \sa_events[11][50] ;
input \sa_events[11][49] ;
input \sa_events[11][48] ;
input \sa_events[11][47] ;
input \sa_events[11][46] ;
input \sa_events[11][45] ;
input \sa_events[11][44] ;
input \sa_events[11][43] ;
input \sa_events[11][42] ;
input \sa_events[11][41] ;
input \sa_events[11][40] ;
input \sa_events[11][39] ;
input \sa_events[11][38] ;
input \sa_events[11][37] ;
input \sa_events[11][36] ;
input \sa_events[11][35] ;
input \sa_events[11][34] ;
input \sa_events[11][33] ;
input \sa_events[11][32] ;
input \sa_events[11][31] ;
input \sa_events[11][30] ;
input \sa_events[11][29] ;
input \sa_events[11][28] ;
input \sa_events[11][27] ;
input \sa_events[11][26] ;
input \sa_events[11][25] ;
input \sa_events[11][24] ;
input \sa_events[11][23] ;
input \sa_events[11][22] ;
input \sa_events[11][21] ;
input \sa_events[11][20] ;
input \sa_events[11][19] ;
input \sa_events[11][18] ;
input \sa_events[11][17] ;
input \sa_events[11][16] ;
input \sa_events[11][15] ;
input \sa_events[11][14] ;
input \sa_events[11][13] ;
input \sa_events[11][12] ;
input \sa_events[11][11] ;
input \sa_events[11][10] ;
input \sa_events[11][9] ;
input \sa_events[11][8] ;
input \sa_events[11][7] ;
input \sa_events[11][6] ;
input \sa_events[11][5] ;
input \sa_events[11][4] ;
input \sa_events[11][3] ;
input \sa_events[11][2] ;
input \sa_events[11][1] ;
input \sa_events[11][0] ;
input \sa_events[10][63] ;
input \sa_events[10][62] ;
input \sa_events[10][61] ;
input \sa_events[10][60] ;
input \sa_events[10][59] ;
input \sa_events[10][58] ;
input \sa_events[10][57] ;
input \sa_events[10][56] ;
input \sa_events[10][55] ;
input \sa_events[10][54] ;
input \sa_events[10][53] ;
input \sa_events[10][52] ;
input \sa_events[10][51] ;
input \sa_events[10][50] ;
input \sa_events[10][49] ;
input \sa_events[10][48] ;
input \sa_events[10][47] ;
input \sa_events[10][46] ;
input \sa_events[10][45] ;
input \sa_events[10][44] ;
input \sa_events[10][43] ;
input \sa_events[10][42] ;
input \sa_events[10][41] ;
input \sa_events[10][40] ;
input \sa_events[10][39] ;
input \sa_events[10][38] ;
input \sa_events[10][37] ;
input \sa_events[10][36] ;
input \sa_events[10][35] ;
input \sa_events[10][34] ;
input \sa_events[10][33] ;
input \sa_events[10][32] ;
input \sa_events[10][31] ;
input \sa_events[10][30] ;
input \sa_events[10][29] ;
input \sa_events[10][28] ;
input \sa_events[10][27] ;
input \sa_events[10][26] ;
input \sa_events[10][25] ;
input \sa_events[10][24] ;
input \sa_events[10][23] ;
input \sa_events[10][22] ;
input \sa_events[10][21] ;
input \sa_events[10][20] ;
input \sa_events[10][19] ;
input \sa_events[10][18] ;
input \sa_events[10][17] ;
input \sa_events[10][16] ;
input \sa_events[10][15] ;
input \sa_events[10][14] ;
input \sa_events[10][13] ;
input \sa_events[10][12] ;
input \sa_events[10][11] ;
input \sa_events[10][10] ;
input \sa_events[10][9] ;
input \sa_events[10][8] ;
input \sa_events[10][7] ;
input \sa_events[10][6] ;
input \sa_events[10][5] ;
input \sa_events[10][4] ;
input \sa_events[10][3] ;
input \sa_events[10][2] ;
input \sa_events[10][1] ;
input \sa_events[10][0] ;
input \sa_events[9][63] ;
input \sa_events[9][62] ;
input \sa_events[9][61] ;
input \sa_events[9][60] ;
input \sa_events[9][59] ;
input \sa_events[9][58] ;
input \sa_events[9][57] ;
input \sa_events[9][56] ;
input \sa_events[9][55] ;
input \sa_events[9][54] ;
input \sa_events[9][53] ;
input \sa_events[9][52] ;
input \sa_events[9][51] ;
input \sa_events[9][50] ;
input \sa_events[9][49] ;
input \sa_events[9][48] ;
input \sa_events[9][47] ;
input \sa_events[9][46] ;
input \sa_events[9][45] ;
input \sa_events[9][44] ;
input \sa_events[9][43] ;
input \sa_events[9][42] ;
input \sa_events[9][41] ;
input \sa_events[9][40] ;
input \sa_events[9][39] ;
input \sa_events[9][38] ;
input \sa_events[9][37] ;
input \sa_events[9][36] ;
input \sa_events[9][35] ;
input \sa_events[9][34] ;
input \sa_events[9][33] ;
input \sa_events[9][32] ;
input \sa_events[9][31] ;
input \sa_events[9][30] ;
input \sa_events[9][29] ;
input \sa_events[9][28] ;
input \sa_events[9][27] ;
input \sa_events[9][26] ;
input \sa_events[9][25] ;
input \sa_events[9][24] ;
input \sa_events[9][23] ;
input \sa_events[9][22] ;
input \sa_events[9][21] ;
input \sa_events[9][20] ;
input \sa_events[9][19] ;
input \sa_events[9][18] ;
input \sa_events[9][17] ;
input \sa_events[9][16] ;
input \sa_events[9][15] ;
input \sa_events[9][14] ;
input \sa_events[9][13] ;
input \sa_events[9][12] ;
input \sa_events[9][11] ;
input \sa_events[9][10] ;
input \sa_events[9][9] ;
input \sa_events[9][8] ;
input \sa_events[9][7] ;
input \sa_events[9][6] ;
input \sa_events[9][5] ;
input \sa_events[9][4] ;
input \sa_events[9][3] ;
input \sa_events[9][2] ;
input \sa_events[9][1] ;
input \sa_events[9][0] ;
input \sa_events[8][63] ;
input \sa_events[8][62] ;
input \sa_events[8][61] ;
input \sa_events[8][60] ;
input \sa_events[8][59] ;
input \sa_events[8][58] ;
input \sa_events[8][57] ;
input \sa_events[8][56] ;
input \sa_events[8][55] ;
input \sa_events[8][54] ;
input \sa_events[8][53] ;
input \sa_events[8][52] ;
input \sa_events[8][51] ;
input \sa_events[8][50] ;
input \sa_events[8][49] ;
input \sa_events[8][48] ;
input \sa_events[8][47] ;
input \sa_events[8][46] ;
input \sa_events[8][45] ;
input \sa_events[8][44] ;
input \sa_events[8][43] ;
input \sa_events[8][42] ;
input \sa_events[8][41] ;
input \sa_events[8][40] ;
input \sa_events[8][39] ;
input \sa_events[8][38] ;
input \sa_events[8][37] ;
input \sa_events[8][36] ;
input \sa_events[8][35] ;
input \sa_events[8][34] ;
input \sa_events[8][33] ;
input \sa_events[8][32] ;
input \sa_events[8][31] ;
input \sa_events[8][30] ;
input \sa_events[8][29] ;
input \sa_events[8][28] ;
input \sa_events[8][27] ;
input \sa_events[8][26] ;
input \sa_events[8][25] ;
input \sa_events[8][24] ;
input \sa_events[8][23] ;
input \sa_events[8][22] ;
input \sa_events[8][21] ;
input \sa_events[8][20] ;
input \sa_events[8][19] ;
input \sa_events[8][18] ;
input \sa_events[8][17] ;
input \sa_events[8][16] ;
input \sa_events[8][15] ;
input \sa_events[8][14] ;
input \sa_events[8][13] ;
input \sa_events[8][12] ;
input \sa_events[8][11] ;
input \sa_events[8][10] ;
input \sa_events[8][9] ;
input \sa_events[8][8] ;
input \sa_events[8][7] ;
input \sa_events[8][6] ;
input \sa_events[8][5] ;
input \sa_events[8][4] ;
input \sa_events[8][3] ;
input \sa_events[8][2] ;
input \sa_events[8][1] ;
input \sa_events[8][0] ;
input \sa_events[7][63] ;
input \sa_events[7][62] ;
input \sa_events[7][61] ;
input \sa_events[7][60] ;
input \sa_events[7][59] ;
input \sa_events[7][58] ;
input \sa_events[7][57] ;
input \sa_events[7][56] ;
input \sa_events[7][55] ;
input \sa_events[7][54] ;
input \sa_events[7][53] ;
input \sa_events[7][52] ;
input \sa_events[7][51] ;
input \sa_events[7][50] ;
input \sa_events[7][49] ;
input \sa_events[7][48] ;
input \sa_events[7][47] ;
input \sa_events[7][46] ;
input \sa_events[7][45] ;
input \sa_events[7][44] ;
input \sa_events[7][43] ;
input \sa_events[7][42] ;
input \sa_events[7][41] ;
input \sa_events[7][40] ;
input \sa_events[7][39] ;
input \sa_events[7][38] ;
input \sa_events[7][37] ;
input \sa_events[7][36] ;
input \sa_events[7][35] ;
input \sa_events[7][34] ;
input \sa_events[7][33] ;
input \sa_events[7][32] ;
input \sa_events[7][31] ;
input \sa_events[7][30] ;
input \sa_events[7][29] ;
input \sa_events[7][28] ;
input \sa_events[7][27] ;
input \sa_events[7][26] ;
input \sa_events[7][25] ;
input \sa_events[7][24] ;
input \sa_events[7][23] ;
input \sa_events[7][22] ;
input \sa_events[7][21] ;
input \sa_events[7][20] ;
input \sa_events[7][19] ;
input \sa_events[7][18] ;
input \sa_events[7][17] ;
input \sa_events[7][16] ;
input \sa_events[7][15] ;
input \sa_events[7][14] ;
input \sa_events[7][13] ;
input \sa_events[7][12] ;
input \sa_events[7][11] ;
input \sa_events[7][10] ;
input \sa_events[7][9] ;
input \sa_events[7][8] ;
input \sa_events[7][7] ;
input \sa_events[7][6] ;
input \sa_events[7][5] ;
input \sa_events[7][4] ;
input \sa_events[7][3] ;
input \sa_events[7][2] ;
input \sa_events[7][1] ;
input \sa_events[7][0] ;
input \sa_events[6][63] ;
input \sa_events[6][62] ;
input \sa_events[6][61] ;
input \sa_events[6][60] ;
input \sa_events[6][59] ;
input \sa_events[6][58] ;
input \sa_events[6][57] ;
input \sa_events[6][56] ;
input \sa_events[6][55] ;
input \sa_events[6][54] ;
input \sa_events[6][53] ;
input \sa_events[6][52] ;
input \sa_events[6][51] ;
input \sa_events[6][50] ;
input \sa_events[6][49] ;
input \sa_events[6][48] ;
input \sa_events[6][47] ;
input \sa_events[6][46] ;
input \sa_events[6][45] ;
input \sa_events[6][44] ;
input \sa_events[6][43] ;
input \sa_events[6][42] ;
input \sa_events[6][41] ;
input \sa_events[6][40] ;
input \sa_events[6][39] ;
input \sa_events[6][38] ;
input \sa_events[6][37] ;
input \sa_events[6][36] ;
input \sa_events[6][35] ;
input \sa_events[6][34] ;
input \sa_events[6][33] ;
input \sa_events[6][32] ;
input \sa_events[6][31] ;
input \sa_events[6][30] ;
input \sa_events[6][29] ;
input \sa_events[6][28] ;
input \sa_events[6][27] ;
input \sa_events[6][26] ;
input \sa_events[6][25] ;
input \sa_events[6][24] ;
input \sa_events[6][23] ;
input \sa_events[6][22] ;
input \sa_events[6][21] ;
input \sa_events[6][20] ;
input \sa_events[6][19] ;
input \sa_events[6][18] ;
input \sa_events[6][17] ;
input \sa_events[6][16] ;
input \sa_events[6][15] ;
input \sa_events[6][14] ;
input \sa_events[6][13] ;
input \sa_events[6][12] ;
input \sa_events[6][11] ;
input \sa_events[6][10] ;
input \sa_events[6][9] ;
input \sa_events[6][8] ;
input \sa_events[6][7] ;
input \sa_events[6][6] ;
input \sa_events[6][5] ;
input \sa_events[6][4] ;
input \sa_events[6][3] ;
input \sa_events[6][2] ;
input \sa_events[6][1] ;
input \sa_events[6][0] ;
input \sa_events[5][63] ;
input \sa_events[5][62] ;
input \sa_events[5][61] ;
input \sa_events[5][60] ;
input \sa_events[5][59] ;
input \sa_events[5][58] ;
input \sa_events[5][57] ;
input \sa_events[5][56] ;
input \sa_events[5][55] ;
input \sa_events[5][54] ;
input \sa_events[5][53] ;
input \sa_events[5][52] ;
input \sa_events[5][51] ;
input \sa_events[5][50] ;
input \sa_events[5][49] ;
input \sa_events[5][48] ;
input \sa_events[5][47] ;
input \sa_events[5][46] ;
input \sa_events[5][45] ;
input \sa_events[5][44] ;
input \sa_events[5][43] ;
input \sa_events[5][42] ;
input \sa_events[5][41] ;
input \sa_events[5][40] ;
input \sa_events[5][39] ;
input \sa_events[5][38] ;
input \sa_events[5][37] ;
input \sa_events[5][36] ;
input \sa_events[5][35] ;
input \sa_events[5][34] ;
input \sa_events[5][33] ;
input \sa_events[5][32] ;
input \sa_events[5][31] ;
input \sa_events[5][30] ;
input \sa_events[5][29] ;
input \sa_events[5][28] ;
input \sa_events[5][27] ;
input \sa_events[5][26] ;
input \sa_events[5][25] ;
input \sa_events[5][24] ;
input \sa_events[5][23] ;
input \sa_events[5][22] ;
input \sa_events[5][21] ;
input \sa_events[5][20] ;
input \sa_events[5][19] ;
input \sa_events[5][18] ;
input \sa_events[5][17] ;
input \sa_events[5][16] ;
input \sa_events[5][15] ;
input \sa_events[5][14] ;
input \sa_events[5][13] ;
input \sa_events[5][12] ;
input \sa_events[5][11] ;
input \sa_events[5][10] ;
input \sa_events[5][9] ;
input \sa_events[5][8] ;
input \sa_events[5][7] ;
input \sa_events[5][6] ;
input \sa_events[5][5] ;
input \sa_events[5][4] ;
input \sa_events[5][3] ;
input \sa_events[5][2] ;
input \sa_events[5][1] ;
input \sa_events[5][0] ;
input \sa_events[4][63] ;
input \sa_events[4][62] ;
input \sa_events[4][61] ;
input \sa_events[4][60] ;
input \sa_events[4][59] ;
input \sa_events[4][58] ;
input \sa_events[4][57] ;
input \sa_events[4][56] ;
input \sa_events[4][55] ;
input \sa_events[4][54] ;
input \sa_events[4][53] ;
input \sa_events[4][52] ;
input \sa_events[4][51] ;
input \sa_events[4][50] ;
input \sa_events[4][49] ;
input \sa_events[4][48] ;
input \sa_events[4][47] ;
input \sa_events[4][46] ;
input \sa_events[4][45] ;
input \sa_events[4][44] ;
input \sa_events[4][43] ;
input \sa_events[4][42] ;
input \sa_events[4][41] ;
input \sa_events[4][40] ;
input \sa_events[4][39] ;
input \sa_events[4][38] ;
input \sa_events[4][37] ;
input \sa_events[4][36] ;
input \sa_events[4][35] ;
input \sa_events[4][34] ;
input \sa_events[4][33] ;
input \sa_events[4][32] ;
input \sa_events[4][31] ;
input \sa_events[4][30] ;
input \sa_events[4][29] ;
input \sa_events[4][28] ;
input \sa_events[4][27] ;
input \sa_events[4][26] ;
input \sa_events[4][25] ;
input \sa_events[4][24] ;
input \sa_events[4][23] ;
input \sa_events[4][22] ;
input \sa_events[4][21] ;
input \sa_events[4][20] ;
input \sa_events[4][19] ;
input \sa_events[4][18] ;
input \sa_events[4][17] ;
input \sa_events[4][16] ;
input \sa_events[4][15] ;
input \sa_events[4][14] ;
input \sa_events[4][13] ;
input \sa_events[4][12] ;
input \sa_events[4][11] ;
input \sa_events[4][10] ;
input \sa_events[4][9] ;
input \sa_events[4][8] ;
input \sa_events[4][7] ;
input \sa_events[4][6] ;
input \sa_events[4][5] ;
input \sa_events[4][4] ;
input \sa_events[4][3] ;
input \sa_events[4][2] ;
input \sa_events[4][1] ;
input \sa_events[4][0] ;
input \sa_events[3][63] ;
input \sa_events[3][62] ;
input \sa_events[3][61] ;
input \sa_events[3][60] ;
input \sa_events[3][59] ;
input \sa_events[3][58] ;
input \sa_events[3][57] ;
input \sa_events[3][56] ;
input \sa_events[3][55] ;
input \sa_events[3][54] ;
input \sa_events[3][53] ;
input \sa_events[3][52] ;
input \sa_events[3][51] ;
input \sa_events[3][50] ;
input \sa_events[3][49] ;
input \sa_events[3][48] ;
input \sa_events[3][47] ;
input \sa_events[3][46] ;
input \sa_events[3][45] ;
input \sa_events[3][44] ;
input \sa_events[3][43] ;
input \sa_events[3][42] ;
input \sa_events[3][41] ;
input \sa_events[3][40] ;
input \sa_events[3][39] ;
input \sa_events[3][38] ;
input \sa_events[3][37] ;
input \sa_events[3][36] ;
input \sa_events[3][35] ;
input \sa_events[3][34] ;
input \sa_events[3][33] ;
input \sa_events[3][32] ;
input \sa_events[3][31] ;
input \sa_events[3][30] ;
input \sa_events[3][29] ;
input \sa_events[3][28] ;
input \sa_events[3][27] ;
input \sa_events[3][26] ;
input \sa_events[3][25] ;
input \sa_events[3][24] ;
input \sa_events[3][23] ;
input \sa_events[3][22] ;
input \sa_events[3][21] ;
input \sa_events[3][20] ;
input \sa_events[3][19] ;
input \sa_events[3][18] ;
input \sa_events[3][17] ;
input \sa_events[3][16] ;
input \sa_events[3][15] ;
input \sa_events[3][14] ;
input \sa_events[3][13] ;
input \sa_events[3][12] ;
input \sa_events[3][11] ;
input \sa_events[3][10] ;
input \sa_events[3][9] ;
input \sa_events[3][8] ;
input \sa_events[3][7] ;
input \sa_events[3][6] ;
input \sa_events[3][5] ;
input \sa_events[3][4] ;
input \sa_events[3][3] ;
input \sa_events[3][2] ;
input \sa_events[3][1] ;
input \sa_events[3][0] ;
input \sa_events[2][63] ;
input \sa_events[2][62] ;
input \sa_events[2][61] ;
input \sa_events[2][60] ;
input \sa_events[2][59] ;
input \sa_events[2][58] ;
input \sa_events[2][57] ;
input \sa_events[2][56] ;
input \sa_events[2][55] ;
input \sa_events[2][54] ;
input \sa_events[2][53] ;
input \sa_events[2][52] ;
input \sa_events[2][51] ;
input \sa_events[2][50] ;
input \sa_events[2][49] ;
input \sa_events[2][48] ;
input \sa_events[2][47] ;
input \sa_events[2][46] ;
input \sa_events[2][45] ;
input \sa_events[2][44] ;
input \sa_events[2][43] ;
input \sa_events[2][42] ;
input \sa_events[2][41] ;
input \sa_events[2][40] ;
input \sa_events[2][39] ;
input \sa_events[2][38] ;
input \sa_events[2][37] ;
input \sa_events[2][36] ;
input \sa_events[2][35] ;
input \sa_events[2][34] ;
input \sa_events[2][33] ;
input \sa_events[2][32] ;
input \sa_events[2][31] ;
input \sa_events[2][30] ;
input \sa_events[2][29] ;
input \sa_events[2][28] ;
input \sa_events[2][27] ;
input \sa_events[2][26] ;
input \sa_events[2][25] ;
input \sa_events[2][24] ;
input \sa_events[2][23] ;
input \sa_events[2][22] ;
input \sa_events[2][21] ;
input \sa_events[2][20] ;
input \sa_events[2][19] ;
input \sa_events[2][18] ;
input \sa_events[2][17] ;
input \sa_events[2][16] ;
input \sa_events[2][15] ;
input \sa_events[2][14] ;
input \sa_events[2][13] ;
input \sa_events[2][12] ;
input \sa_events[2][11] ;
input \sa_events[2][10] ;
input \sa_events[2][9] ;
input \sa_events[2][8] ;
input \sa_events[2][7] ;
input \sa_events[2][6] ;
input \sa_events[2][5] ;
input \sa_events[2][4] ;
input \sa_events[2][3] ;
input \sa_events[2][2] ;
input \sa_events[2][1] ;
input \sa_events[2][0] ;
input \sa_events[1][63] ;
input \sa_events[1][62] ;
input \sa_events[1][61] ;
input \sa_events[1][60] ;
input \sa_events[1][59] ;
input \sa_events[1][58] ;
input \sa_events[1][57] ;
input \sa_events[1][56] ;
input \sa_events[1][55] ;
input \sa_events[1][54] ;
input \sa_events[1][53] ;
input \sa_events[1][52] ;
input \sa_events[1][51] ;
input \sa_events[1][50] ;
input \sa_events[1][49] ;
input \sa_events[1][48] ;
input \sa_events[1][47] ;
input \sa_events[1][46] ;
input \sa_events[1][45] ;
input \sa_events[1][44] ;
input \sa_events[1][43] ;
input \sa_events[1][42] ;
input \sa_events[1][41] ;
input \sa_events[1][40] ;
input \sa_events[1][39] ;
input \sa_events[1][38] ;
input \sa_events[1][37] ;
input \sa_events[1][36] ;
input \sa_events[1][35] ;
input \sa_events[1][34] ;
input \sa_events[1][33] ;
input \sa_events[1][32] ;
input \sa_events[1][31] ;
input \sa_events[1][30] ;
input \sa_events[1][29] ;
input \sa_events[1][28] ;
input \sa_events[1][27] ;
input \sa_events[1][26] ;
input \sa_events[1][25] ;
input \sa_events[1][24] ;
input \sa_events[1][23] ;
input \sa_events[1][22] ;
input \sa_events[1][21] ;
input \sa_events[1][20] ;
input \sa_events[1][19] ;
input \sa_events[1][18] ;
input \sa_events[1][17] ;
input \sa_events[1][16] ;
input \sa_events[1][15] ;
input \sa_events[1][14] ;
input \sa_events[1][13] ;
input \sa_events[1][12] ;
input \sa_events[1][11] ;
input \sa_events[1][10] ;
input \sa_events[1][9] ;
input \sa_events[1][8] ;
input \sa_events[1][7] ;
input \sa_events[1][6] ;
input \sa_events[1][5] ;
input \sa_events[1][4] ;
input \sa_events[1][3] ;
input \sa_events[1][2] ;
input \sa_events[1][1] ;
input \sa_events[1][0] ;
input \sa_events[0][63] ;
input \sa_events[0][62] ;
input \sa_events[0][61] ;
input \sa_events[0][60] ;
input \sa_events[0][59] ;
input \sa_events[0][58] ;
input \sa_events[0][57] ;
input \sa_events[0][56] ;
input \sa_events[0][55] ;
input \sa_events[0][54] ;
input \sa_events[0][53] ;
input \sa_events[0][52] ;
input \sa_events[0][51] ;
input \sa_events[0][50] ;
input \sa_events[0][49] ;
input \sa_events[0][48] ;
input \sa_events[0][47] ;
input \sa_events[0][46] ;
input \sa_events[0][45] ;
input \sa_events[0][44] ;
input \sa_events[0][43] ;
input \sa_events[0][42] ;
input \sa_events[0][41] ;
input \sa_events[0][40] ;
input \sa_events[0][39] ;
input \sa_events[0][38] ;
input \sa_events[0][37] ;
input \sa_events[0][36] ;
input \sa_events[0][35] ;
input \sa_events[0][34] ;
input \sa_events[0][33] ;
input \sa_events[0][32] ;
input \sa_events[0][31] ;
input \sa_events[0][30] ;
input \sa_events[0][29] ;
input \sa_events[0][28] ;
input \sa_events[0][27] ;
input \sa_events[0][26] ;
input \sa_events[0][25] ;
input \sa_events[0][24] ;
input \sa_events[0][23] ;
input \sa_events[0][22] ;
input \sa_events[0][21] ;
input \sa_events[0][20] ;
input \sa_events[0][19] ;
input \sa_events[0][18] ;
input \sa_events[0][17] ;
input \sa_events[0][16] ;
input \sa_events[0][15] ;
input \sa_events[0][14] ;
input \sa_events[0][13] ;
input \sa_events[0][12] ;
input \sa_events[0][11] ;
input \sa_events[0][10] ;
input \sa_events[0][9] ;
input \sa_events[0][8] ;
input \sa_events[0][7] ;
input \sa_events[0][6] ;
input \sa_events[0][5] ;
input \sa_events[0][4] ;
input \sa_events[0][3] ;
input \sa_events[0][2] ;
input \sa_events[0][1] ;
input \sa_events[0][0] ;
input sa_clear;
input sa_snap;
wire [0:49] _zy_simnet_sa_count_0_w$;
wire [0:49] _zy_simnet_sa_snapshot_1_w$;
wire [63:0] sa_mux1;
wire sa_mux2;
wire [5:0] mux2_sel;
ixc_assign_50 _zz_strnp_3 ( _zy_simnet_sa_snapshot_1_w$[0:49], 
	sa_snapshot[49:0]);
ixc_assign_50 _zz_strnp_2 ( _zy_simnet_sa_count_0_w$[0:49], sa_count[49:0]);
ixc_assign _zz_strnp_1 ( sa_mux2, n9);
Q_MX08 U3 ( .S0(mux2_sel[3]), .S1(mux2_sel[4]), .S2(mux2_sel[5]), .A0(n8), .A1(n7), .A2(n6), .A3(n5), .A4(n4), .A5(n3), .A6(n2), .A7(n1), .Z(n9));
Q_MX08 U4 ( .S0(mux2_sel[0]), .S1(mux2_sel[1]), .S2(mux2_sel[2]), .A0(sa_mux1[0]), .A1(sa_mux1[1]), .A2(sa_mux1[2]), .A3(sa_mux1[3]), .A4(sa_mux1[4]), .A5(sa_mux1[5]), .A6(sa_mux1[6]), .A7(sa_mux1[7]), .Z(n8));
Q_MX08 U5 ( .S0(mux2_sel[0]), .S1(mux2_sel[1]), .S2(mux2_sel[2]), .A0(sa_mux1[8]), .A1(sa_mux1[9]), .A2(sa_mux1[10]), .A3(sa_mux1[11]), .A4(sa_mux1[12]), .A5(sa_mux1[13]), .A6(sa_mux1[14]), .A7(sa_mux1[15]), .Z(n7));
Q_MX08 U6 ( .S0(mux2_sel[0]), .S1(mux2_sel[1]), .S2(mux2_sel[2]), .A0(sa_mux1[16]), .A1(sa_mux1[17]), .A2(sa_mux1[18]), .A3(sa_mux1[19]), .A4(sa_mux1[20]), .A5(sa_mux1[21]), .A6(sa_mux1[22]), .A7(sa_mux1[23]), .Z(n6));
Q_MX08 U7 ( .S0(mux2_sel[0]), .S1(mux2_sel[1]), .S2(mux2_sel[2]), .A0(sa_mux1[24]), .A1(sa_mux1[25]), .A2(sa_mux1[26]), .A3(sa_mux1[27]), .A4(sa_mux1[28]), .A5(sa_mux1[29]), .A6(sa_mux1[30]), .A7(sa_mux1[31]), .Z(n5));
Q_MX08 U8 ( .S0(mux2_sel[0]), .S1(mux2_sel[1]), .S2(mux2_sel[2]), .A0(sa_mux1[32]), .A1(sa_mux1[33]), .A2(sa_mux1[34]), .A3(sa_mux1[35]), .A4(sa_mux1[36]), .A5(sa_mux1[37]), .A6(sa_mux1[38]), .A7(sa_mux1[39]), .Z(n4));
Q_MX08 U9 ( .S0(mux2_sel[0]), .S1(mux2_sel[1]), .S2(mux2_sel[2]), .A0(sa_mux1[40]), .A1(sa_mux1[41]), .A2(sa_mux1[42]), .A3(sa_mux1[43]), .A4(sa_mux1[44]), .A5(sa_mux1[45]), .A6(sa_mux1[46]), .A7(sa_mux1[47]), .Z(n3));
Q_MX08 U10 ( .S0(mux2_sel[0]), .S1(mux2_sel[1]), .S2(mux2_sel[2]), .A0(sa_mux1[48]), .A1(sa_mux1[49]), .A2(sa_mux1[50]), .A3(sa_mux1[51]), .A4(sa_mux1[52]), .A5(sa_mux1[53]), .A6(sa_mux1[54]), .A7(sa_mux1[55]), .Z(n2));
Q_MX08 U11 ( .S0(mux2_sel[0]), .S1(mux2_sel[1]), .S2(mux2_sel[2]), .A0(sa_mux1[56]), .A1(sa_mux1[57]), .A2(sa_mux1[58]), .A3(sa_mux1[59]), .A4(sa_mux1[60]), .A5(sa_mux1[61]), .A6(sa_mux1[62]), .A7(sa_mux1[63]), .Z(n1));
ixc_assign_6 _zz_strnp_0 ( mux2_sel[5:0], sa_event_sel[5:0]);
Q_AD01HF U13 ( .A0(sa_count[1]), .B0(sa_count[0]), .S(n10), .CO(n11));
Q_AD01HF U14 ( .A0(sa_count[2]), .B0(n11), .S(n12), .CO(n13));
Q_AD01HF U15 ( .A0(sa_count[3]), .B0(n13), .S(n14), .CO(n15));
Q_AD01HF U16 ( .A0(sa_count[4]), .B0(n15), .S(n16), .CO(n17));
Q_AD01HF U17 ( .A0(sa_count[5]), .B0(n17), .S(n18), .CO(n19));
Q_AD01HF U18 ( .A0(sa_count[6]), .B0(n19), .S(n20), .CO(n21));
Q_AD01HF U19 ( .A0(sa_count[7]), .B0(n21), .S(n22), .CO(n23));
Q_AD01HF U20 ( .A0(sa_count[8]), .B0(n23), .S(n24), .CO(n25));
Q_AD01HF U21 ( .A0(sa_count[9]), .B0(n25), .S(n26), .CO(n27));
Q_AD01HF U22 ( .A0(sa_count[10]), .B0(n27), .S(n28), .CO(n29));
Q_AD01HF U23 ( .A0(sa_count[11]), .B0(n29), .S(n30), .CO(n31));
Q_AD01HF U24 ( .A0(sa_count[12]), .B0(n31), .S(n32), .CO(n33));
Q_AD01HF U25 ( .A0(sa_count[13]), .B0(n33), .S(n34), .CO(n35));
Q_AD01HF U26 ( .A0(sa_count[14]), .B0(n35), .S(n36), .CO(n37));
Q_AD01HF U27 ( .A0(sa_count[15]), .B0(n37), .S(n38), .CO(n39));
Q_AD01HF U28 ( .A0(sa_count[16]), .B0(n39), .S(n40), .CO(n41));
Q_AD01HF U29 ( .A0(sa_count[17]), .B0(n41), .S(n42), .CO(n43));
Q_AD01HF U30 ( .A0(sa_count[18]), .B0(n43), .S(n44), .CO(n45));
Q_AD01HF U31 ( .A0(sa_count[19]), .B0(n45), .S(n46), .CO(n47));
Q_AD01HF U32 ( .A0(sa_count[20]), .B0(n47), .S(n48), .CO(n49));
Q_AD01HF U33 ( .A0(sa_count[21]), .B0(n49), .S(n50), .CO(n51));
Q_AD01HF U34 ( .A0(sa_count[22]), .B0(n51), .S(n52), .CO(n53));
Q_AD01HF U35 ( .A0(sa_count[23]), .B0(n53), .S(n54), .CO(n55));
Q_AD01HF U36 ( .A0(sa_count[24]), .B0(n55), .S(n56), .CO(n57));
Q_AD01HF U37 ( .A0(sa_count[25]), .B0(n57), .S(n58), .CO(n59));
Q_AD01HF U38 ( .A0(sa_count[26]), .B0(n59), .S(n60), .CO(n61));
Q_AD01HF U39 ( .A0(sa_count[27]), .B0(n61), .S(n62), .CO(n63));
Q_AD01HF U40 ( .A0(sa_count[28]), .B0(n63), .S(n64), .CO(n65));
Q_AD01HF U41 ( .A0(sa_count[29]), .B0(n65), .S(n66), .CO(n67));
Q_AD01HF U42 ( .A0(sa_count[30]), .B0(n67), .S(n68), .CO(n69));
Q_AD01HF U43 ( .A0(sa_count[31]), .B0(n69), .S(n70), .CO(n71));
Q_AD01HF U44 ( .A0(sa_count[32]), .B0(n71), .S(n72), .CO(n73));
Q_AD01HF U45 ( .A0(sa_count[33]), .B0(n73), .S(n74), .CO(n75));
Q_AD01HF U46 ( .A0(sa_count[34]), .B0(n75), .S(n76), .CO(n77));
Q_AD01HF U47 ( .A0(sa_count[35]), .B0(n77), .S(n78), .CO(n79));
Q_AD01HF U48 ( .A0(sa_count[36]), .B0(n79), .S(n80), .CO(n81));
Q_AD01HF U49 ( .A0(sa_count[37]), .B0(n81), .S(n82), .CO(n83));
Q_AD01HF U50 ( .A0(sa_count[38]), .B0(n83), .S(n84), .CO(n85));
Q_AD01HF U51 ( .A0(sa_count[39]), .B0(n85), .S(n86), .CO(n87));
Q_AD01HF U52 ( .A0(sa_count[40]), .B0(n87), .S(n88), .CO(n89));
Q_AD01HF U53 ( .A0(sa_count[41]), .B0(n89), .S(n90), .CO(n91));
Q_AD01HF U54 ( .A0(sa_count[42]), .B0(n91), .S(n92), .CO(n93));
Q_AD01HF U55 ( .A0(sa_count[43]), .B0(n93), .S(n94), .CO(n95));
Q_AD01HF U56 ( .A0(sa_count[44]), .B0(n95), .S(n96), .CO(n97));
Q_AD01HF U57 ( .A0(sa_count[45]), .B0(n97), .S(n98), .CO(n99));
Q_AD01HF U58 ( .A0(sa_count[46]), .B0(n99), .S(n100), .CO(n101));
Q_AD01HF U59 ( .A0(sa_count[47]), .B0(n101), .S(n102), .CO(n103));
Q_AD01HF U60 ( .A0(sa_count[48]), .B0(n103), .S(n104), .CO(n105));
Q_XOR2 U61 ( .A0(sa_count[49]), .A1(n105), .Z(n106));
Q_NR02 U62 ( .A0(sa_clear), .A1(sa_count[0]), .Z(n107));
Q_AN02 U63 ( .A0(n158), .A1(n10), .Z(n108));
Q_AN02 U64 ( .A0(n158), .A1(n12), .Z(n109));
Q_AN02 U65 ( .A0(n158), .A1(n14), .Z(n110));
Q_AN02 U66 ( .A0(n158), .A1(n16), .Z(n111));
Q_AN02 U67 ( .A0(n158), .A1(n18), .Z(n112));
Q_AN02 U68 ( .A0(n158), .A1(n20), .Z(n113));
Q_AN02 U69 ( .A0(n158), .A1(n22), .Z(n114));
Q_AN02 U70 ( .A0(n158), .A1(n24), .Z(n115));
Q_AN02 U71 ( .A0(n158), .A1(n26), .Z(n116));
Q_AN02 U72 ( .A0(n158), .A1(n28), .Z(n117));
Q_AN02 U73 ( .A0(n158), .A1(n30), .Z(n118));
Q_AN02 U74 ( .A0(n158), .A1(n32), .Z(n119));
Q_AN02 U75 ( .A0(n158), .A1(n34), .Z(n120));
Q_AN02 U76 ( .A0(n158), .A1(n36), .Z(n121));
Q_AN02 U77 ( .A0(n158), .A1(n38), .Z(n122));
Q_AN02 U78 ( .A0(n158), .A1(n40), .Z(n123));
Q_AN02 U79 ( .A0(n158), .A1(n42), .Z(n124));
Q_AN02 U80 ( .A0(n158), .A1(n44), .Z(n125));
Q_AN02 U81 ( .A0(n158), .A1(n46), .Z(n126));
Q_AN02 U82 ( .A0(n158), .A1(n48), .Z(n127));
Q_AN02 U83 ( .A0(n158), .A1(n50), .Z(n128));
Q_AN02 U84 ( .A0(n158), .A1(n52), .Z(n129));
Q_AN02 U85 ( .A0(n158), .A1(n54), .Z(n130));
Q_AN02 U86 ( .A0(n158), .A1(n56), .Z(n131));
Q_AN02 U87 ( .A0(n158), .A1(n58), .Z(n132));
Q_AN02 U88 ( .A0(n158), .A1(n60), .Z(n133));
Q_AN02 U89 ( .A0(n158), .A1(n62), .Z(n134));
Q_AN02 U90 ( .A0(n158), .A1(n64), .Z(n135));
Q_AN02 U91 ( .A0(n158), .A1(n66), .Z(n136));
Q_AN02 U92 ( .A0(n158), .A1(n68), .Z(n137));
Q_AN02 U93 ( .A0(n158), .A1(n70), .Z(n138));
Q_AN02 U94 ( .A0(n158), .A1(n72), .Z(n139));
Q_AN02 U95 ( .A0(n158), .A1(n74), .Z(n140));
Q_AN02 U96 ( .A0(n158), .A1(n76), .Z(n141));
Q_AN02 U97 ( .A0(n158), .A1(n78), .Z(n142));
Q_AN02 U98 ( .A0(n158), .A1(n80), .Z(n143));
Q_AN02 U99 ( .A0(n158), .A1(n82), .Z(n144));
Q_AN02 U100 ( .A0(n158), .A1(n84), .Z(n145));
Q_AN02 U101 ( .A0(n158), .A1(n86), .Z(n146));
Q_AN02 U102 ( .A0(n158), .A1(n88), .Z(n147));
Q_AN02 U103 ( .A0(n158), .A1(n90), .Z(n148));
Q_AN02 U104 ( .A0(n158), .A1(n92), .Z(n149));
Q_AN02 U105 ( .A0(n158), .A1(n94), .Z(n150));
Q_AN02 U106 ( .A0(n158), .A1(n96), .Z(n151));
Q_AN02 U107 ( .A0(n158), .A1(n98), .Z(n152));
Q_AN02 U108 ( .A0(n158), .A1(n100), .Z(n153));
Q_AN02 U109 ( .A0(n158), .A1(n102), .Z(n154));
Q_AN02 U110 ( .A0(n158), .A1(n104), .Z(n155));
Q_AN02 U111 ( .A0(n158), .A1(n106), .Z(n156));
Q_INV U112 ( .A(n157), .Z(n159));
Q_NR02 U113 ( .A0(sa_clear), .A1(sa_mux2), .Z(n157));
Q_INV U114 ( .A(sa_clear), .Z(n158));
Q_MX04 U115 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][0] ), .A1(\sa_events[13][0] ), .A2(\sa_events[14][0] ), .A3(\sa_events[15][0] ), .Z(n160));
Q_MX04 U116 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][0] ), .A1(\sa_events[9][0] ), .A2(\sa_events[10][0] ), .A3(\sa_events[11][0] ), .Z(n161));
Q_MX04 U117 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][0] ), .A1(\sa_events[5][0] ), .A2(\sa_events[6][0] ), .A3(\sa_events[7][0] ), .Z(n162));
Q_MX04 U118 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][0] ), .A1(\sa_events[1][0] ), .A2(\sa_events[2][0] ), .A3(\sa_events[3][0] ), .Z(n163));
Q_MX04 U119 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n163), .A1(n162), .A2(n161), .A3(n160), .Z(sa_mux1[0]));
Q_MX04 U120 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][1] ), .A1(\sa_events[13][1] ), .A2(\sa_events[14][1] ), .A3(\sa_events[15][1] ), .Z(n164));
Q_MX04 U121 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][1] ), .A1(\sa_events[9][1] ), .A2(\sa_events[10][1] ), .A3(\sa_events[11][1] ), .Z(n165));
Q_MX04 U122 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][1] ), .A1(\sa_events[5][1] ), .A2(\sa_events[6][1] ), .A3(\sa_events[7][1] ), .Z(n166));
Q_MX04 U123 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][1] ), .A1(\sa_events[1][1] ), .A2(\sa_events[2][1] ), .A3(\sa_events[3][1] ), .Z(n167));
Q_MX04 U124 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n167), .A1(n166), .A2(n165), .A3(n164), .Z(sa_mux1[1]));
Q_MX04 U125 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][2] ), .A1(\sa_events[13][2] ), .A2(\sa_events[14][2] ), .A3(\sa_events[15][2] ), .Z(n168));
Q_MX04 U126 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][2] ), .A1(\sa_events[9][2] ), .A2(\sa_events[10][2] ), .A3(\sa_events[11][2] ), .Z(n169));
Q_MX04 U127 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][2] ), .A1(\sa_events[5][2] ), .A2(\sa_events[6][2] ), .A3(\sa_events[7][2] ), .Z(n170));
Q_MX04 U128 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][2] ), .A1(\sa_events[1][2] ), .A2(\sa_events[2][2] ), .A3(\sa_events[3][2] ), .Z(n171));
Q_MX04 U129 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n171), .A1(n170), .A2(n169), .A3(n168), .Z(sa_mux1[2]));
Q_MX04 U130 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][3] ), .A1(\sa_events[13][3] ), .A2(\sa_events[14][3] ), .A3(\sa_events[15][3] ), .Z(n172));
Q_MX04 U131 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][3] ), .A1(\sa_events[9][3] ), .A2(\sa_events[10][3] ), .A3(\sa_events[11][3] ), .Z(n173));
Q_MX04 U132 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][3] ), .A1(\sa_events[5][3] ), .A2(\sa_events[6][3] ), .A3(\sa_events[7][3] ), .Z(n174));
Q_MX04 U133 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][3] ), .A1(\sa_events[1][3] ), .A2(\sa_events[2][3] ), .A3(\sa_events[3][3] ), .Z(n175));
Q_MX04 U134 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n175), .A1(n174), .A2(n173), .A3(n172), .Z(sa_mux1[3]));
Q_MX04 U135 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][4] ), .A1(\sa_events[13][4] ), .A2(\sa_events[14][4] ), .A3(\sa_events[15][4] ), .Z(n176));
Q_MX04 U136 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][4] ), .A1(\sa_events[9][4] ), .A2(\sa_events[10][4] ), .A3(\sa_events[11][4] ), .Z(n177));
Q_MX04 U137 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][4] ), .A1(\sa_events[5][4] ), .A2(\sa_events[6][4] ), .A3(\sa_events[7][4] ), .Z(n178));
Q_MX04 U138 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][4] ), .A1(\sa_events[1][4] ), .A2(\sa_events[2][4] ), .A3(\sa_events[3][4] ), .Z(n179));
Q_MX04 U139 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n179), .A1(n178), .A2(n177), .A3(n176), .Z(sa_mux1[4]));
Q_MX04 U140 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][5] ), .A1(\sa_events[13][5] ), .A2(\sa_events[14][5] ), .A3(\sa_events[15][5] ), .Z(n180));
Q_MX04 U141 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][5] ), .A1(\sa_events[9][5] ), .A2(\sa_events[10][5] ), .A3(\sa_events[11][5] ), .Z(n181));
Q_MX04 U142 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][5] ), .A1(\sa_events[5][5] ), .A2(\sa_events[6][5] ), .A3(\sa_events[7][5] ), .Z(n182));
Q_MX04 U143 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][5] ), .A1(\sa_events[1][5] ), .A2(\sa_events[2][5] ), .A3(\sa_events[3][5] ), .Z(n183));
Q_MX04 U144 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n183), .A1(n182), .A2(n181), .A3(n180), .Z(sa_mux1[5]));
Q_MX04 U145 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][6] ), .A1(\sa_events[13][6] ), .A2(\sa_events[14][6] ), .A3(\sa_events[15][6] ), .Z(n184));
Q_MX04 U146 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][6] ), .A1(\sa_events[9][6] ), .A2(\sa_events[10][6] ), .A3(\sa_events[11][6] ), .Z(n185));
Q_MX04 U147 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][6] ), .A1(\sa_events[5][6] ), .A2(\sa_events[6][6] ), .A3(\sa_events[7][6] ), .Z(n186));
Q_MX04 U148 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][6] ), .A1(\sa_events[1][6] ), .A2(\sa_events[2][6] ), .A3(\sa_events[3][6] ), .Z(n187));
Q_MX04 U149 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n187), .A1(n186), .A2(n185), .A3(n184), .Z(sa_mux1[6]));
Q_MX04 U150 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][7] ), .A1(\sa_events[13][7] ), .A2(\sa_events[14][7] ), .A3(\sa_events[15][7] ), .Z(n188));
Q_MX04 U151 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][7] ), .A1(\sa_events[9][7] ), .A2(\sa_events[10][7] ), .A3(\sa_events[11][7] ), .Z(n189));
Q_MX04 U152 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][7] ), .A1(\sa_events[5][7] ), .A2(\sa_events[6][7] ), .A3(\sa_events[7][7] ), .Z(n190));
Q_MX04 U153 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][7] ), .A1(\sa_events[1][7] ), .A2(\sa_events[2][7] ), .A3(\sa_events[3][7] ), .Z(n191));
Q_MX04 U154 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n191), .A1(n190), .A2(n189), .A3(n188), .Z(sa_mux1[7]));
Q_MX04 U155 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][8] ), .A1(\sa_events[13][8] ), .A2(\sa_events[14][8] ), .A3(\sa_events[15][8] ), .Z(n192));
Q_MX04 U156 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][8] ), .A1(\sa_events[9][8] ), .A2(\sa_events[10][8] ), .A3(\sa_events[11][8] ), .Z(n193));
Q_MX04 U157 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][8] ), .A1(\sa_events[5][8] ), .A2(\sa_events[6][8] ), .A3(\sa_events[7][8] ), .Z(n194));
Q_MX04 U158 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][8] ), .A1(\sa_events[1][8] ), .A2(\sa_events[2][8] ), .A3(\sa_events[3][8] ), .Z(n195));
Q_MX04 U159 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n195), .A1(n194), .A2(n193), .A3(n192), .Z(sa_mux1[8]));
Q_MX04 U160 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][9] ), .A1(\sa_events[13][9] ), .A2(\sa_events[14][9] ), .A3(\sa_events[15][9] ), .Z(n196));
Q_MX04 U161 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][9] ), .A1(\sa_events[9][9] ), .A2(\sa_events[10][9] ), .A3(\sa_events[11][9] ), .Z(n197));
Q_MX04 U162 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][9] ), .A1(\sa_events[5][9] ), .A2(\sa_events[6][9] ), .A3(\sa_events[7][9] ), .Z(n198));
Q_MX04 U163 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][9] ), .A1(\sa_events[1][9] ), .A2(\sa_events[2][9] ), .A3(\sa_events[3][9] ), .Z(n199));
Q_MX04 U164 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n199), .A1(n198), .A2(n197), .A3(n196), .Z(sa_mux1[9]));
Q_MX04 U165 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][10] ), .A1(\sa_events[13][10] ), .A2(\sa_events[14][10] ), .A3(\sa_events[15][10] ), .Z(n200));
Q_MX04 U166 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][10] ), .A1(\sa_events[9][10] ), .A2(\sa_events[10][10] ), .A3(\sa_events[11][10] ), .Z(n201));
Q_MX04 U167 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][10] ), .A1(\sa_events[5][10] ), .A2(\sa_events[6][10] ), .A3(\sa_events[7][10] ), .Z(n202));
Q_MX04 U168 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][10] ), .A1(\sa_events[1][10] ), .A2(\sa_events[2][10] ), .A3(\sa_events[3][10] ), .Z(n203));
Q_MX04 U169 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n203), .A1(n202), .A2(n201), .A3(n200), .Z(sa_mux1[10]));
Q_MX04 U170 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][11] ), .A1(\sa_events[13][11] ), .A2(\sa_events[14][11] ), .A3(\sa_events[15][11] ), .Z(n204));
Q_MX04 U171 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][11] ), .A1(\sa_events[9][11] ), .A2(\sa_events[10][11] ), .A3(\sa_events[11][11] ), .Z(n205));
Q_MX04 U172 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][11] ), .A1(\sa_events[5][11] ), .A2(\sa_events[6][11] ), .A3(\sa_events[7][11] ), .Z(n206));
Q_MX04 U173 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][11] ), .A1(\sa_events[1][11] ), .A2(\sa_events[2][11] ), .A3(\sa_events[3][11] ), .Z(n207));
Q_MX04 U174 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n207), .A1(n206), .A2(n205), .A3(n204), .Z(sa_mux1[11]));
Q_MX04 U175 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][12] ), .A1(\sa_events[13][12] ), .A2(\sa_events[14][12] ), .A3(\sa_events[15][12] ), .Z(n208));
Q_MX04 U176 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][12] ), .A1(\sa_events[9][12] ), .A2(\sa_events[10][12] ), .A3(\sa_events[11][12] ), .Z(n209));
Q_MX04 U177 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][12] ), .A1(\sa_events[5][12] ), .A2(\sa_events[6][12] ), .A3(\sa_events[7][12] ), .Z(n210));
Q_MX04 U178 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][12] ), .A1(\sa_events[1][12] ), .A2(\sa_events[2][12] ), .A3(\sa_events[3][12] ), .Z(n211));
Q_MX04 U179 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n211), .A1(n210), .A2(n209), .A3(n208), .Z(sa_mux1[12]));
Q_MX04 U180 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][13] ), .A1(\sa_events[13][13] ), .A2(\sa_events[14][13] ), .A3(\sa_events[15][13] ), .Z(n212));
Q_MX04 U181 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][13] ), .A1(\sa_events[9][13] ), .A2(\sa_events[10][13] ), .A3(\sa_events[11][13] ), .Z(n213));
Q_MX04 U182 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][13] ), .A1(\sa_events[5][13] ), .A2(\sa_events[6][13] ), .A3(\sa_events[7][13] ), .Z(n214));
Q_MX04 U183 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][13] ), .A1(\sa_events[1][13] ), .A2(\sa_events[2][13] ), .A3(\sa_events[3][13] ), .Z(n215));
Q_MX04 U184 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n215), .A1(n214), .A2(n213), .A3(n212), .Z(sa_mux1[13]));
Q_MX04 U185 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][14] ), .A1(\sa_events[13][14] ), .A2(\sa_events[14][14] ), .A3(\sa_events[15][14] ), .Z(n216));
Q_MX04 U186 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][14] ), .A1(\sa_events[9][14] ), .A2(\sa_events[10][14] ), .A3(\sa_events[11][14] ), .Z(n217));
Q_MX04 U187 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][14] ), .A1(\sa_events[5][14] ), .A2(\sa_events[6][14] ), .A3(\sa_events[7][14] ), .Z(n218));
Q_MX04 U188 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][14] ), .A1(\sa_events[1][14] ), .A2(\sa_events[2][14] ), .A3(\sa_events[3][14] ), .Z(n219));
Q_MX04 U189 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n219), .A1(n218), .A2(n217), .A3(n216), .Z(sa_mux1[14]));
Q_MX04 U190 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][15] ), .A1(\sa_events[13][15] ), .A2(\sa_events[14][15] ), .A3(\sa_events[15][15] ), .Z(n220));
Q_MX04 U191 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][15] ), .A1(\sa_events[9][15] ), .A2(\sa_events[10][15] ), .A3(\sa_events[11][15] ), .Z(n221));
Q_MX04 U192 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][15] ), .A1(\sa_events[5][15] ), .A2(\sa_events[6][15] ), .A3(\sa_events[7][15] ), .Z(n222));
Q_MX04 U193 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][15] ), .A1(\sa_events[1][15] ), .A2(\sa_events[2][15] ), .A3(\sa_events[3][15] ), .Z(n223));
Q_MX04 U194 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n223), .A1(n222), .A2(n221), .A3(n220), .Z(sa_mux1[15]));
Q_MX04 U195 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][16] ), .A1(\sa_events[13][16] ), .A2(\sa_events[14][16] ), .A3(\sa_events[15][16] ), .Z(n224));
Q_MX04 U196 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][16] ), .A1(\sa_events[9][16] ), .A2(\sa_events[10][16] ), .A3(\sa_events[11][16] ), .Z(n225));
Q_MX04 U197 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][16] ), .A1(\sa_events[5][16] ), .A2(\sa_events[6][16] ), .A3(\sa_events[7][16] ), .Z(n226));
Q_MX04 U198 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][16] ), .A1(\sa_events[1][16] ), .A2(\sa_events[2][16] ), .A3(\sa_events[3][16] ), .Z(n227));
Q_MX04 U199 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n227), .A1(n226), .A2(n225), .A3(n224), .Z(sa_mux1[16]));
Q_MX04 U200 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][17] ), .A1(\sa_events[13][17] ), .A2(\sa_events[14][17] ), .A3(\sa_events[15][17] ), .Z(n228));
Q_MX04 U201 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][17] ), .A1(\sa_events[9][17] ), .A2(\sa_events[10][17] ), .A3(\sa_events[11][17] ), .Z(n229));
Q_MX04 U202 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][17] ), .A1(\sa_events[5][17] ), .A2(\sa_events[6][17] ), .A3(\sa_events[7][17] ), .Z(n230));
Q_MX04 U203 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][17] ), .A1(\sa_events[1][17] ), .A2(\sa_events[2][17] ), .A3(\sa_events[3][17] ), .Z(n231));
Q_MX04 U204 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n231), .A1(n230), .A2(n229), .A3(n228), .Z(sa_mux1[17]));
Q_MX04 U205 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][18] ), .A1(\sa_events[13][18] ), .A2(\sa_events[14][18] ), .A3(\sa_events[15][18] ), .Z(n232));
Q_MX04 U206 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][18] ), .A1(\sa_events[9][18] ), .A2(\sa_events[10][18] ), .A3(\sa_events[11][18] ), .Z(n233));
Q_MX04 U207 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][18] ), .A1(\sa_events[5][18] ), .A2(\sa_events[6][18] ), .A3(\sa_events[7][18] ), .Z(n234));
Q_MX04 U208 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][18] ), .A1(\sa_events[1][18] ), .A2(\sa_events[2][18] ), .A3(\sa_events[3][18] ), .Z(n235));
Q_MX04 U209 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n235), .A1(n234), .A2(n233), .A3(n232), .Z(sa_mux1[18]));
Q_MX04 U210 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][19] ), .A1(\sa_events[13][19] ), .A2(\sa_events[14][19] ), .A3(\sa_events[15][19] ), .Z(n236));
Q_MX04 U211 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][19] ), .A1(\sa_events[9][19] ), .A2(\sa_events[10][19] ), .A3(\sa_events[11][19] ), .Z(n237));
Q_MX04 U212 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][19] ), .A1(\sa_events[5][19] ), .A2(\sa_events[6][19] ), .A3(\sa_events[7][19] ), .Z(n238));
Q_MX04 U213 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][19] ), .A1(\sa_events[1][19] ), .A2(\sa_events[2][19] ), .A3(\sa_events[3][19] ), .Z(n239));
Q_MX04 U214 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n239), .A1(n238), .A2(n237), .A3(n236), .Z(sa_mux1[19]));
Q_MX04 U215 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][20] ), .A1(\sa_events[13][20] ), .A2(\sa_events[14][20] ), .A3(\sa_events[15][20] ), .Z(n240));
Q_MX04 U216 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][20] ), .A1(\sa_events[9][20] ), .A2(\sa_events[10][20] ), .A3(\sa_events[11][20] ), .Z(n241));
Q_MX04 U217 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][20] ), .A1(\sa_events[5][20] ), .A2(\sa_events[6][20] ), .A3(\sa_events[7][20] ), .Z(n242));
Q_MX04 U218 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][20] ), .A1(\sa_events[1][20] ), .A2(\sa_events[2][20] ), .A3(\sa_events[3][20] ), .Z(n243));
Q_MX04 U219 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n243), .A1(n242), .A2(n241), .A3(n240), .Z(sa_mux1[20]));
Q_MX04 U220 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][21] ), .A1(\sa_events[13][21] ), .A2(\sa_events[14][21] ), .A3(\sa_events[15][21] ), .Z(n244));
Q_MX04 U221 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][21] ), .A1(\sa_events[9][21] ), .A2(\sa_events[10][21] ), .A3(\sa_events[11][21] ), .Z(n245));
Q_MX04 U222 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][21] ), .A1(\sa_events[5][21] ), .A2(\sa_events[6][21] ), .A3(\sa_events[7][21] ), .Z(n246));
Q_MX04 U223 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][21] ), .A1(\sa_events[1][21] ), .A2(\sa_events[2][21] ), .A3(\sa_events[3][21] ), .Z(n247));
Q_MX04 U224 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n247), .A1(n246), .A2(n245), .A3(n244), .Z(sa_mux1[21]));
Q_MX04 U225 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][22] ), .A1(\sa_events[13][22] ), .A2(\sa_events[14][22] ), .A3(\sa_events[15][22] ), .Z(n248));
Q_MX04 U226 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][22] ), .A1(\sa_events[9][22] ), .A2(\sa_events[10][22] ), .A3(\sa_events[11][22] ), .Z(n249));
Q_MX04 U227 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][22] ), .A1(\sa_events[5][22] ), .A2(\sa_events[6][22] ), .A3(\sa_events[7][22] ), .Z(n250));
Q_MX04 U228 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][22] ), .A1(\sa_events[1][22] ), .A2(\sa_events[2][22] ), .A3(\sa_events[3][22] ), .Z(n251));
Q_MX04 U229 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n251), .A1(n250), .A2(n249), .A3(n248), .Z(sa_mux1[22]));
Q_MX04 U230 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][23] ), .A1(\sa_events[13][23] ), .A2(\sa_events[14][23] ), .A3(\sa_events[15][23] ), .Z(n252));
Q_MX04 U231 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][23] ), .A1(\sa_events[9][23] ), .A2(\sa_events[10][23] ), .A3(\sa_events[11][23] ), .Z(n253));
Q_MX04 U232 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][23] ), .A1(\sa_events[5][23] ), .A2(\sa_events[6][23] ), .A3(\sa_events[7][23] ), .Z(n254));
Q_MX04 U233 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][23] ), .A1(\sa_events[1][23] ), .A2(\sa_events[2][23] ), .A3(\sa_events[3][23] ), .Z(n255));
Q_MX04 U234 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n255), .A1(n254), .A2(n253), .A3(n252), .Z(sa_mux1[23]));
Q_MX04 U235 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][24] ), .A1(\sa_events[13][24] ), .A2(\sa_events[14][24] ), .A3(\sa_events[15][24] ), .Z(n256));
Q_MX04 U236 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][24] ), .A1(\sa_events[9][24] ), .A2(\sa_events[10][24] ), .A3(\sa_events[11][24] ), .Z(n257));
Q_MX04 U237 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][24] ), .A1(\sa_events[5][24] ), .A2(\sa_events[6][24] ), .A3(\sa_events[7][24] ), .Z(n258));
Q_MX04 U238 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][24] ), .A1(\sa_events[1][24] ), .A2(\sa_events[2][24] ), .A3(\sa_events[3][24] ), .Z(n259));
Q_MX04 U239 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n259), .A1(n258), .A2(n257), .A3(n256), .Z(sa_mux1[24]));
Q_MX04 U240 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][25] ), .A1(\sa_events[13][25] ), .A2(\sa_events[14][25] ), .A3(\sa_events[15][25] ), .Z(n260));
Q_MX04 U241 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][25] ), .A1(\sa_events[9][25] ), .A2(\sa_events[10][25] ), .A3(\sa_events[11][25] ), .Z(n261));
Q_MX04 U242 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][25] ), .A1(\sa_events[5][25] ), .A2(\sa_events[6][25] ), .A3(\sa_events[7][25] ), .Z(n262));
Q_MX04 U243 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][25] ), .A1(\sa_events[1][25] ), .A2(\sa_events[2][25] ), .A3(\sa_events[3][25] ), .Z(n263));
Q_MX04 U244 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n263), .A1(n262), .A2(n261), .A3(n260), .Z(sa_mux1[25]));
Q_MX04 U245 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][26] ), .A1(\sa_events[13][26] ), .A2(\sa_events[14][26] ), .A3(\sa_events[15][26] ), .Z(n264));
Q_MX04 U246 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][26] ), .A1(\sa_events[9][26] ), .A2(\sa_events[10][26] ), .A3(\sa_events[11][26] ), .Z(n265));
Q_MX04 U247 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][26] ), .A1(\sa_events[5][26] ), .A2(\sa_events[6][26] ), .A3(\sa_events[7][26] ), .Z(n266));
Q_MX04 U248 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][26] ), .A1(\sa_events[1][26] ), .A2(\sa_events[2][26] ), .A3(\sa_events[3][26] ), .Z(n267));
Q_MX04 U249 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n267), .A1(n266), .A2(n265), .A3(n264), .Z(sa_mux1[26]));
Q_MX04 U250 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][27] ), .A1(\sa_events[13][27] ), .A2(\sa_events[14][27] ), .A3(\sa_events[15][27] ), .Z(n268));
Q_MX04 U251 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][27] ), .A1(\sa_events[9][27] ), .A2(\sa_events[10][27] ), .A3(\sa_events[11][27] ), .Z(n269));
Q_MX04 U252 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][27] ), .A1(\sa_events[5][27] ), .A2(\sa_events[6][27] ), .A3(\sa_events[7][27] ), .Z(n270));
Q_MX04 U253 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][27] ), .A1(\sa_events[1][27] ), .A2(\sa_events[2][27] ), .A3(\sa_events[3][27] ), .Z(n271));
Q_MX04 U254 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n271), .A1(n270), .A2(n269), .A3(n268), .Z(sa_mux1[27]));
Q_MX04 U255 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][28] ), .A1(\sa_events[13][28] ), .A2(\sa_events[14][28] ), .A3(\sa_events[15][28] ), .Z(n272));
Q_MX04 U256 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][28] ), .A1(\sa_events[9][28] ), .A2(\sa_events[10][28] ), .A3(\sa_events[11][28] ), .Z(n273));
Q_MX04 U257 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][28] ), .A1(\sa_events[5][28] ), .A2(\sa_events[6][28] ), .A3(\sa_events[7][28] ), .Z(n274));
Q_MX04 U258 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][28] ), .A1(\sa_events[1][28] ), .A2(\sa_events[2][28] ), .A3(\sa_events[3][28] ), .Z(n275));
Q_MX04 U259 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n275), .A1(n274), .A2(n273), .A3(n272), .Z(sa_mux1[28]));
Q_MX04 U260 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][29] ), .A1(\sa_events[13][29] ), .A2(\sa_events[14][29] ), .A3(\sa_events[15][29] ), .Z(n276));
Q_MX04 U261 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][29] ), .A1(\sa_events[9][29] ), .A2(\sa_events[10][29] ), .A3(\sa_events[11][29] ), .Z(n277));
Q_MX04 U262 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][29] ), .A1(\sa_events[5][29] ), .A2(\sa_events[6][29] ), .A3(\sa_events[7][29] ), .Z(n278));
Q_MX04 U263 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][29] ), .A1(\sa_events[1][29] ), .A2(\sa_events[2][29] ), .A3(\sa_events[3][29] ), .Z(n279));
Q_MX04 U264 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n279), .A1(n278), .A2(n277), .A3(n276), .Z(sa_mux1[29]));
Q_MX04 U265 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][30] ), .A1(\sa_events[13][30] ), .A2(\sa_events[14][30] ), .A3(\sa_events[15][30] ), .Z(n280));
Q_MX04 U266 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][30] ), .A1(\sa_events[9][30] ), .A2(\sa_events[10][30] ), .A3(\sa_events[11][30] ), .Z(n281));
Q_MX04 U267 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][30] ), .A1(\sa_events[5][30] ), .A2(\sa_events[6][30] ), .A3(\sa_events[7][30] ), .Z(n282));
Q_MX04 U268 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][30] ), .A1(\sa_events[1][30] ), .A2(\sa_events[2][30] ), .A3(\sa_events[3][30] ), .Z(n283));
Q_MX04 U269 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n283), .A1(n282), .A2(n281), .A3(n280), .Z(sa_mux1[30]));
Q_MX04 U270 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][31] ), .A1(\sa_events[13][31] ), .A2(\sa_events[14][31] ), .A3(\sa_events[15][31] ), .Z(n284));
Q_MX04 U271 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][31] ), .A1(\sa_events[9][31] ), .A2(\sa_events[10][31] ), .A3(\sa_events[11][31] ), .Z(n285));
Q_MX04 U272 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][31] ), .A1(\sa_events[5][31] ), .A2(\sa_events[6][31] ), .A3(\sa_events[7][31] ), .Z(n286));
Q_MX04 U273 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][31] ), .A1(\sa_events[1][31] ), .A2(\sa_events[2][31] ), .A3(\sa_events[3][31] ), .Z(n287));
Q_MX04 U274 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n287), .A1(n286), .A2(n285), .A3(n284), .Z(sa_mux1[31]));
Q_MX04 U275 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][32] ), .A1(\sa_events[13][32] ), .A2(\sa_events[14][32] ), .A3(\sa_events[15][32] ), .Z(n288));
Q_MX04 U276 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][32] ), .A1(\sa_events[9][32] ), .A2(\sa_events[10][32] ), .A3(\sa_events[11][32] ), .Z(n289));
Q_MX04 U277 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][32] ), .A1(\sa_events[5][32] ), .A2(\sa_events[6][32] ), .A3(\sa_events[7][32] ), .Z(n290));
Q_MX04 U278 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][32] ), .A1(\sa_events[1][32] ), .A2(\sa_events[2][32] ), .A3(\sa_events[3][32] ), .Z(n291));
Q_MX04 U279 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n291), .A1(n290), .A2(n289), .A3(n288), .Z(sa_mux1[32]));
Q_MX04 U280 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][33] ), .A1(\sa_events[13][33] ), .A2(\sa_events[14][33] ), .A3(\sa_events[15][33] ), .Z(n292));
Q_MX04 U281 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][33] ), .A1(\sa_events[9][33] ), .A2(\sa_events[10][33] ), .A3(\sa_events[11][33] ), .Z(n293));
Q_MX04 U282 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][33] ), .A1(\sa_events[5][33] ), .A2(\sa_events[6][33] ), .A3(\sa_events[7][33] ), .Z(n294));
Q_MX04 U283 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][33] ), .A1(\sa_events[1][33] ), .A2(\sa_events[2][33] ), .A3(\sa_events[3][33] ), .Z(n295));
Q_MX04 U284 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n295), .A1(n294), .A2(n293), .A3(n292), .Z(sa_mux1[33]));
Q_MX04 U285 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][34] ), .A1(\sa_events[13][34] ), .A2(\sa_events[14][34] ), .A3(\sa_events[15][34] ), .Z(n296));
Q_MX04 U286 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][34] ), .A1(\sa_events[9][34] ), .A2(\sa_events[10][34] ), .A3(\sa_events[11][34] ), .Z(n297));
Q_MX04 U287 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][34] ), .A1(\sa_events[5][34] ), .A2(\sa_events[6][34] ), .A3(\sa_events[7][34] ), .Z(n298));
Q_MX04 U288 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][34] ), .A1(\sa_events[1][34] ), .A2(\sa_events[2][34] ), .A3(\sa_events[3][34] ), .Z(n299));
Q_MX04 U289 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n299), .A1(n298), .A2(n297), .A3(n296), .Z(sa_mux1[34]));
Q_MX04 U290 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][35] ), .A1(\sa_events[13][35] ), .A2(\sa_events[14][35] ), .A3(\sa_events[15][35] ), .Z(n300));
Q_MX04 U291 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][35] ), .A1(\sa_events[9][35] ), .A2(\sa_events[10][35] ), .A3(\sa_events[11][35] ), .Z(n301));
Q_MX04 U292 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][35] ), .A1(\sa_events[5][35] ), .A2(\sa_events[6][35] ), .A3(\sa_events[7][35] ), .Z(n302));
Q_MX04 U293 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][35] ), .A1(\sa_events[1][35] ), .A2(\sa_events[2][35] ), .A3(\sa_events[3][35] ), .Z(n303));
Q_MX04 U294 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n303), .A1(n302), .A2(n301), .A3(n300), .Z(sa_mux1[35]));
Q_MX04 U295 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][36] ), .A1(\sa_events[13][36] ), .A2(\sa_events[14][36] ), .A3(\sa_events[15][36] ), .Z(n304));
Q_MX04 U296 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][36] ), .A1(\sa_events[9][36] ), .A2(\sa_events[10][36] ), .A3(\sa_events[11][36] ), .Z(n305));
Q_MX04 U297 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][36] ), .A1(\sa_events[5][36] ), .A2(\sa_events[6][36] ), .A3(\sa_events[7][36] ), .Z(n306));
Q_MX04 U298 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][36] ), .A1(\sa_events[1][36] ), .A2(\sa_events[2][36] ), .A3(\sa_events[3][36] ), .Z(n307));
Q_MX04 U299 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n307), .A1(n306), .A2(n305), .A3(n304), .Z(sa_mux1[36]));
Q_MX04 U300 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][37] ), .A1(\sa_events[13][37] ), .A2(\sa_events[14][37] ), .A3(\sa_events[15][37] ), .Z(n308));
Q_MX04 U301 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][37] ), .A1(\sa_events[9][37] ), .A2(\sa_events[10][37] ), .A3(\sa_events[11][37] ), .Z(n309));
Q_MX04 U302 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][37] ), .A1(\sa_events[5][37] ), .A2(\sa_events[6][37] ), .A3(\sa_events[7][37] ), .Z(n310));
Q_MX04 U303 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][37] ), .A1(\sa_events[1][37] ), .A2(\sa_events[2][37] ), .A3(\sa_events[3][37] ), .Z(n311));
Q_MX04 U304 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n311), .A1(n310), .A2(n309), .A3(n308), .Z(sa_mux1[37]));
Q_MX04 U305 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][38] ), .A1(\sa_events[13][38] ), .A2(\sa_events[14][38] ), .A3(\sa_events[15][38] ), .Z(n312));
Q_MX04 U306 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][38] ), .A1(\sa_events[9][38] ), .A2(\sa_events[10][38] ), .A3(\sa_events[11][38] ), .Z(n313));
Q_MX04 U307 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][38] ), .A1(\sa_events[5][38] ), .A2(\sa_events[6][38] ), .A3(\sa_events[7][38] ), .Z(n314));
Q_MX04 U308 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][38] ), .A1(\sa_events[1][38] ), .A2(\sa_events[2][38] ), .A3(\sa_events[3][38] ), .Z(n315));
Q_MX04 U309 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n315), .A1(n314), .A2(n313), .A3(n312), .Z(sa_mux1[38]));
Q_MX04 U310 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][39] ), .A1(\sa_events[13][39] ), .A2(\sa_events[14][39] ), .A3(\sa_events[15][39] ), .Z(n316));
Q_MX04 U311 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][39] ), .A1(\sa_events[9][39] ), .A2(\sa_events[10][39] ), .A3(\sa_events[11][39] ), .Z(n317));
Q_MX04 U312 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][39] ), .A1(\sa_events[5][39] ), .A2(\sa_events[6][39] ), .A3(\sa_events[7][39] ), .Z(n318));
Q_MX04 U313 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][39] ), .A1(\sa_events[1][39] ), .A2(\sa_events[2][39] ), .A3(\sa_events[3][39] ), .Z(n319));
Q_MX04 U314 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n319), .A1(n318), .A2(n317), .A3(n316), .Z(sa_mux1[39]));
Q_MX04 U315 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][40] ), .A1(\sa_events[13][40] ), .A2(\sa_events[14][40] ), .A3(\sa_events[15][40] ), .Z(n320));
Q_MX04 U316 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][40] ), .A1(\sa_events[9][40] ), .A2(\sa_events[10][40] ), .A3(\sa_events[11][40] ), .Z(n321));
Q_MX04 U317 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][40] ), .A1(\sa_events[5][40] ), .A2(\sa_events[6][40] ), .A3(\sa_events[7][40] ), .Z(n322));
Q_MX04 U318 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][40] ), .A1(\sa_events[1][40] ), .A2(\sa_events[2][40] ), .A3(\sa_events[3][40] ), .Z(n323));
Q_MX04 U319 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n323), .A1(n322), .A2(n321), .A3(n320), .Z(sa_mux1[40]));
Q_MX04 U320 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][41] ), .A1(\sa_events[13][41] ), .A2(\sa_events[14][41] ), .A3(\sa_events[15][41] ), .Z(n324));
Q_MX04 U321 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][41] ), .A1(\sa_events[9][41] ), .A2(\sa_events[10][41] ), .A3(\sa_events[11][41] ), .Z(n325));
Q_MX04 U322 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][41] ), .A1(\sa_events[5][41] ), .A2(\sa_events[6][41] ), .A3(\sa_events[7][41] ), .Z(n326));
Q_MX04 U323 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][41] ), .A1(\sa_events[1][41] ), .A2(\sa_events[2][41] ), .A3(\sa_events[3][41] ), .Z(n327));
Q_MX04 U324 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n327), .A1(n326), .A2(n325), .A3(n324), .Z(sa_mux1[41]));
Q_MX04 U325 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][42] ), .A1(\sa_events[13][42] ), .A2(\sa_events[14][42] ), .A3(\sa_events[15][42] ), .Z(n328));
Q_MX04 U326 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][42] ), .A1(\sa_events[9][42] ), .A2(\sa_events[10][42] ), .A3(\sa_events[11][42] ), .Z(n329));
Q_MX04 U327 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][42] ), .A1(\sa_events[5][42] ), .A2(\sa_events[6][42] ), .A3(\sa_events[7][42] ), .Z(n330));
Q_MX04 U328 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][42] ), .A1(\sa_events[1][42] ), .A2(\sa_events[2][42] ), .A3(\sa_events[3][42] ), .Z(n331));
Q_MX04 U329 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n331), .A1(n330), .A2(n329), .A3(n328), .Z(sa_mux1[42]));
Q_MX04 U330 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][43] ), .A1(\sa_events[13][43] ), .A2(\sa_events[14][43] ), .A3(\sa_events[15][43] ), .Z(n332));
Q_MX04 U331 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][43] ), .A1(\sa_events[9][43] ), .A2(\sa_events[10][43] ), .A3(\sa_events[11][43] ), .Z(n333));
Q_MX04 U332 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][43] ), .A1(\sa_events[5][43] ), .A2(\sa_events[6][43] ), .A3(\sa_events[7][43] ), .Z(n334));
Q_MX04 U333 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][43] ), .A1(\sa_events[1][43] ), .A2(\sa_events[2][43] ), .A3(\sa_events[3][43] ), .Z(n335));
Q_MX04 U334 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n335), .A1(n334), .A2(n333), .A3(n332), .Z(sa_mux1[43]));
Q_MX04 U335 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][44] ), .A1(\sa_events[13][44] ), .A2(\sa_events[14][44] ), .A3(\sa_events[15][44] ), .Z(n336));
Q_MX04 U336 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][44] ), .A1(\sa_events[9][44] ), .A2(\sa_events[10][44] ), .A3(\sa_events[11][44] ), .Z(n337));
Q_MX04 U337 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][44] ), .A1(\sa_events[5][44] ), .A2(\sa_events[6][44] ), .A3(\sa_events[7][44] ), .Z(n338));
Q_MX04 U338 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][44] ), .A1(\sa_events[1][44] ), .A2(\sa_events[2][44] ), .A3(\sa_events[3][44] ), .Z(n339));
Q_MX04 U339 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n339), .A1(n338), .A2(n337), .A3(n336), .Z(sa_mux1[44]));
Q_MX04 U340 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][45] ), .A1(\sa_events[13][45] ), .A2(\sa_events[14][45] ), .A3(\sa_events[15][45] ), .Z(n340));
Q_MX04 U341 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][45] ), .A1(\sa_events[9][45] ), .A2(\sa_events[10][45] ), .A3(\sa_events[11][45] ), .Z(n341));
Q_MX04 U342 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][45] ), .A1(\sa_events[5][45] ), .A2(\sa_events[6][45] ), .A3(\sa_events[7][45] ), .Z(n342));
Q_MX04 U343 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][45] ), .A1(\sa_events[1][45] ), .A2(\sa_events[2][45] ), .A3(\sa_events[3][45] ), .Z(n343));
Q_MX04 U344 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n343), .A1(n342), .A2(n341), .A3(n340), .Z(sa_mux1[45]));
Q_MX04 U345 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][46] ), .A1(\sa_events[13][46] ), .A2(\sa_events[14][46] ), .A3(\sa_events[15][46] ), .Z(n344));
Q_MX04 U346 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][46] ), .A1(\sa_events[9][46] ), .A2(\sa_events[10][46] ), .A3(\sa_events[11][46] ), .Z(n345));
Q_MX04 U347 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][46] ), .A1(\sa_events[5][46] ), .A2(\sa_events[6][46] ), .A3(\sa_events[7][46] ), .Z(n346));
Q_MX04 U348 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][46] ), .A1(\sa_events[1][46] ), .A2(\sa_events[2][46] ), .A3(\sa_events[3][46] ), .Z(n347));
Q_MX04 U349 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n347), .A1(n346), .A2(n345), .A3(n344), .Z(sa_mux1[46]));
Q_MX04 U350 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][47] ), .A1(\sa_events[13][47] ), .A2(\sa_events[14][47] ), .A3(\sa_events[15][47] ), .Z(n348));
Q_MX04 U351 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][47] ), .A1(\sa_events[9][47] ), .A2(\sa_events[10][47] ), .A3(\sa_events[11][47] ), .Z(n349));
Q_MX04 U352 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][47] ), .A1(\sa_events[5][47] ), .A2(\sa_events[6][47] ), .A3(\sa_events[7][47] ), .Z(n350));
Q_MX04 U353 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][47] ), .A1(\sa_events[1][47] ), .A2(\sa_events[2][47] ), .A3(\sa_events[3][47] ), .Z(n351));
Q_MX04 U354 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n351), .A1(n350), .A2(n349), .A3(n348), .Z(sa_mux1[47]));
Q_MX04 U355 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][48] ), .A1(\sa_events[13][48] ), .A2(\sa_events[14][48] ), .A3(\sa_events[15][48] ), .Z(n352));
Q_MX04 U356 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][48] ), .A1(\sa_events[9][48] ), .A2(\sa_events[10][48] ), .A3(\sa_events[11][48] ), .Z(n353));
Q_MX04 U357 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][48] ), .A1(\sa_events[5][48] ), .A2(\sa_events[6][48] ), .A3(\sa_events[7][48] ), .Z(n354));
Q_MX04 U358 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][48] ), .A1(\sa_events[1][48] ), .A2(\sa_events[2][48] ), .A3(\sa_events[3][48] ), .Z(n355));
Q_MX04 U359 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n355), .A1(n354), .A2(n353), .A3(n352), .Z(sa_mux1[48]));
Q_MX04 U360 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][49] ), .A1(\sa_events[13][49] ), .A2(\sa_events[14][49] ), .A3(\sa_events[15][49] ), .Z(n356));
Q_MX04 U361 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][49] ), .A1(\sa_events[9][49] ), .A2(\sa_events[10][49] ), .A3(\sa_events[11][49] ), .Z(n357));
Q_MX04 U362 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][49] ), .A1(\sa_events[5][49] ), .A2(\sa_events[6][49] ), .A3(\sa_events[7][49] ), .Z(n358));
Q_MX04 U363 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][49] ), .A1(\sa_events[1][49] ), .A2(\sa_events[2][49] ), .A3(\sa_events[3][49] ), .Z(n359));
Q_MX04 U364 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n359), .A1(n358), .A2(n357), .A3(n356), .Z(sa_mux1[49]));
Q_MX04 U365 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][50] ), .A1(\sa_events[13][50] ), .A2(\sa_events[14][50] ), .A3(\sa_events[15][50] ), .Z(n360));
Q_MX04 U366 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][50] ), .A1(\sa_events[9][50] ), .A2(\sa_events[10][50] ), .A3(\sa_events[11][50] ), .Z(n361));
Q_MX04 U367 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][50] ), .A1(\sa_events[5][50] ), .A2(\sa_events[6][50] ), .A3(\sa_events[7][50] ), .Z(n362));
Q_MX04 U368 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][50] ), .A1(\sa_events[1][50] ), .A2(\sa_events[2][50] ), .A3(\sa_events[3][50] ), .Z(n363));
Q_MX04 U369 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n363), .A1(n362), .A2(n361), .A3(n360), .Z(sa_mux1[50]));
Q_MX04 U370 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][51] ), .A1(\sa_events[13][51] ), .A2(\sa_events[14][51] ), .A3(\sa_events[15][51] ), .Z(n364));
Q_MX04 U371 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][51] ), .A1(\sa_events[9][51] ), .A2(\sa_events[10][51] ), .A3(\sa_events[11][51] ), .Z(n365));
Q_MX04 U372 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][51] ), .A1(\sa_events[5][51] ), .A2(\sa_events[6][51] ), .A3(\sa_events[7][51] ), .Z(n366));
Q_MX04 U373 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][51] ), .A1(\sa_events[1][51] ), .A2(\sa_events[2][51] ), .A3(\sa_events[3][51] ), .Z(n367));
Q_MX04 U374 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n367), .A1(n366), .A2(n365), .A3(n364), .Z(sa_mux1[51]));
Q_MX04 U375 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][52] ), .A1(\sa_events[13][52] ), .A2(\sa_events[14][52] ), .A3(\sa_events[15][52] ), .Z(n368));
Q_MX04 U376 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][52] ), .A1(\sa_events[9][52] ), .A2(\sa_events[10][52] ), .A3(\sa_events[11][52] ), .Z(n369));
Q_MX04 U377 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][52] ), .A1(\sa_events[5][52] ), .A2(\sa_events[6][52] ), .A3(\sa_events[7][52] ), .Z(n370));
Q_MX04 U378 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][52] ), .A1(\sa_events[1][52] ), .A2(\sa_events[2][52] ), .A3(\sa_events[3][52] ), .Z(n371));
Q_MX04 U379 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n371), .A1(n370), .A2(n369), .A3(n368), .Z(sa_mux1[52]));
Q_MX04 U380 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][53] ), .A1(\sa_events[13][53] ), .A2(\sa_events[14][53] ), .A3(\sa_events[15][53] ), .Z(n372));
Q_MX04 U381 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][53] ), .A1(\sa_events[9][53] ), .A2(\sa_events[10][53] ), .A3(\sa_events[11][53] ), .Z(n373));
Q_MX04 U382 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][53] ), .A1(\sa_events[5][53] ), .A2(\sa_events[6][53] ), .A3(\sa_events[7][53] ), .Z(n374));
Q_MX04 U383 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][53] ), .A1(\sa_events[1][53] ), .A2(\sa_events[2][53] ), .A3(\sa_events[3][53] ), .Z(n375));
Q_MX04 U384 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n375), .A1(n374), .A2(n373), .A3(n372), .Z(sa_mux1[53]));
Q_MX04 U385 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][54] ), .A1(\sa_events[13][54] ), .A2(\sa_events[14][54] ), .A3(\sa_events[15][54] ), .Z(n376));
Q_MX04 U386 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][54] ), .A1(\sa_events[9][54] ), .A2(\sa_events[10][54] ), .A3(\sa_events[11][54] ), .Z(n377));
Q_MX04 U387 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][54] ), .A1(\sa_events[5][54] ), .A2(\sa_events[6][54] ), .A3(\sa_events[7][54] ), .Z(n378));
Q_MX04 U388 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][54] ), .A1(\sa_events[1][54] ), .A2(\sa_events[2][54] ), .A3(\sa_events[3][54] ), .Z(n379));
Q_MX04 U389 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n379), .A1(n378), .A2(n377), .A3(n376), .Z(sa_mux1[54]));
Q_MX04 U390 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][55] ), .A1(\sa_events[13][55] ), .A2(\sa_events[14][55] ), .A3(\sa_events[15][55] ), .Z(n380));
Q_MX04 U391 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][55] ), .A1(\sa_events[9][55] ), .A2(\sa_events[10][55] ), .A3(\sa_events[11][55] ), .Z(n381));
Q_MX04 U392 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][55] ), .A1(\sa_events[5][55] ), .A2(\sa_events[6][55] ), .A3(\sa_events[7][55] ), .Z(n382));
Q_MX04 U393 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][55] ), .A1(\sa_events[1][55] ), .A2(\sa_events[2][55] ), .A3(\sa_events[3][55] ), .Z(n383));
Q_MX04 U394 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n383), .A1(n382), .A2(n381), .A3(n380), .Z(sa_mux1[55]));
Q_MX04 U395 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][56] ), .A1(\sa_events[13][56] ), .A2(\sa_events[14][56] ), .A3(\sa_events[15][56] ), .Z(n384));
Q_MX04 U396 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][56] ), .A1(\sa_events[9][56] ), .A2(\sa_events[10][56] ), .A3(\sa_events[11][56] ), .Z(n385));
Q_MX04 U397 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][56] ), .A1(\sa_events[5][56] ), .A2(\sa_events[6][56] ), .A3(\sa_events[7][56] ), .Z(n386));
Q_MX04 U398 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][56] ), .A1(\sa_events[1][56] ), .A2(\sa_events[2][56] ), .A3(\sa_events[3][56] ), .Z(n387));
Q_MX04 U399 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n387), .A1(n386), .A2(n385), .A3(n384), .Z(sa_mux1[56]));
Q_MX04 U400 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][57] ), .A1(\sa_events[13][57] ), .A2(\sa_events[14][57] ), .A3(\sa_events[15][57] ), .Z(n388));
Q_MX04 U401 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][57] ), .A1(\sa_events[9][57] ), .A2(\sa_events[10][57] ), .A3(\sa_events[11][57] ), .Z(n389));
Q_MX04 U402 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][57] ), .A1(\sa_events[5][57] ), .A2(\sa_events[6][57] ), .A3(\sa_events[7][57] ), .Z(n390));
Q_MX04 U403 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][57] ), .A1(\sa_events[1][57] ), .A2(\sa_events[2][57] ), .A3(\sa_events[3][57] ), .Z(n391));
Q_MX04 U404 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n391), .A1(n390), .A2(n389), .A3(n388), .Z(sa_mux1[57]));
Q_MX04 U405 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][58] ), .A1(\sa_events[13][58] ), .A2(\sa_events[14][58] ), .A3(\sa_events[15][58] ), .Z(n392));
Q_MX04 U406 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][58] ), .A1(\sa_events[9][58] ), .A2(\sa_events[10][58] ), .A3(\sa_events[11][58] ), .Z(n393));
Q_MX04 U407 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][58] ), .A1(\sa_events[5][58] ), .A2(\sa_events[6][58] ), .A3(\sa_events[7][58] ), .Z(n394));
Q_MX04 U408 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][58] ), .A1(\sa_events[1][58] ), .A2(\sa_events[2][58] ), .A3(\sa_events[3][58] ), .Z(n395));
Q_MX04 U409 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n395), .A1(n394), .A2(n393), .A3(n392), .Z(sa_mux1[58]));
Q_MX04 U410 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][59] ), .A1(\sa_events[13][59] ), .A2(\sa_events[14][59] ), .A3(\sa_events[15][59] ), .Z(n396));
Q_MX04 U411 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][59] ), .A1(\sa_events[9][59] ), .A2(\sa_events[10][59] ), .A3(\sa_events[11][59] ), .Z(n397));
Q_MX04 U412 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][59] ), .A1(\sa_events[5][59] ), .A2(\sa_events[6][59] ), .A3(\sa_events[7][59] ), .Z(n398));
Q_MX04 U413 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][59] ), .A1(\sa_events[1][59] ), .A2(\sa_events[2][59] ), .A3(\sa_events[3][59] ), .Z(n399));
Q_MX04 U414 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n399), .A1(n398), .A2(n397), .A3(n396), .Z(sa_mux1[59]));
Q_MX04 U415 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][60] ), .A1(\sa_events[13][60] ), .A2(\sa_events[14][60] ), .A3(\sa_events[15][60] ), .Z(n400));
Q_MX04 U416 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][60] ), .A1(\sa_events[9][60] ), .A2(\sa_events[10][60] ), .A3(\sa_events[11][60] ), .Z(n401));
Q_MX04 U417 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][60] ), .A1(\sa_events[5][60] ), .A2(\sa_events[6][60] ), .A3(\sa_events[7][60] ), .Z(n402));
Q_MX04 U418 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][60] ), .A1(\sa_events[1][60] ), .A2(\sa_events[2][60] ), .A3(\sa_events[3][60] ), .Z(n403));
Q_MX04 U419 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n403), .A1(n402), .A2(n401), .A3(n400), .Z(sa_mux1[60]));
Q_MX04 U420 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][61] ), .A1(\sa_events[13][61] ), .A2(\sa_events[14][61] ), .A3(\sa_events[15][61] ), .Z(n404));
Q_MX04 U421 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][61] ), .A1(\sa_events[9][61] ), .A2(\sa_events[10][61] ), .A3(\sa_events[11][61] ), .Z(n405));
Q_MX04 U422 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][61] ), .A1(\sa_events[5][61] ), .A2(\sa_events[6][61] ), .A3(\sa_events[7][61] ), .Z(n406));
Q_MX04 U423 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][61] ), .A1(\sa_events[1][61] ), .A2(\sa_events[2][61] ), .A3(\sa_events[3][61] ), .Z(n407));
Q_MX04 U424 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n407), .A1(n406), .A2(n405), .A3(n404), .Z(sa_mux1[61]));
Q_MX04 U425 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][62] ), .A1(\sa_events[13][62] ), .A2(\sa_events[14][62] ), .A3(\sa_events[15][62] ), .Z(n408));
Q_MX04 U426 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][62] ), .A1(\sa_events[9][62] ), .A2(\sa_events[10][62] ), .A3(\sa_events[11][62] ), .Z(n409));
Q_MX04 U427 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][62] ), .A1(\sa_events[5][62] ), .A2(\sa_events[6][62] ), .A3(\sa_events[7][62] ), .Z(n410));
Q_MX04 U428 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][62] ), .A1(\sa_events[1][62] ), .A2(\sa_events[2][62] ), .A3(\sa_events[3][62] ), .Z(n411));
Q_MX04 U429 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n411), .A1(n410), .A2(n409), .A3(n408), .Z(sa_mux1[62]));
Q_MX04 U430 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[12][63] ), .A1(\sa_events[13][63] ), .A2(\sa_events[14][63] ), .A3(\sa_events[15][63] ), .Z(n412));
Q_MX04 U431 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[8][63] ), .A1(\sa_events[9][63] ), .A2(\sa_events[10][63] ), .A3(\sa_events[11][63] ), .Z(n413));
Q_MX04 U432 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[4][63] ), .A1(\sa_events[5][63] ), .A2(\sa_events[6][63] ), .A3(\sa_events[7][63] ), .Z(n414));
Q_MX04 U433 ( .S0(sa_event_sel[6]), .S1(sa_event_sel[7]), .A0(\sa_events[0][63] ), .A1(\sa_events[1][63] ), .A2(\sa_events[2][63] ), .A3(\sa_events[3][63] ), .Z(n415));
Q_MX04 U434 ( .S0(sa_event_sel[8]), .S1(sa_event_sel[9]), .A0(n415), .A1(n414), .A2(n413), .A3(n412), .Z(sa_mux1[63]));
Q_FDP4EP \sa_count_REG[0] ( .CK(clk), .CE(n159), .R(n416), .D(n107), .Q(sa_count[0]));
Q_INV U436 ( .A(rst_n), .Z(n416));
Q_FDP4EP \sa_count_REG[1] ( .CK(clk), .CE(n159), .R(n416), .D(n108), .Q(sa_count[1]));
Q_FDP4EP \sa_count_REG[2] ( .CK(clk), .CE(n159), .R(n416), .D(n109), .Q(sa_count[2]));
Q_FDP4EP \sa_count_REG[3] ( .CK(clk), .CE(n159), .R(n416), .D(n110), .Q(sa_count[3]));
Q_FDP4EP \sa_count_REG[4] ( .CK(clk), .CE(n159), .R(n416), .D(n111), .Q(sa_count[4]));
Q_FDP4EP \sa_count_REG[5] ( .CK(clk), .CE(n159), .R(n416), .D(n112), .Q(sa_count[5]));
Q_FDP4EP \sa_count_REG[6] ( .CK(clk), .CE(n159), .R(n416), .D(n113), .Q(sa_count[6]));
Q_FDP4EP \sa_count_REG[7] ( .CK(clk), .CE(n159), .R(n416), .D(n114), .Q(sa_count[7]));
Q_FDP4EP \sa_count_REG[8] ( .CK(clk), .CE(n159), .R(n416), .D(n115), .Q(sa_count[8]));
Q_FDP4EP \sa_count_REG[9] ( .CK(clk), .CE(n159), .R(n416), .D(n116), .Q(sa_count[9]));
Q_FDP4EP \sa_count_REG[10] ( .CK(clk), .CE(n159), .R(n416), .D(n117), .Q(sa_count[10]));
Q_FDP4EP \sa_count_REG[11] ( .CK(clk), .CE(n159), .R(n416), .D(n118), .Q(sa_count[11]));
Q_FDP4EP \sa_count_REG[12] ( .CK(clk), .CE(n159), .R(n416), .D(n119), .Q(sa_count[12]));
Q_FDP4EP \sa_count_REG[13] ( .CK(clk), .CE(n159), .R(n416), .D(n120), .Q(sa_count[13]));
Q_FDP4EP \sa_count_REG[14] ( .CK(clk), .CE(n159), .R(n416), .D(n121), .Q(sa_count[14]));
Q_FDP4EP \sa_count_REG[15] ( .CK(clk), .CE(n159), .R(n416), .D(n122), .Q(sa_count[15]));
Q_FDP4EP \sa_count_REG[16] ( .CK(clk), .CE(n159), .R(n416), .D(n123), .Q(sa_count[16]));
Q_FDP4EP \sa_count_REG[17] ( .CK(clk), .CE(n159), .R(n416), .D(n124), .Q(sa_count[17]));
Q_FDP4EP \sa_count_REG[18] ( .CK(clk), .CE(n159), .R(n416), .D(n125), .Q(sa_count[18]));
Q_FDP4EP \sa_count_REG[19] ( .CK(clk), .CE(n159), .R(n416), .D(n126), .Q(sa_count[19]));
Q_FDP4EP \sa_count_REG[20] ( .CK(clk), .CE(n159), .R(n416), .D(n127), .Q(sa_count[20]));
Q_FDP4EP \sa_count_REG[21] ( .CK(clk), .CE(n159), .R(n416), .D(n128), .Q(sa_count[21]));
Q_FDP4EP \sa_count_REG[22] ( .CK(clk), .CE(n159), .R(n416), .D(n129), .Q(sa_count[22]));
Q_FDP4EP \sa_count_REG[23] ( .CK(clk), .CE(n159), .R(n416), .D(n130), .Q(sa_count[23]));
Q_FDP4EP \sa_count_REG[24] ( .CK(clk), .CE(n159), .R(n416), .D(n131), .Q(sa_count[24]));
Q_FDP4EP \sa_count_REG[25] ( .CK(clk), .CE(n159), .R(n416), .D(n132), .Q(sa_count[25]));
Q_FDP4EP \sa_count_REG[26] ( .CK(clk), .CE(n159), .R(n416), .D(n133), .Q(sa_count[26]));
Q_FDP4EP \sa_count_REG[27] ( .CK(clk), .CE(n159), .R(n416), .D(n134), .Q(sa_count[27]));
Q_FDP4EP \sa_count_REG[28] ( .CK(clk), .CE(n159), .R(n416), .D(n135), .Q(sa_count[28]));
Q_FDP4EP \sa_count_REG[29] ( .CK(clk), .CE(n159), .R(n416), .D(n136), .Q(sa_count[29]));
Q_FDP4EP \sa_count_REG[30] ( .CK(clk), .CE(n159), .R(n416), .D(n137), .Q(sa_count[30]));
Q_FDP4EP \sa_count_REG[31] ( .CK(clk), .CE(n159), .R(n416), .D(n138), .Q(sa_count[31]));
Q_FDP4EP \sa_count_REG[32] ( .CK(clk), .CE(n159), .R(n416), .D(n139), .Q(sa_count[32]));
Q_FDP4EP \sa_count_REG[33] ( .CK(clk), .CE(n159), .R(n416), .D(n140), .Q(sa_count[33]));
Q_FDP4EP \sa_count_REG[34] ( .CK(clk), .CE(n159), .R(n416), .D(n141), .Q(sa_count[34]));
Q_FDP4EP \sa_count_REG[35] ( .CK(clk), .CE(n159), .R(n416), .D(n142), .Q(sa_count[35]));
Q_FDP4EP \sa_count_REG[36] ( .CK(clk), .CE(n159), .R(n416), .D(n143), .Q(sa_count[36]));
Q_FDP4EP \sa_count_REG[37] ( .CK(clk), .CE(n159), .R(n416), .D(n144), .Q(sa_count[37]));
Q_FDP4EP \sa_count_REG[38] ( .CK(clk), .CE(n159), .R(n416), .D(n145), .Q(sa_count[38]));
Q_FDP4EP \sa_count_REG[39] ( .CK(clk), .CE(n159), .R(n416), .D(n146), .Q(sa_count[39]));
Q_FDP4EP \sa_count_REG[40] ( .CK(clk), .CE(n159), .R(n416), .D(n147), .Q(sa_count[40]));
Q_FDP4EP \sa_count_REG[41] ( .CK(clk), .CE(n159), .R(n416), .D(n148), .Q(sa_count[41]));
Q_FDP4EP \sa_count_REG[42] ( .CK(clk), .CE(n159), .R(n416), .D(n149), .Q(sa_count[42]));
Q_FDP4EP \sa_count_REG[43] ( .CK(clk), .CE(n159), .R(n416), .D(n150), .Q(sa_count[43]));
Q_FDP4EP \sa_count_REG[44] ( .CK(clk), .CE(n159), .R(n416), .D(n151), .Q(sa_count[44]));
Q_FDP4EP \sa_count_REG[45] ( .CK(clk), .CE(n159), .R(n416), .D(n152), .Q(sa_count[45]));
Q_FDP4EP \sa_count_REG[46] ( .CK(clk), .CE(n159), .R(n416), .D(n153), .Q(sa_count[46]));
Q_FDP4EP \sa_count_REG[47] ( .CK(clk), .CE(n159), .R(n416), .D(n154), .Q(sa_count[47]));
Q_FDP4EP \sa_count_REG[48] ( .CK(clk), .CE(n159), .R(n416), .D(n155), .Q(sa_count[48]));
Q_FDP4EP \sa_count_REG[49] ( .CK(clk), .CE(n159), .R(n416), .D(n156), .Q(sa_count[49]));
Q_FDP4EP \sa_snapshot_REG[0] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[0]), .Q(sa_snapshot[0]));
Q_FDP4EP \sa_snapshot_REG[1] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[1]), .Q(sa_snapshot[1]));
Q_FDP4EP \sa_snapshot_REG[2] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[2]), .Q(sa_snapshot[2]));
Q_FDP4EP \sa_snapshot_REG[3] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[3]), .Q(sa_snapshot[3]));
Q_FDP4EP \sa_snapshot_REG[4] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[4]), .Q(sa_snapshot[4]));
Q_FDP4EP \sa_snapshot_REG[5] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[5]), .Q(sa_snapshot[5]));
Q_FDP4EP \sa_snapshot_REG[6] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[6]), .Q(sa_snapshot[6]));
Q_FDP4EP \sa_snapshot_REG[7] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[7]), .Q(sa_snapshot[7]));
Q_FDP4EP \sa_snapshot_REG[8] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[8]), .Q(sa_snapshot[8]));
Q_FDP4EP \sa_snapshot_REG[9] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[9]), .Q(sa_snapshot[9]));
Q_FDP4EP \sa_snapshot_REG[10] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[10]), .Q(sa_snapshot[10]));
Q_FDP4EP \sa_snapshot_REG[11] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[11]), .Q(sa_snapshot[11]));
Q_FDP4EP \sa_snapshot_REG[12] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[12]), .Q(sa_snapshot[12]));
Q_FDP4EP \sa_snapshot_REG[13] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[13]), .Q(sa_snapshot[13]));
Q_FDP4EP \sa_snapshot_REG[14] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[14]), .Q(sa_snapshot[14]));
Q_FDP4EP \sa_snapshot_REG[15] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[15]), .Q(sa_snapshot[15]));
Q_FDP4EP \sa_snapshot_REG[16] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[16]), .Q(sa_snapshot[16]));
Q_FDP4EP \sa_snapshot_REG[17] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[17]), .Q(sa_snapshot[17]));
Q_FDP4EP \sa_snapshot_REG[18] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[18]), .Q(sa_snapshot[18]));
Q_FDP4EP \sa_snapshot_REG[19] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[19]), .Q(sa_snapshot[19]));
Q_FDP4EP \sa_snapshot_REG[20] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[20]), .Q(sa_snapshot[20]));
Q_FDP4EP \sa_snapshot_REG[21] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[21]), .Q(sa_snapshot[21]));
Q_FDP4EP \sa_snapshot_REG[22] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[22]), .Q(sa_snapshot[22]));
Q_FDP4EP \sa_snapshot_REG[23] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[23]), .Q(sa_snapshot[23]));
Q_FDP4EP \sa_snapshot_REG[24] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[24]), .Q(sa_snapshot[24]));
Q_FDP4EP \sa_snapshot_REG[25] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[25]), .Q(sa_snapshot[25]));
Q_FDP4EP \sa_snapshot_REG[26] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[26]), .Q(sa_snapshot[26]));
Q_FDP4EP \sa_snapshot_REG[27] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[27]), .Q(sa_snapshot[27]));
Q_FDP4EP \sa_snapshot_REG[28] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[28]), .Q(sa_snapshot[28]));
Q_FDP4EP \sa_snapshot_REG[29] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[29]), .Q(sa_snapshot[29]));
Q_FDP4EP \sa_snapshot_REG[30] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[30]), .Q(sa_snapshot[30]));
Q_FDP4EP \sa_snapshot_REG[31] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[31]), .Q(sa_snapshot[31]));
Q_FDP4EP \sa_snapshot_REG[32] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[32]), .Q(sa_snapshot[32]));
Q_FDP4EP \sa_snapshot_REG[33] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[33]), .Q(sa_snapshot[33]));
Q_FDP4EP \sa_snapshot_REG[34] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[34]), .Q(sa_snapshot[34]));
Q_FDP4EP \sa_snapshot_REG[35] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[35]), .Q(sa_snapshot[35]));
Q_FDP4EP \sa_snapshot_REG[36] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[36]), .Q(sa_snapshot[36]));
Q_FDP4EP \sa_snapshot_REG[37] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[37]), .Q(sa_snapshot[37]));
Q_FDP4EP \sa_snapshot_REG[38] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[38]), .Q(sa_snapshot[38]));
Q_FDP4EP \sa_snapshot_REG[39] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[39]), .Q(sa_snapshot[39]));
Q_FDP4EP \sa_snapshot_REG[40] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[40]), .Q(sa_snapshot[40]));
Q_FDP4EP \sa_snapshot_REG[41] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[41]), .Q(sa_snapshot[41]));
Q_FDP4EP \sa_snapshot_REG[42] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[42]), .Q(sa_snapshot[42]));
Q_FDP4EP \sa_snapshot_REG[43] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[43]), .Q(sa_snapshot[43]));
Q_FDP4EP \sa_snapshot_REG[44] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[44]), .Q(sa_snapshot[44]));
Q_FDP4EP \sa_snapshot_REG[45] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[45]), .Q(sa_snapshot[45]));
Q_FDP4EP \sa_snapshot_REG[46] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[46]), .Q(sa_snapshot[46]));
Q_FDP4EP \sa_snapshot_REG[47] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[47]), .Q(sa_snapshot[47]));
Q_FDP4EP \sa_snapshot_REG[48] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[48]), .Q(sa_snapshot[48]));
Q_FDP4EP \sa_snapshot_REG[49] ( .CK(clk), .CE(sa_snap), .R(n416), .D(sa_count[49]), .Q(sa_snapshot[49]));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "sa_events 1 63 0 15 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
endmodule
