library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
use work.cr_kme_regfilePKG.all ;
entity cr_kme_drbg_reggen is
  port (
    set_drbg_expired_int : out std_logic ;
    kdf_drbg_ctrl : out std_logic_vector(1 downto 0) ;
    seed0_valid : out std_logic ;
    seed0_internal_state_key : out std_logic_vector(255 downto 0) ;
    seed0_internal_state_value : out std_logic_vector(127 downto 0) ;
    seed0_reseed_interval : out std_logic_vector(47 downto 0) ;
    seed1_valid : out std_logic ;
    seed1_internal_state_key : out std_logic_vector(255 downto 0) ;
    seed1_internal_state_value : out std_logic_vector(127 downto 0) ;
    seed1_reseed_interval : out std_logic_vector(47 downto 0) ;
    clk : in std_logic ;
    rst_n : in std_logic ;
    wr_stb : in std_logic ;
    wr_data : in std_logic_vector(31 downto 0) ;
    reg_addr : in std_logic_vector(10 downto 0) ;
    o_kdf_drbg_ctrl : in std_logic_vector(1 downto 0) ;
    o_kdf_drbg_seed_0_reseed_interval_0 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_reseed_interval_1 : in std_logic_vector(15 downto 0) ;
    o_kdf_drbg_seed_0_state_key_127_96 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_159_128 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_191_160 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_223_192 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_255_224 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_31_0 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_63_32 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_key_95_64 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_value_127_96 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_value_31_0 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_value_63_32 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_0_state_value_95_64 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_reseed_interval_0 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_reseed_interval_1 : in std_logic_vector(15 downto 0) ;
    o_kdf_drbg_seed_1_state_key_127_96 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_159_128 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_191_160 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_223_192 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_255_224 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_31_0 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_63_32 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_key_95_64 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_value_127_96 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_value_31_0 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_value_63_32 : in std_logic_vector(31 downto 0) ;
    o_kdf_drbg_seed_1_state_value_95_64 : in std_logic_vector(31 downto 0) ;
    seed0_invalidate : in std_logic ;
  seed1_invalidate : in std_logic ) ;
  attribute _2_state_: integer;
end cr_kme_drbg_reggen ;
