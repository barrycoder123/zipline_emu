
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_tlvp2_rsm_core ( pt_ob_rd, tlvp_rsm_usr_ob_ren, tlvp_rsm_ob_wen, 
	.tlvp_rsm_ob_wdata( {\tlvp_rsm_ob_wdata.tvalid , 
	\tlvp_rsm_ob_wdata.tlast , \tlvp_rsm_ob_wdata.tid [0], 
	\tlvp_rsm_ob_wdata.tstrb [7], \tlvp_rsm_ob_wdata.tstrb [6], 
	\tlvp_rsm_ob_wdata.tstrb [5], \tlvp_rsm_ob_wdata.tstrb [4], 
	\tlvp_rsm_ob_wdata.tstrb [3], \tlvp_rsm_ob_wdata.tstrb [2], 
	\tlvp_rsm_ob_wdata.tstrb [1], \tlvp_rsm_ob_wdata.tstrb [0], 
	\tlvp_rsm_ob_wdata.tuser [7], \tlvp_rsm_ob_wdata.tuser [6], 
	\tlvp_rsm_ob_wdata.tuser [5], \tlvp_rsm_ob_wdata.tuser [4], 
	\tlvp_rsm_ob_wdata.tuser [3], \tlvp_rsm_ob_wdata.tuser [2], 
	\tlvp_rsm_ob_wdata.tuser [1], \tlvp_rsm_ob_wdata.tuser [0], 
	\tlvp_rsm_ob_wdata.tdata [63], \tlvp_rsm_ob_wdata.tdata [62], 
	\tlvp_rsm_ob_wdata.tdata [61], \tlvp_rsm_ob_wdata.tdata [60], 
	\tlvp_rsm_ob_wdata.tdata [59], \tlvp_rsm_ob_wdata.tdata [58], 
	\tlvp_rsm_ob_wdata.tdata [57], \tlvp_rsm_ob_wdata.tdata [56], 
	\tlvp_rsm_ob_wdata.tdata [55], \tlvp_rsm_ob_wdata.tdata [54], 
	\tlvp_rsm_ob_wdata.tdata [53], \tlvp_rsm_ob_wdata.tdata [52], 
	\tlvp_rsm_ob_wdata.tdata [51], \tlvp_rsm_ob_wdata.tdata [50], 
	\tlvp_rsm_ob_wdata.tdata [49], \tlvp_rsm_ob_wdata.tdata [48], 
	\tlvp_rsm_ob_wdata.tdata [47], \tlvp_rsm_ob_wdata.tdata [46], 
	\tlvp_rsm_ob_wdata.tdata [45], \tlvp_rsm_ob_wdata.tdata [44], 
	\tlvp_rsm_ob_wdata.tdata [43], \tlvp_rsm_ob_wdata.tdata [42], 
	\tlvp_rsm_ob_wdata.tdata [41], \tlvp_rsm_ob_wdata.tdata [40], 
	\tlvp_rsm_ob_wdata.tdata [39], \tlvp_rsm_ob_wdata.tdata [38], 
	\tlvp_rsm_ob_wdata.tdata [37], \tlvp_rsm_ob_wdata.tdata [36], 
	\tlvp_rsm_ob_wdata.tdata [35], \tlvp_rsm_ob_wdata.tdata [34], 
	\tlvp_rsm_ob_wdata.tdata [33], \tlvp_rsm_ob_wdata.tdata [32], 
	\tlvp_rsm_ob_wdata.tdata [31], \tlvp_rsm_ob_wdata.tdata [30], 
	\tlvp_rsm_ob_wdata.tdata [29], \tlvp_rsm_ob_wdata.tdata [28], 
	\tlvp_rsm_ob_wdata.tdata [27], \tlvp_rsm_ob_wdata.tdata [26], 
	\tlvp_rsm_ob_wdata.tdata [25], \tlvp_rsm_ob_wdata.tdata [24], 
	\tlvp_rsm_ob_wdata.tdata [23], \tlvp_rsm_ob_wdata.tdata [22], 
	\tlvp_rsm_ob_wdata.tdata [21], \tlvp_rsm_ob_wdata.tdata [20], 
	\tlvp_rsm_ob_wdata.tdata [19], \tlvp_rsm_ob_wdata.tdata [18], 
	\tlvp_rsm_ob_wdata.tdata [17], \tlvp_rsm_ob_wdata.tdata [16], 
	\tlvp_rsm_ob_wdata.tdata [15], \tlvp_rsm_ob_wdata.tdata [14], 
	\tlvp_rsm_ob_wdata.tdata [13], \tlvp_rsm_ob_wdata.tdata [12], 
	\tlvp_rsm_ob_wdata.tdata [11], \tlvp_rsm_ob_wdata.tdata [10], 
	\tlvp_rsm_ob_wdata.tdata [9], \tlvp_rsm_ob_wdata.tdata [8], 
	\tlvp_rsm_ob_wdata.tdata [7], \tlvp_rsm_ob_wdata.tdata [6], 
	\tlvp_rsm_ob_wdata.tdata [5], \tlvp_rsm_ob_wdata.tdata [4], 
	\tlvp_rsm_ob_wdata.tdata [3], \tlvp_rsm_ob_wdata.tdata [2], 
	\tlvp_rsm_ob_wdata.tdata [1], \tlvp_rsm_ob_wdata.tdata [0]} ), clk, 
	rst_n, pt_ob_empty, pt_ob_aempty, .pt_ob_tlv( {\pt_ob_tlv.insert , 
	\pt_ob_tlv.ordern [12], \pt_ob_tlv.ordern [11], 
	\pt_ob_tlv.ordern [10], \pt_ob_tlv.ordern [9], \pt_ob_tlv.ordern [8], 
	\pt_ob_tlv.ordern [7], \pt_ob_tlv.ordern [6], \pt_ob_tlv.ordern [5], 
	\pt_ob_tlv.ordern [4], \pt_ob_tlv.ordern [3], \pt_ob_tlv.ordern [2], 
	\pt_ob_tlv.ordern [1], \pt_ob_tlv.ordern [0], \pt_ob_tlv.typen [7], 
	\pt_ob_tlv.typen [6], \pt_ob_tlv.typen [5], \pt_ob_tlv.typen [4], 
	\pt_ob_tlv.typen [3], \pt_ob_tlv.typen [2], \pt_ob_tlv.typen [1], 
	\pt_ob_tlv.typen [0], \pt_ob_tlv.sot , \pt_ob_tlv.eot , 
	\pt_ob_tlv.tlast , \pt_ob_tlv.tid [0], \pt_ob_tlv.tstrb [7], 
	\pt_ob_tlv.tstrb [6], \pt_ob_tlv.tstrb [5], \pt_ob_tlv.tstrb [4], 
	\pt_ob_tlv.tstrb [3], \pt_ob_tlv.tstrb [2], \pt_ob_tlv.tstrb [1], 
	\pt_ob_tlv.tstrb [0], \pt_ob_tlv.tuser [7], \pt_ob_tlv.tuser [6], 
	\pt_ob_tlv.tuser [5], \pt_ob_tlv.tuser [4], \pt_ob_tlv.tuser [3], 
	\pt_ob_tlv.tuser [2], \pt_ob_tlv.tuser [1], \pt_ob_tlv.tuser [0], 
	\pt_ob_tlv.tdata [63], \pt_ob_tlv.tdata [62], \pt_ob_tlv.tdata [61], 
	\pt_ob_tlv.tdata [60], \pt_ob_tlv.tdata [59], \pt_ob_tlv.tdata [58], 
	\pt_ob_tlv.tdata [57], \pt_ob_tlv.tdata [56], \pt_ob_tlv.tdata [55], 
	\pt_ob_tlv.tdata [54], \pt_ob_tlv.tdata [53], \pt_ob_tlv.tdata [52], 
	\pt_ob_tlv.tdata [51], \pt_ob_tlv.tdata [50], \pt_ob_tlv.tdata [49], 
	\pt_ob_tlv.tdata [48], \pt_ob_tlv.tdata [47], \pt_ob_tlv.tdata [46], 
	\pt_ob_tlv.tdata [45], \pt_ob_tlv.tdata [44], \pt_ob_tlv.tdata [43], 
	\pt_ob_tlv.tdata [42], \pt_ob_tlv.tdata [41], \pt_ob_tlv.tdata [40], 
	\pt_ob_tlv.tdata [39], \pt_ob_tlv.tdata [38], \pt_ob_tlv.tdata [37], 
	\pt_ob_tlv.tdata [36], \pt_ob_tlv.tdata [35], \pt_ob_tlv.tdata [34], 
	\pt_ob_tlv.tdata [33], \pt_ob_tlv.tdata [32], \pt_ob_tlv.tdata [31], 
	\pt_ob_tlv.tdata [30], \pt_ob_tlv.tdata [29], \pt_ob_tlv.tdata [28], 
	\pt_ob_tlv.tdata [27], \pt_ob_tlv.tdata [26], \pt_ob_tlv.tdata [25], 
	\pt_ob_tlv.tdata [24], \pt_ob_tlv.tdata [23], \pt_ob_tlv.tdata [22], 
	\pt_ob_tlv.tdata [21], \pt_ob_tlv.tdata [20], \pt_ob_tlv.tdata [19], 
	\pt_ob_tlv.tdata [18], \pt_ob_tlv.tdata [17], \pt_ob_tlv.tdata [16], 
	\pt_ob_tlv.tdata [15], \pt_ob_tlv.tdata [14], \pt_ob_tlv.tdata [13], 
	\pt_ob_tlv.tdata [12], \pt_ob_tlv.tdata [11], \pt_ob_tlv.tdata [10], 
	\pt_ob_tlv.tdata [9], \pt_ob_tlv.tdata [8], \pt_ob_tlv.tdata [7], 
	\pt_ob_tlv.tdata [6], \pt_ob_tlv.tdata [5], \pt_ob_tlv.tdata [4], 
	\pt_ob_tlv.tdata [3], \pt_ob_tlv.tdata [2], \pt_ob_tlv.tdata [1], 
	\pt_ob_tlv.tdata [0]} ), .tlvp_rsm_usr_ob_rdata( {
	\tlvp_rsm_usr_ob_rdata.insert , \tlvp_rsm_usr_ob_rdata.ordern [12], 
	\tlvp_rsm_usr_ob_rdata.ordern [11], 
	\tlvp_rsm_usr_ob_rdata.ordern [10], 
	\tlvp_rsm_usr_ob_rdata.ordern [9], \tlvp_rsm_usr_ob_rdata.ordern [8], 
	\tlvp_rsm_usr_ob_rdata.ordern [7], \tlvp_rsm_usr_ob_rdata.ordern [6], 
	\tlvp_rsm_usr_ob_rdata.ordern [5], \tlvp_rsm_usr_ob_rdata.ordern [4], 
	\tlvp_rsm_usr_ob_rdata.ordern [3], \tlvp_rsm_usr_ob_rdata.ordern [2], 
	\tlvp_rsm_usr_ob_rdata.ordern [1], \tlvp_rsm_usr_ob_rdata.ordern [0], 
	\tlvp_rsm_usr_ob_rdata.typen [7], \tlvp_rsm_usr_ob_rdata.typen [6], 
	\tlvp_rsm_usr_ob_rdata.typen [5], \tlvp_rsm_usr_ob_rdata.typen [4], 
	\tlvp_rsm_usr_ob_rdata.typen [3], \tlvp_rsm_usr_ob_rdata.typen [2], 
	\tlvp_rsm_usr_ob_rdata.typen [1], \tlvp_rsm_usr_ob_rdata.typen [0], 
	\tlvp_rsm_usr_ob_rdata.sot , \tlvp_rsm_usr_ob_rdata.eot , 
	\tlvp_rsm_usr_ob_rdata.tlast , \tlvp_rsm_usr_ob_rdata.tid [0], 
	\tlvp_rsm_usr_ob_rdata.tstrb [7], \tlvp_rsm_usr_ob_rdata.tstrb [6], 
	\tlvp_rsm_usr_ob_rdata.tstrb [5], \tlvp_rsm_usr_ob_rdata.tstrb [4], 
	\tlvp_rsm_usr_ob_rdata.tstrb [3], \tlvp_rsm_usr_ob_rdata.tstrb [2], 
	\tlvp_rsm_usr_ob_rdata.tstrb [1], \tlvp_rsm_usr_ob_rdata.tstrb [0], 
	\tlvp_rsm_usr_ob_rdata.tuser [7], \tlvp_rsm_usr_ob_rdata.tuser [6], 
	\tlvp_rsm_usr_ob_rdata.tuser [5], \tlvp_rsm_usr_ob_rdata.tuser [4], 
	\tlvp_rsm_usr_ob_rdata.tuser [3], \tlvp_rsm_usr_ob_rdata.tuser [2], 
	\tlvp_rsm_usr_ob_rdata.tuser [1], \tlvp_rsm_usr_ob_rdata.tuser [0], 
	\tlvp_rsm_usr_ob_rdata.tdata [63], \tlvp_rsm_usr_ob_rdata.tdata [62], 
	\tlvp_rsm_usr_ob_rdata.tdata [61], \tlvp_rsm_usr_ob_rdata.tdata [60], 
	\tlvp_rsm_usr_ob_rdata.tdata [59], \tlvp_rsm_usr_ob_rdata.tdata [58], 
	\tlvp_rsm_usr_ob_rdata.tdata [57], \tlvp_rsm_usr_ob_rdata.tdata [56], 
	\tlvp_rsm_usr_ob_rdata.tdata [55], \tlvp_rsm_usr_ob_rdata.tdata [54], 
	\tlvp_rsm_usr_ob_rdata.tdata [53], \tlvp_rsm_usr_ob_rdata.tdata [52], 
	\tlvp_rsm_usr_ob_rdata.tdata [51], \tlvp_rsm_usr_ob_rdata.tdata [50], 
	\tlvp_rsm_usr_ob_rdata.tdata [49], \tlvp_rsm_usr_ob_rdata.tdata [48], 
	\tlvp_rsm_usr_ob_rdata.tdata [47], \tlvp_rsm_usr_ob_rdata.tdata [46], 
	\tlvp_rsm_usr_ob_rdata.tdata [45], \tlvp_rsm_usr_ob_rdata.tdata [44], 
	\tlvp_rsm_usr_ob_rdata.tdata [43], \tlvp_rsm_usr_ob_rdata.tdata [42], 
	\tlvp_rsm_usr_ob_rdata.tdata [41], \tlvp_rsm_usr_ob_rdata.tdata [40], 
	\tlvp_rsm_usr_ob_rdata.tdata [39], \tlvp_rsm_usr_ob_rdata.tdata [38], 
	\tlvp_rsm_usr_ob_rdata.tdata [37], \tlvp_rsm_usr_ob_rdata.tdata [36], 
	\tlvp_rsm_usr_ob_rdata.tdata [35], \tlvp_rsm_usr_ob_rdata.tdata [34], 
	\tlvp_rsm_usr_ob_rdata.tdata [33], \tlvp_rsm_usr_ob_rdata.tdata [32], 
	\tlvp_rsm_usr_ob_rdata.tdata [31], \tlvp_rsm_usr_ob_rdata.tdata [30], 
	\tlvp_rsm_usr_ob_rdata.tdata [29], \tlvp_rsm_usr_ob_rdata.tdata [28], 
	\tlvp_rsm_usr_ob_rdata.tdata [27], \tlvp_rsm_usr_ob_rdata.tdata [26], 
	\tlvp_rsm_usr_ob_rdata.tdata [25], \tlvp_rsm_usr_ob_rdata.tdata [24], 
	\tlvp_rsm_usr_ob_rdata.tdata [23], \tlvp_rsm_usr_ob_rdata.tdata [22], 
	\tlvp_rsm_usr_ob_rdata.tdata [21], \tlvp_rsm_usr_ob_rdata.tdata [20], 
	\tlvp_rsm_usr_ob_rdata.tdata [19], \tlvp_rsm_usr_ob_rdata.tdata [18], 
	\tlvp_rsm_usr_ob_rdata.tdata [17], \tlvp_rsm_usr_ob_rdata.tdata [16], 
	\tlvp_rsm_usr_ob_rdata.tdata [15], \tlvp_rsm_usr_ob_rdata.tdata [14], 
	\tlvp_rsm_usr_ob_rdata.tdata [13], \tlvp_rsm_usr_ob_rdata.tdata [12], 
	\tlvp_rsm_usr_ob_rdata.tdata [11], \tlvp_rsm_usr_ob_rdata.tdata [10], 
	\tlvp_rsm_usr_ob_rdata.tdata [9], \tlvp_rsm_usr_ob_rdata.tdata [8], 
	\tlvp_rsm_usr_ob_rdata.tdata [7], \tlvp_rsm_usr_ob_rdata.tdata [6], 
	\tlvp_rsm_usr_ob_rdata.tdata [5], \tlvp_rsm_usr_ob_rdata.tdata [4], 
	\tlvp_rsm_usr_ob_rdata.tdata [3], \tlvp_rsm_usr_ob_rdata.tdata [2], 
	\tlvp_rsm_usr_ob_rdata.tdata [1], \tlvp_rsm_usr_ob_rdata.tdata [0]} ), 
	usr_ob_empty, usr_ob_aempty, tlvp_ob_full, tlvp_ob_afull);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output pt_ob_rd;
output tlvp_rsm_usr_ob_ren;
output tlvp_rsm_ob_wen;
output \tlvp_rsm_ob_wdata.tvalid ;
output \tlvp_rsm_ob_wdata.tlast ;
output [0:0] \tlvp_rsm_ob_wdata.tid ;
output [7:0] \tlvp_rsm_ob_wdata.tstrb ;
output [7:0] \tlvp_rsm_ob_wdata.tuser ;
output [63:0] \tlvp_rsm_ob_wdata.tdata ;
wire [82:0] tlvp_rsm_ob_wdata;
input clk;
input rst_n;
input pt_ob_empty;
input pt_ob_aempty;
input \pt_ob_tlv.insert ;
input [12:0] \pt_ob_tlv.ordern ;
input [7:0] \pt_ob_tlv.typen ;
input \pt_ob_tlv.sot ;
input \pt_ob_tlv.eot ;
input \pt_ob_tlv.tlast ;
input [0:0] \pt_ob_tlv.tid ;
input [7:0] \pt_ob_tlv.tstrb ;
input [7:0] \pt_ob_tlv.tuser ;
input [63:0] \pt_ob_tlv.tdata ;
wire [105:0] pt_ob_tlv;
input \tlvp_rsm_usr_ob_rdata.insert ;
input [12:0] \tlvp_rsm_usr_ob_rdata.ordern ;
input [7:0] \tlvp_rsm_usr_ob_rdata.typen ;
input \tlvp_rsm_usr_ob_rdata.sot ;
input \tlvp_rsm_usr_ob_rdata.eot ;
input \tlvp_rsm_usr_ob_rdata.tlast ;
input [0:0] \tlvp_rsm_usr_ob_rdata.tid ;
input [7:0] \tlvp_rsm_usr_ob_rdata.tstrb ;
input [7:0] \tlvp_rsm_usr_ob_rdata.tuser ;
input [63:0] \tlvp_rsm_usr_ob_rdata.tdata ;
wire [105:0] tlvp_rsm_usr_ob_rdata;
input usr_ob_empty;
input usr_ob_aempty;
input tlvp_ob_full;
input tlvp_ob_afull;
wire _zy_simnet_pt_ob_rd_0_w$;
wire _zy_simnet_tlvp_rsm_usr_ob_ren_1_w$;
wire _zy_simnet_tlvp_rsm_ob_wen_2_w$;
wire [0:82] _zy_simnet_tlvp_rsm_ob_wdata_3_w$;
wire [63:0] tlvp_rsm_usr_ob_rdata_dw0;
wire [1:0] tlvp_rsm_bip2;
wire tlvp_rsm_usr_ob_valid;
wire [105:0] tlvp_rsm_usr_ob_tlv;
wire tlvp_rsm_usr_ob_wen;
wire tlvp_rsm_usr_ob_sel;
wire tlvp_rsm_pt_valid;
wire [105:0] tlvp_rsm_pt_tlv;
wire tlvp_rsm_pt_wen;
wire tlvp_rsm_pt_sel;
wire [105:0] tlvp_rsm_ob_datain;
wire [12:0] tlvp_rsm_nxt_ordern;
wire [7:0] tlvp_rsm_last_typen;
wire tlvp_rsm_pt_next;
wire tlvp_rsm_usr_ob_next;
wire tlvp_rsm_usr_insert;
wire [1:0] tlvp_rsm_selector;
wire [12:0] tlvp_rsm_usr_ob_tlv_ordern;
wire [12:0] tlvp_rsm_pt_tlv_ordern;
wire [31:0] current_state;
wire [31:0] next_state;
supply0 n1;
wire [1:0] \tlvp_rsm_usr_ob_rdata_dw0.tlv_bip2 ;
wire [18:0] \tlvp_rsm_usr_ob_rdata_dw0.resv0 ;
wire [10:0] \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num ;
wire [3:0] \tlvp_rsm_usr_ob_rdata_dw0.resv1 ;
wire [3:0] \tlvp_rsm_usr_ob_rdata_dw0.tlv_eng_id ;
wire [7:0] \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num ;
wire [7:0] \tlvp_rsm_usr_ob_rdata_dw0.tlv_len ;
wire [7:0] \tlvp_rsm_usr_ob_rdata_dw0.tlv_type ;
wire \tlvp_rsm_usr_ob_tlv.insert ;
wire [12:0] \tlvp_rsm_usr_ob_tlv.ordern ;
wire [7:0] \tlvp_rsm_usr_ob_tlv.typen ;
wire \tlvp_rsm_usr_ob_tlv.sot ;
wire \tlvp_rsm_usr_ob_tlv.eot ;
wire \tlvp_rsm_usr_ob_tlv.tlast ;
wire [0:0] \tlvp_rsm_usr_ob_tlv.tid ;
wire [7:0] \tlvp_rsm_usr_ob_tlv.tstrb ;
wire [7:0] \tlvp_rsm_usr_ob_tlv.tuser ;
wire [63:0] \tlvp_rsm_usr_ob_tlv.tdata ;
wire \tlvp_rsm_pt_tlv.insert ;
wire [12:0] \tlvp_rsm_pt_tlv.ordern ;
wire [7:0] \tlvp_rsm_pt_tlv.typen ;
wire \tlvp_rsm_pt_tlv.sot ;
wire \tlvp_rsm_pt_tlv.eot ;
wire \tlvp_rsm_pt_tlv.tlast ;
wire [0:0] \tlvp_rsm_pt_tlv.tid ;
wire [7:0] \tlvp_rsm_pt_tlv.tstrb ;
wire [7:0] \tlvp_rsm_pt_tlv.tuser ;
wire [63:0] \tlvp_rsm_pt_tlv.tdata ;
wire \tlvp_rsm_ob_datain.insert ;
wire [12:0] \tlvp_rsm_ob_datain.ordern ;
wire [7:0] \tlvp_rsm_ob_datain.typen ;
wire \tlvp_rsm_ob_datain.sot ;
wire \tlvp_rsm_ob_datain.eot ;
wire \tlvp_rsm_ob_datain.tlast ;
wire [0:0] \tlvp_rsm_ob_datain.tid ;
wire [7:0] \tlvp_rsm_ob_datain.tstrb ;
wire [7:0] \tlvp_rsm_ob_datain.tuser ;
wire [63:0] \tlvp_rsm_ob_datain.tdata ;
tran (tlvp_rsm_ob_wdata[82], \tlvp_rsm_ob_wdata.tvalid );
tran (tlvp_rsm_ob_wdata[81], \tlvp_rsm_ob_wdata.tlast );
tran (tlvp_rsm_ob_wdata[80], \tlvp_rsm_ob_wdata.tid [0]);
tran (tlvp_rsm_ob_wdata[79], \tlvp_rsm_ob_wdata.tstrb [7]);
tran (tlvp_rsm_ob_wdata[78], \tlvp_rsm_ob_wdata.tstrb [6]);
tran (tlvp_rsm_ob_wdata[77], \tlvp_rsm_ob_wdata.tstrb [5]);
tran (tlvp_rsm_ob_wdata[76], \tlvp_rsm_ob_wdata.tstrb [4]);
tran (tlvp_rsm_ob_wdata[75], \tlvp_rsm_ob_wdata.tstrb [3]);
tran (tlvp_rsm_ob_wdata[74], \tlvp_rsm_ob_wdata.tstrb [2]);
tran (tlvp_rsm_ob_wdata[73], \tlvp_rsm_ob_wdata.tstrb [1]);
tran (tlvp_rsm_ob_wdata[72], \tlvp_rsm_ob_wdata.tstrb [0]);
tran (tlvp_rsm_ob_wdata[71], \tlvp_rsm_ob_wdata.tuser [7]);
tran (tlvp_rsm_ob_wdata[70], \tlvp_rsm_ob_wdata.tuser [6]);
tran (tlvp_rsm_ob_wdata[69], \tlvp_rsm_ob_wdata.tuser [5]);
tran (tlvp_rsm_ob_wdata[68], \tlvp_rsm_ob_wdata.tuser [4]);
tran (tlvp_rsm_ob_wdata[67], \tlvp_rsm_ob_wdata.tuser [3]);
tran (tlvp_rsm_ob_wdata[66], \tlvp_rsm_ob_wdata.tuser [2]);
tran (tlvp_rsm_ob_wdata[65], \tlvp_rsm_ob_wdata.tuser [1]);
tran (tlvp_rsm_ob_wdata[64], \tlvp_rsm_ob_wdata.tuser [0]);
tran (tlvp_rsm_ob_wdata[63], \tlvp_rsm_ob_wdata.tdata [63]);
tran (tlvp_rsm_ob_wdata[62], \tlvp_rsm_ob_wdata.tdata [62]);
tran (tlvp_rsm_ob_wdata[61], \tlvp_rsm_ob_wdata.tdata [61]);
tran (tlvp_rsm_ob_wdata[60], \tlvp_rsm_ob_wdata.tdata [60]);
tran (tlvp_rsm_ob_wdata[59], \tlvp_rsm_ob_wdata.tdata [59]);
tran (tlvp_rsm_ob_wdata[58], \tlvp_rsm_ob_wdata.tdata [58]);
tran (tlvp_rsm_ob_wdata[57], \tlvp_rsm_ob_wdata.tdata [57]);
tran (tlvp_rsm_ob_wdata[56], \tlvp_rsm_ob_wdata.tdata [56]);
tran (tlvp_rsm_ob_wdata[55], \tlvp_rsm_ob_wdata.tdata [55]);
tran (tlvp_rsm_ob_wdata[54], \tlvp_rsm_ob_wdata.tdata [54]);
tran (tlvp_rsm_ob_wdata[53], \tlvp_rsm_ob_wdata.tdata [53]);
tran (tlvp_rsm_ob_wdata[52], \tlvp_rsm_ob_wdata.tdata [52]);
tran (tlvp_rsm_ob_wdata[51], \tlvp_rsm_ob_wdata.tdata [51]);
tran (tlvp_rsm_ob_wdata[50], \tlvp_rsm_ob_wdata.tdata [50]);
tran (tlvp_rsm_ob_wdata[49], \tlvp_rsm_ob_wdata.tdata [49]);
tran (tlvp_rsm_ob_wdata[48], \tlvp_rsm_ob_wdata.tdata [48]);
tran (tlvp_rsm_ob_wdata[47], \tlvp_rsm_ob_wdata.tdata [47]);
tran (tlvp_rsm_ob_wdata[46], \tlvp_rsm_ob_wdata.tdata [46]);
tran (tlvp_rsm_ob_wdata[45], \tlvp_rsm_ob_wdata.tdata [45]);
tran (tlvp_rsm_ob_wdata[44], \tlvp_rsm_ob_wdata.tdata [44]);
tran (tlvp_rsm_ob_wdata[43], \tlvp_rsm_ob_wdata.tdata [43]);
tran (tlvp_rsm_ob_wdata[42], \tlvp_rsm_ob_wdata.tdata [42]);
tran (tlvp_rsm_ob_wdata[41], \tlvp_rsm_ob_wdata.tdata [41]);
tran (tlvp_rsm_ob_wdata[40], \tlvp_rsm_ob_wdata.tdata [40]);
tran (tlvp_rsm_ob_wdata[39], \tlvp_rsm_ob_wdata.tdata [39]);
tran (tlvp_rsm_ob_wdata[38], \tlvp_rsm_ob_wdata.tdata [38]);
tran (tlvp_rsm_ob_wdata[37], \tlvp_rsm_ob_wdata.tdata [37]);
tran (tlvp_rsm_ob_wdata[36], \tlvp_rsm_ob_wdata.tdata [36]);
tran (tlvp_rsm_ob_wdata[35], \tlvp_rsm_ob_wdata.tdata [35]);
tran (tlvp_rsm_ob_wdata[34], \tlvp_rsm_ob_wdata.tdata [34]);
tran (tlvp_rsm_ob_wdata[33], \tlvp_rsm_ob_wdata.tdata [33]);
tran (tlvp_rsm_ob_wdata[32], \tlvp_rsm_ob_wdata.tdata [32]);
tran (tlvp_rsm_ob_wdata[31], \tlvp_rsm_ob_wdata.tdata [31]);
tran (tlvp_rsm_ob_wdata[30], \tlvp_rsm_ob_wdata.tdata [30]);
tran (tlvp_rsm_ob_wdata[29], \tlvp_rsm_ob_wdata.tdata [29]);
tran (tlvp_rsm_ob_wdata[28], \tlvp_rsm_ob_wdata.tdata [28]);
tran (tlvp_rsm_ob_wdata[27], \tlvp_rsm_ob_wdata.tdata [27]);
tran (tlvp_rsm_ob_wdata[26], \tlvp_rsm_ob_wdata.tdata [26]);
tran (tlvp_rsm_ob_wdata[25], \tlvp_rsm_ob_wdata.tdata [25]);
tran (tlvp_rsm_ob_wdata[24], \tlvp_rsm_ob_wdata.tdata [24]);
tran (tlvp_rsm_ob_wdata[23], \tlvp_rsm_ob_wdata.tdata [23]);
tran (tlvp_rsm_ob_wdata[22], \tlvp_rsm_ob_wdata.tdata [22]);
tran (tlvp_rsm_ob_wdata[21], \tlvp_rsm_ob_wdata.tdata [21]);
tran (tlvp_rsm_ob_wdata[20], \tlvp_rsm_ob_wdata.tdata [20]);
tran (tlvp_rsm_ob_wdata[19], \tlvp_rsm_ob_wdata.tdata [19]);
tran (tlvp_rsm_ob_wdata[18], \tlvp_rsm_ob_wdata.tdata [18]);
tran (tlvp_rsm_ob_wdata[17], \tlvp_rsm_ob_wdata.tdata [17]);
tran (tlvp_rsm_ob_wdata[16], \tlvp_rsm_ob_wdata.tdata [16]);
tran (tlvp_rsm_ob_wdata[15], \tlvp_rsm_ob_wdata.tdata [15]);
tran (tlvp_rsm_ob_wdata[14], \tlvp_rsm_ob_wdata.tdata [14]);
tran (tlvp_rsm_ob_wdata[13], \tlvp_rsm_ob_wdata.tdata [13]);
tran (tlvp_rsm_ob_wdata[12], \tlvp_rsm_ob_wdata.tdata [12]);
tran (tlvp_rsm_ob_wdata[11], \tlvp_rsm_ob_wdata.tdata [11]);
tran (tlvp_rsm_ob_wdata[10], \tlvp_rsm_ob_wdata.tdata [10]);
tran (tlvp_rsm_ob_wdata[9], \tlvp_rsm_ob_wdata.tdata [9]);
tran (tlvp_rsm_ob_wdata[8], \tlvp_rsm_ob_wdata.tdata [8]);
tran (tlvp_rsm_ob_wdata[7], \tlvp_rsm_ob_wdata.tdata [7]);
tran (tlvp_rsm_ob_wdata[6], \tlvp_rsm_ob_wdata.tdata [6]);
tran (tlvp_rsm_ob_wdata[5], \tlvp_rsm_ob_wdata.tdata [5]);
tran (tlvp_rsm_ob_wdata[4], \tlvp_rsm_ob_wdata.tdata [4]);
tran (tlvp_rsm_ob_wdata[3], \tlvp_rsm_ob_wdata.tdata [3]);
tran (tlvp_rsm_ob_wdata[2], \tlvp_rsm_ob_wdata.tdata [2]);
tran (tlvp_rsm_ob_wdata[1], \tlvp_rsm_ob_wdata.tdata [1]);
tran (tlvp_rsm_ob_wdata[0], \tlvp_rsm_ob_wdata.tdata [0]);
tran (pt_ob_tlv[105], \pt_ob_tlv.insert );
tran (pt_ob_tlv[104], \pt_ob_tlv.ordern [12]);
tran (pt_ob_tlv[103], \pt_ob_tlv.ordern [11]);
tran (pt_ob_tlv[102], \pt_ob_tlv.ordern [10]);
tran (pt_ob_tlv[101], \pt_ob_tlv.ordern [9]);
tran (pt_ob_tlv[100], \pt_ob_tlv.ordern [8]);
tran (pt_ob_tlv[99], \pt_ob_tlv.ordern [7]);
tran (pt_ob_tlv[98], \pt_ob_tlv.ordern [6]);
tran (pt_ob_tlv[97], \pt_ob_tlv.ordern [5]);
tran (pt_ob_tlv[96], \pt_ob_tlv.ordern [4]);
tran (pt_ob_tlv[95], \pt_ob_tlv.ordern [3]);
tran (pt_ob_tlv[94], \pt_ob_tlv.ordern [2]);
tran (pt_ob_tlv[93], \pt_ob_tlv.ordern [1]);
tran (pt_ob_tlv[92], \pt_ob_tlv.ordern [0]);
tran (pt_ob_tlv[91], \pt_ob_tlv.typen [7]);
tran (pt_ob_tlv[90], \pt_ob_tlv.typen [6]);
tran (pt_ob_tlv[89], \pt_ob_tlv.typen [5]);
tran (pt_ob_tlv[88], \pt_ob_tlv.typen [4]);
tran (pt_ob_tlv[87], \pt_ob_tlv.typen [3]);
tran (pt_ob_tlv[86], \pt_ob_tlv.typen [2]);
tran (pt_ob_tlv[85], \pt_ob_tlv.typen [1]);
tran (pt_ob_tlv[84], \pt_ob_tlv.typen [0]);
tran (pt_ob_tlv[83], \pt_ob_tlv.sot );
tran (pt_ob_tlv[82], \pt_ob_tlv.eot );
tran (pt_ob_tlv[81], \pt_ob_tlv.tlast );
tran (pt_ob_tlv[80], \pt_ob_tlv.tid [0]);
tran (pt_ob_tlv[79], \pt_ob_tlv.tstrb [7]);
tran (pt_ob_tlv[78], \pt_ob_tlv.tstrb [6]);
tran (pt_ob_tlv[77], \pt_ob_tlv.tstrb [5]);
tran (pt_ob_tlv[76], \pt_ob_tlv.tstrb [4]);
tran (pt_ob_tlv[75], \pt_ob_tlv.tstrb [3]);
tran (pt_ob_tlv[74], \pt_ob_tlv.tstrb [2]);
tran (pt_ob_tlv[73], \pt_ob_tlv.tstrb [1]);
tran (pt_ob_tlv[72], \pt_ob_tlv.tstrb [0]);
tran (pt_ob_tlv[71], \pt_ob_tlv.tuser [7]);
tran (pt_ob_tlv[70], \pt_ob_tlv.tuser [6]);
tran (pt_ob_tlv[69], \pt_ob_tlv.tuser [5]);
tran (pt_ob_tlv[68], \pt_ob_tlv.tuser [4]);
tran (pt_ob_tlv[67], \pt_ob_tlv.tuser [3]);
tran (pt_ob_tlv[66], \pt_ob_tlv.tuser [2]);
tran (pt_ob_tlv[65], \pt_ob_tlv.tuser [1]);
tran (pt_ob_tlv[64], \pt_ob_tlv.tuser [0]);
tran (pt_ob_tlv[63], \pt_ob_tlv.tdata [63]);
tran (pt_ob_tlv[62], \pt_ob_tlv.tdata [62]);
tran (pt_ob_tlv[61], \pt_ob_tlv.tdata [61]);
tran (pt_ob_tlv[60], \pt_ob_tlv.tdata [60]);
tran (pt_ob_tlv[59], \pt_ob_tlv.tdata [59]);
tran (pt_ob_tlv[58], \pt_ob_tlv.tdata [58]);
tran (pt_ob_tlv[57], \pt_ob_tlv.tdata [57]);
tran (pt_ob_tlv[56], \pt_ob_tlv.tdata [56]);
tran (pt_ob_tlv[55], \pt_ob_tlv.tdata [55]);
tran (pt_ob_tlv[54], \pt_ob_tlv.tdata [54]);
tran (pt_ob_tlv[53], \pt_ob_tlv.tdata [53]);
tran (pt_ob_tlv[52], \pt_ob_tlv.tdata [52]);
tran (pt_ob_tlv[51], \pt_ob_tlv.tdata [51]);
tran (pt_ob_tlv[50], \pt_ob_tlv.tdata [50]);
tran (pt_ob_tlv[49], \pt_ob_tlv.tdata [49]);
tran (pt_ob_tlv[48], \pt_ob_tlv.tdata [48]);
tran (pt_ob_tlv[47], \pt_ob_tlv.tdata [47]);
tran (pt_ob_tlv[46], \pt_ob_tlv.tdata [46]);
tran (pt_ob_tlv[45], \pt_ob_tlv.tdata [45]);
tran (pt_ob_tlv[44], \pt_ob_tlv.tdata [44]);
tran (pt_ob_tlv[43], \pt_ob_tlv.tdata [43]);
tran (pt_ob_tlv[42], \pt_ob_tlv.tdata [42]);
tran (pt_ob_tlv[41], \pt_ob_tlv.tdata [41]);
tran (pt_ob_tlv[40], \pt_ob_tlv.tdata [40]);
tran (pt_ob_tlv[39], \pt_ob_tlv.tdata [39]);
tran (pt_ob_tlv[38], \pt_ob_tlv.tdata [38]);
tran (pt_ob_tlv[37], \pt_ob_tlv.tdata [37]);
tran (pt_ob_tlv[36], \pt_ob_tlv.tdata [36]);
tran (pt_ob_tlv[35], \pt_ob_tlv.tdata [35]);
tran (pt_ob_tlv[34], \pt_ob_tlv.tdata [34]);
tran (pt_ob_tlv[33], \pt_ob_tlv.tdata [33]);
tran (pt_ob_tlv[32], \pt_ob_tlv.tdata [32]);
tran (pt_ob_tlv[31], \pt_ob_tlv.tdata [31]);
tran (pt_ob_tlv[30], \pt_ob_tlv.tdata [30]);
tran (pt_ob_tlv[29], \pt_ob_tlv.tdata [29]);
tran (pt_ob_tlv[28], \pt_ob_tlv.tdata [28]);
tran (pt_ob_tlv[27], \pt_ob_tlv.tdata [27]);
tran (pt_ob_tlv[26], \pt_ob_tlv.tdata [26]);
tran (pt_ob_tlv[25], \pt_ob_tlv.tdata [25]);
tran (pt_ob_tlv[24], \pt_ob_tlv.tdata [24]);
tran (pt_ob_tlv[23], \pt_ob_tlv.tdata [23]);
tran (pt_ob_tlv[22], \pt_ob_tlv.tdata [22]);
tran (pt_ob_tlv[21], \pt_ob_tlv.tdata [21]);
tran (pt_ob_tlv[20], \pt_ob_tlv.tdata [20]);
tran (pt_ob_tlv[19], \pt_ob_tlv.tdata [19]);
tran (pt_ob_tlv[18], \pt_ob_tlv.tdata [18]);
tran (pt_ob_tlv[17], \pt_ob_tlv.tdata [17]);
tran (pt_ob_tlv[16], \pt_ob_tlv.tdata [16]);
tran (pt_ob_tlv[15], \pt_ob_tlv.tdata [15]);
tran (pt_ob_tlv[14], \pt_ob_tlv.tdata [14]);
tran (pt_ob_tlv[13], \pt_ob_tlv.tdata [13]);
tran (pt_ob_tlv[12], \pt_ob_tlv.tdata [12]);
tran (pt_ob_tlv[11], \pt_ob_tlv.tdata [11]);
tran (pt_ob_tlv[10], \pt_ob_tlv.tdata [10]);
tran (pt_ob_tlv[9], \pt_ob_tlv.tdata [9]);
tran (pt_ob_tlv[8], \pt_ob_tlv.tdata [8]);
tran (pt_ob_tlv[7], \pt_ob_tlv.tdata [7]);
tran (pt_ob_tlv[6], \pt_ob_tlv.tdata [6]);
tran (pt_ob_tlv[5], \pt_ob_tlv.tdata [5]);
tran (pt_ob_tlv[4], \pt_ob_tlv.tdata [4]);
tran (pt_ob_tlv[3], \pt_ob_tlv.tdata [3]);
tran (pt_ob_tlv[2], \pt_ob_tlv.tdata [2]);
tran (pt_ob_tlv[1], \pt_ob_tlv.tdata [1]);
tran (pt_ob_tlv[0], \pt_ob_tlv.tdata [0]);
tran (tlvp_rsm_usr_ob_rdata[105], \tlvp_rsm_usr_ob_rdata.insert );
tran (tlvp_rsm_usr_ob_rdata[104], \tlvp_rsm_usr_ob_rdata.ordern [12]);
tran (tlvp_rsm_usr_ob_rdata[103], \tlvp_rsm_usr_ob_rdata.ordern [11]);
tran (tlvp_rsm_usr_ob_rdata[102], \tlvp_rsm_usr_ob_rdata.ordern [10]);
tran (tlvp_rsm_usr_ob_rdata[101], \tlvp_rsm_usr_ob_rdata.ordern [9]);
tran (tlvp_rsm_usr_ob_rdata[100], \tlvp_rsm_usr_ob_rdata.ordern [8]);
tran (tlvp_rsm_usr_ob_rdata[99], \tlvp_rsm_usr_ob_rdata.ordern [7]);
tran (tlvp_rsm_usr_ob_rdata[98], \tlvp_rsm_usr_ob_rdata.ordern [6]);
tran (tlvp_rsm_usr_ob_rdata[97], \tlvp_rsm_usr_ob_rdata.ordern [5]);
tran (tlvp_rsm_usr_ob_rdata[96], \tlvp_rsm_usr_ob_rdata.ordern [4]);
tran (tlvp_rsm_usr_ob_rdata[95], \tlvp_rsm_usr_ob_rdata.ordern [3]);
tran (tlvp_rsm_usr_ob_rdata[94], \tlvp_rsm_usr_ob_rdata.ordern [2]);
tran (tlvp_rsm_usr_ob_rdata[93], \tlvp_rsm_usr_ob_rdata.ordern [1]);
tran (tlvp_rsm_usr_ob_rdata[92], \tlvp_rsm_usr_ob_rdata.ordern [0]);
tran (tlvp_rsm_usr_ob_rdata[91], \tlvp_rsm_usr_ob_rdata.typen [7]);
tran (tlvp_rsm_usr_ob_rdata[90], \tlvp_rsm_usr_ob_rdata.typen [6]);
tran (tlvp_rsm_usr_ob_rdata[89], \tlvp_rsm_usr_ob_rdata.typen [5]);
tran (tlvp_rsm_usr_ob_rdata[88], \tlvp_rsm_usr_ob_rdata.typen [4]);
tran (tlvp_rsm_usr_ob_rdata[87], \tlvp_rsm_usr_ob_rdata.typen [3]);
tran (tlvp_rsm_usr_ob_rdata[86], \tlvp_rsm_usr_ob_rdata.typen [2]);
tran (tlvp_rsm_usr_ob_rdata[85], \tlvp_rsm_usr_ob_rdata.typen [1]);
tran (tlvp_rsm_usr_ob_rdata[84], \tlvp_rsm_usr_ob_rdata.typen [0]);
tran (tlvp_rsm_usr_ob_rdata[83], \tlvp_rsm_usr_ob_rdata.sot );
tran (tlvp_rsm_usr_ob_rdata[82], \tlvp_rsm_usr_ob_rdata.eot );
tran (tlvp_rsm_usr_ob_rdata[81], \tlvp_rsm_usr_ob_rdata.tlast );
tran (tlvp_rsm_usr_ob_rdata[80], \tlvp_rsm_usr_ob_rdata.tid [0]);
tran (tlvp_rsm_usr_ob_rdata[79], \tlvp_rsm_usr_ob_rdata.tstrb [7]);
tran (tlvp_rsm_usr_ob_rdata[78], \tlvp_rsm_usr_ob_rdata.tstrb [6]);
tran (tlvp_rsm_usr_ob_rdata[77], \tlvp_rsm_usr_ob_rdata.tstrb [5]);
tran (tlvp_rsm_usr_ob_rdata[76], \tlvp_rsm_usr_ob_rdata.tstrb [4]);
tran (tlvp_rsm_usr_ob_rdata[75], \tlvp_rsm_usr_ob_rdata.tstrb [3]);
tran (tlvp_rsm_usr_ob_rdata[74], \tlvp_rsm_usr_ob_rdata.tstrb [2]);
tran (tlvp_rsm_usr_ob_rdata[73], \tlvp_rsm_usr_ob_rdata.tstrb [1]);
tran (tlvp_rsm_usr_ob_rdata[72], \tlvp_rsm_usr_ob_rdata.tstrb [0]);
tran (tlvp_rsm_usr_ob_rdata[71], \tlvp_rsm_usr_ob_rdata.tuser [7]);
tran (tlvp_rsm_usr_ob_rdata[70], \tlvp_rsm_usr_ob_rdata.tuser [6]);
tran (tlvp_rsm_usr_ob_rdata[69], \tlvp_rsm_usr_ob_rdata.tuser [5]);
tran (tlvp_rsm_usr_ob_rdata[68], \tlvp_rsm_usr_ob_rdata.tuser [4]);
tran (tlvp_rsm_usr_ob_rdata[67], \tlvp_rsm_usr_ob_rdata.tuser [3]);
tran (tlvp_rsm_usr_ob_rdata[66], \tlvp_rsm_usr_ob_rdata.tuser [2]);
tran (tlvp_rsm_usr_ob_rdata[65], \tlvp_rsm_usr_ob_rdata.tuser [1]);
tran (tlvp_rsm_usr_ob_rdata[64], \tlvp_rsm_usr_ob_rdata.tuser [0]);
tran (tlvp_rsm_usr_ob_rdata[63], \tlvp_rsm_usr_ob_rdata.tdata [63]);
tran (tlvp_rsm_usr_ob_rdata[62], \tlvp_rsm_usr_ob_rdata.tdata [62]);
tran (tlvp_rsm_usr_ob_rdata[61], \tlvp_rsm_usr_ob_rdata.tdata [61]);
tran (tlvp_rsm_usr_ob_rdata[60], \tlvp_rsm_usr_ob_rdata.tdata [60]);
tran (tlvp_rsm_usr_ob_rdata[59], \tlvp_rsm_usr_ob_rdata.tdata [59]);
tran (tlvp_rsm_usr_ob_rdata[58], \tlvp_rsm_usr_ob_rdata.tdata [58]);
tran (tlvp_rsm_usr_ob_rdata[57], \tlvp_rsm_usr_ob_rdata.tdata [57]);
tran (tlvp_rsm_usr_ob_rdata[56], \tlvp_rsm_usr_ob_rdata.tdata [56]);
tran (tlvp_rsm_usr_ob_rdata[55], \tlvp_rsm_usr_ob_rdata.tdata [55]);
tran (tlvp_rsm_usr_ob_rdata[54], \tlvp_rsm_usr_ob_rdata.tdata [54]);
tran (tlvp_rsm_usr_ob_rdata[53], \tlvp_rsm_usr_ob_rdata.tdata [53]);
tran (tlvp_rsm_usr_ob_rdata[52], \tlvp_rsm_usr_ob_rdata.tdata [52]);
tran (tlvp_rsm_usr_ob_rdata[51], \tlvp_rsm_usr_ob_rdata.tdata [51]);
tran (tlvp_rsm_usr_ob_rdata[50], \tlvp_rsm_usr_ob_rdata.tdata [50]);
tran (tlvp_rsm_usr_ob_rdata[49], \tlvp_rsm_usr_ob_rdata.tdata [49]);
tran (tlvp_rsm_usr_ob_rdata[48], \tlvp_rsm_usr_ob_rdata.tdata [48]);
tran (tlvp_rsm_usr_ob_rdata[47], \tlvp_rsm_usr_ob_rdata.tdata [47]);
tran (tlvp_rsm_usr_ob_rdata[46], \tlvp_rsm_usr_ob_rdata.tdata [46]);
tran (tlvp_rsm_usr_ob_rdata[45], \tlvp_rsm_usr_ob_rdata.tdata [45]);
tran (tlvp_rsm_usr_ob_rdata[44], \tlvp_rsm_usr_ob_rdata.tdata [44]);
tran (tlvp_rsm_usr_ob_rdata[43], \tlvp_rsm_usr_ob_rdata.tdata [43]);
tran (tlvp_rsm_usr_ob_rdata[42], \tlvp_rsm_usr_ob_rdata.tdata [42]);
tran (tlvp_rsm_usr_ob_rdata[41], \tlvp_rsm_usr_ob_rdata.tdata [41]);
tran (tlvp_rsm_usr_ob_rdata[40], \tlvp_rsm_usr_ob_rdata.tdata [40]);
tran (tlvp_rsm_usr_ob_rdata[39], \tlvp_rsm_usr_ob_rdata.tdata [39]);
tran (tlvp_rsm_usr_ob_rdata[38], \tlvp_rsm_usr_ob_rdata.tdata [38]);
tran (tlvp_rsm_usr_ob_rdata[37], \tlvp_rsm_usr_ob_rdata.tdata [37]);
tran (tlvp_rsm_usr_ob_rdata[36], \tlvp_rsm_usr_ob_rdata.tdata [36]);
tran (tlvp_rsm_usr_ob_rdata[35], \tlvp_rsm_usr_ob_rdata.tdata [35]);
tran (tlvp_rsm_usr_ob_rdata[34], \tlvp_rsm_usr_ob_rdata.tdata [34]);
tran (tlvp_rsm_usr_ob_rdata[33], \tlvp_rsm_usr_ob_rdata.tdata [33]);
tran (tlvp_rsm_usr_ob_rdata[32], \tlvp_rsm_usr_ob_rdata.tdata [32]);
tran (tlvp_rsm_usr_ob_rdata[31], \tlvp_rsm_usr_ob_rdata.tdata [31]);
tran (tlvp_rsm_usr_ob_rdata[30], \tlvp_rsm_usr_ob_rdata.tdata [30]);
tran (tlvp_rsm_usr_ob_rdata[29], \tlvp_rsm_usr_ob_rdata.tdata [29]);
tran (tlvp_rsm_usr_ob_rdata[28], \tlvp_rsm_usr_ob_rdata.tdata [28]);
tran (tlvp_rsm_usr_ob_rdata[27], \tlvp_rsm_usr_ob_rdata.tdata [27]);
tran (tlvp_rsm_usr_ob_rdata[26], \tlvp_rsm_usr_ob_rdata.tdata [26]);
tran (tlvp_rsm_usr_ob_rdata[25], \tlvp_rsm_usr_ob_rdata.tdata [25]);
tran (tlvp_rsm_usr_ob_rdata[24], \tlvp_rsm_usr_ob_rdata.tdata [24]);
tran (tlvp_rsm_usr_ob_rdata[23], \tlvp_rsm_usr_ob_rdata.tdata [23]);
tran (tlvp_rsm_usr_ob_rdata[22], \tlvp_rsm_usr_ob_rdata.tdata [22]);
tran (tlvp_rsm_usr_ob_rdata[21], \tlvp_rsm_usr_ob_rdata.tdata [21]);
tran (tlvp_rsm_usr_ob_rdata[20], \tlvp_rsm_usr_ob_rdata.tdata [20]);
tran (tlvp_rsm_usr_ob_rdata[19], \tlvp_rsm_usr_ob_rdata.tdata [19]);
tran (tlvp_rsm_usr_ob_rdata[18], \tlvp_rsm_usr_ob_rdata.tdata [18]);
tran (tlvp_rsm_usr_ob_rdata[17], \tlvp_rsm_usr_ob_rdata.tdata [17]);
tran (tlvp_rsm_usr_ob_rdata[16], \tlvp_rsm_usr_ob_rdata.tdata [16]);
tran (tlvp_rsm_usr_ob_rdata[15], \tlvp_rsm_usr_ob_rdata.tdata [15]);
tran (tlvp_rsm_usr_ob_rdata[14], \tlvp_rsm_usr_ob_rdata.tdata [14]);
tran (tlvp_rsm_usr_ob_rdata[13], \tlvp_rsm_usr_ob_rdata.tdata [13]);
tran (tlvp_rsm_usr_ob_rdata[12], \tlvp_rsm_usr_ob_rdata.tdata [12]);
tran (tlvp_rsm_usr_ob_rdata[11], \tlvp_rsm_usr_ob_rdata.tdata [11]);
tran (tlvp_rsm_usr_ob_rdata[10], \tlvp_rsm_usr_ob_rdata.tdata [10]);
tran (tlvp_rsm_usr_ob_rdata[9], \tlvp_rsm_usr_ob_rdata.tdata [9]);
tran (tlvp_rsm_usr_ob_rdata[8], \tlvp_rsm_usr_ob_rdata.tdata [8]);
tran (tlvp_rsm_usr_ob_rdata[7], \tlvp_rsm_usr_ob_rdata.tdata [7]);
tran (tlvp_rsm_usr_ob_rdata[6], \tlvp_rsm_usr_ob_rdata.tdata [6]);
tran (tlvp_rsm_usr_ob_rdata[5], \tlvp_rsm_usr_ob_rdata.tdata [5]);
tran (tlvp_rsm_usr_ob_rdata[4], \tlvp_rsm_usr_ob_rdata.tdata [4]);
tran (tlvp_rsm_usr_ob_rdata[3], \tlvp_rsm_usr_ob_rdata.tdata [3]);
tran (tlvp_rsm_usr_ob_rdata[2], \tlvp_rsm_usr_ob_rdata.tdata [2]);
tran (tlvp_rsm_usr_ob_rdata[1], \tlvp_rsm_usr_ob_rdata.tdata [1]);
tran (tlvp_rsm_usr_ob_rdata[0], \tlvp_rsm_usr_ob_rdata.tdata [0]);
tran (tlvp_rsm_ob_datain[0], \tlvp_rsm_ob_datain.tdata [0]);
tran (tlvp_rsm_ob_datain[1], \tlvp_rsm_ob_datain.tdata [1]);
tran (tlvp_rsm_ob_datain[2], \tlvp_rsm_ob_datain.tdata [2]);
tran (tlvp_rsm_ob_datain[3], \tlvp_rsm_ob_datain.tdata [3]);
tran (tlvp_rsm_ob_datain[4], \tlvp_rsm_ob_datain.tdata [4]);
tran (tlvp_rsm_ob_datain[5], \tlvp_rsm_ob_datain.tdata [5]);
tran (tlvp_rsm_ob_datain[6], \tlvp_rsm_ob_datain.tdata [6]);
tran (tlvp_rsm_ob_datain[7], \tlvp_rsm_ob_datain.tdata [7]);
tran (tlvp_rsm_ob_datain[8], \tlvp_rsm_ob_datain.tdata [8]);
tran (tlvp_rsm_ob_datain[9], \tlvp_rsm_ob_datain.tdata [9]);
tran (tlvp_rsm_ob_datain[10], \tlvp_rsm_ob_datain.tdata [10]);
tran (tlvp_rsm_ob_datain[11], \tlvp_rsm_ob_datain.tdata [11]);
tran (tlvp_rsm_ob_datain[12], \tlvp_rsm_ob_datain.tdata [12]);
tran (tlvp_rsm_ob_datain[13], \tlvp_rsm_ob_datain.tdata [13]);
tran (tlvp_rsm_ob_datain[14], \tlvp_rsm_ob_datain.tdata [14]);
tran (tlvp_rsm_ob_datain[15], \tlvp_rsm_ob_datain.tdata [15]);
tran (tlvp_rsm_ob_datain[16], \tlvp_rsm_ob_datain.tdata [16]);
tran (tlvp_rsm_ob_datain[17], \tlvp_rsm_ob_datain.tdata [17]);
tran (tlvp_rsm_ob_datain[18], \tlvp_rsm_ob_datain.tdata [18]);
tran (tlvp_rsm_ob_datain[19], \tlvp_rsm_ob_datain.tdata [19]);
tran (tlvp_rsm_ob_datain[20], \tlvp_rsm_ob_datain.tdata [20]);
tran (tlvp_rsm_ob_datain[21], \tlvp_rsm_ob_datain.tdata [21]);
tran (tlvp_rsm_ob_datain[22], \tlvp_rsm_ob_datain.tdata [22]);
tran (tlvp_rsm_ob_datain[23], \tlvp_rsm_ob_datain.tdata [23]);
tran (tlvp_rsm_ob_datain[24], \tlvp_rsm_ob_datain.tdata [24]);
tran (tlvp_rsm_ob_datain[25], \tlvp_rsm_ob_datain.tdata [25]);
tran (tlvp_rsm_ob_datain[26], \tlvp_rsm_ob_datain.tdata [26]);
tran (tlvp_rsm_ob_datain[27], \tlvp_rsm_ob_datain.tdata [27]);
tran (tlvp_rsm_ob_datain[28], \tlvp_rsm_ob_datain.tdata [28]);
tran (tlvp_rsm_ob_datain[29], \tlvp_rsm_ob_datain.tdata [29]);
tran (tlvp_rsm_ob_datain[30], \tlvp_rsm_ob_datain.tdata [30]);
tran (tlvp_rsm_ob_datain[31], \tlvp_rsm_ob_datain.tdata [31]);
tran (tlvp_rsm_ob_datain[32], \tlvp_rsm_ob_datain.tdata [32]);
tran (tlvp_rsm_ob_datain[33], \tlvp_rsm_ob_datain.tdata [33]);
tran (tlvp_rsm_ob_datain[34], \tlvp_rsm_ob_datain.tdata [34]);
tran (tlvp_rsm_ob_datain[35], \tlvp_rsm_ob_datain.tdata [35]);
tran (tlvp_rsm_ob_datain[36], \tlvp_rsm_ob_datain.tdata [36]);
tran (tlvp_rsm_ob_datain[37], \tlvp_rsm_ob_datain.tdata [37]);
tran (tlvp_rsm_ob_datain[38], \tlvp_rsm_ob_datain.tdata [38]);
tran (tlvp_rsm_ob_datain[39], \tlvp_rsm_ob_datain.tdata [39]);
tran (tlvp_rsm_ob_datain[40], \tlvp_rsm_ob_datain.tdata [40]);
tran (tlvp_rsm_ob_datain[41], \tlvp_rsm_ob_datain.tdata [41]);
tran (tlvp_rsm_ob_datain[42], \tlvp_rsm_ob_datain.tdata [42]);
tran (tlvp_rsm_ob_datain[43], \tlvp_rsm_ob_datain.tdata [43]);
tran (tlvp_rsm_ob_datain[44], \tlvp_rsm_ob_datain.tdata [44]);
tran (tlvp_rsm_ob_datain[45], \tlvp_rsm_ob_datain.tdata [45]);
tran (tlvp_rsm_ob_datain[46], \tlvp_rsm_ob_datain.tdata [46]);
tran (tlvp_rsm_ob_datain[47], \tlvp_rsm_ob_datain.tdata [47]);
tran (tlvp_rsm_ob_datain[48], \tlvp_rsm_ob_datain.tdata [48]);
tran (tlvp_rsm_ob_datain[49], \tlvp_rsm_ob_datain.tdata [49]);
tran (tlvp_rsm_ob_datain[50], \tlvp_rsm_ob_datain.tdata [50]);
tran (tlvp_rsm_ob_datain[51], \tlvp_rsm_ob_datain.tdata [51]);
tran (tlvp_rsm_ob_datain[52], \tlvp_rsm_ob_datain.tdata [52]);
tran (tlvp_rsm_ob_datain[53], \tlvp_rsm_ob_datain.tdata [53]);
tran (tlvp_rsm_ob_datain[54], \tlvp_rsm_ob_datain.tdata [54]);
tran (tlvp_rsm_ob_datain[55], \tlvp_rsm_ob_datain.tdata [55]);
tran (tlvp_rsm_ob_datain[56], \tlvp_rsm_ob_datain.tdata [56]);
tran (tlvp_rsm_ob_datain[57], \tlvp_rsm_ob_datain.tdata [57]);
tran (tlvp_rsm_ob_datain[58], \tlvp_rsm_ob_datain.tdata [58]);
tran (tlvp_rsm_ob_datain[59], \tlvp_rsm_ob_datain.tdata [59]);
tran (tlvp_rsm_ob_datain[60], \tlvp_rsm_ob_datain.tdata [60]);
tran (tlvp_rsm_ob_datain[61], \tlvp_rsm_ob_datain.tdata [61]);
tran (tlvp_rsm_ob_datain[62], \tlvp_rsm_ob_datain.tdata [62]);
tran (tlvp_rsm_ob_datain[63], \tlvp_rsm_ob_datain.tdata [63]);
tran (tlvp_rsm_ob_datain[64], \tlvp_rsm_ob_datain.tuser [0]);
tran (tlvp_rsm_ob_datain[65], \tlvp_rsm_ob_datain.tuser [1]);
tran (tlvp_rsm_ob_datain[66], \tlvp_rsm_ob_datain.tuser [2]);
tran (tlvp_rsm_ob_datain[67], \tlvp_rsm_ob_datain.tuser [3]);
tran (tlvp_rsm_ob_datain[68], \tlvp_rsm_ob_datain.tuser [4]);
tran (tlvp_rsm_ob_datain[69], \tlvp_rsm_ob_datain.tuser [5]);
tran (tlvp_rsm_ob_datain[70], \tlvp_rsm_ob_datain.tuser [6]);
tran (tlvp_rsm_ob_datain[71], \tlvp_rsm_ob_datain.tuser [7]);
tran (tlvp_rsm_ob_datain[72], \tlvp_rsm_ob_datain.tstrb [0]);
tran (tlvp_rsm_ob_datain[73], \tlvp_rsm_ob_datain.tstrb [1]);
tran (tlvp_rsm_ob_datain[74], \tlvp_rsm_ob_datain.tstrb [2]);
tran (tlvp_rsm_ob_datain[75], \tlvp_rsm_ob_datain.tstrb [3]);
tran (tlvp_rsm_ob_datain[76], \tlvp_rsm_ob_datain.tstrb [4]);
tran (tlvp_rsm_ob_datain[77], \tlvp_rsm_ob_datain.tstrb [5]);
tran (tlvp_rsm_ob_datain[78], \tlvp_rsm_ob_datain.tstrb [6]);
tran (tlvp_rsm_ob_datain[79], \tlvp_rsm_ob_datain.tstrb [7]);
tran (tlvp_rsm_ob_datain[80], \tlvp_rsm_ob_datain.tid [0]);
tran (tlvp_rsm_ob_datain[81], \tlvp_rsm_ob_datain.tlast );
tran (tlvp_rsm_ob_datain[82], \tlvp_rsm_ob_datain.eot );
tran (tlvp_rsm_ob_datain[83], \tlvp_rsm_ob_datain.sot );
tran (tlvp_rsm_ob_datain[84], \tlvp_rsm_ob_datain.typen [0]);
tran (tlvp_rsm_ob_datain[85], \tlvp_rsm_ob_datain.typen [1]);
tran (tlvp_rsm_ob_datain[86], \tlvp_rsm_ob_datain.typen [2]);
tran (tlvp_rsm_ob_datain[87], \tlvp_rsm_ob_datain.typen [3]);
tran (tlvp_rsm_ob_datain[88], \tlvp_rsm_ob_datain.typen [4]);
tran (tlvp_rsm_ob_datain[89], \tlvp_rsm_ob_datain.typen [5]);
tran (tlvp_rsm_ob_datain[90], \tlvp_rsm_ob_datain.typen [6]);
tran (tlvp_rsm_ob_datain[91], \tlvp_rsm_ob_datain.typen [7]);
tran (tlvp_rsm_ob_datain[92], \tlvp_rsm_ob_datain.ordern [0]);
tran (tlvp_rsm_ob_datain[93], \tlvp_rsm_ob_datain.ordern [1]);
tran (tlvp_rsm_ob_datain[94], \tlvp_rsm_ob_datain.ordern [2]);
tran (tlvp_rsm_ob_datain[95], \tlvp_rsm_ob_datain.ordern [3]);
tran (tlvp_rsm_ob_datain[96], \tlvp_rsm_ob_datain.ordern [4]);
tran (tlvp_rsm_ob_datain[97], \tlvp_rsm_ob_datain.ordern [5]);
tran (tlvp_rsm_ob_datain[98], \tlvp_rsm_ob_datain.ordern [6]);
tran (tlvp_rsm_ob_datain[99], \tlvp_rsm_ob_datain.ordern [7]);
tran (tlvp_rsm_ob_datain[100], \tlvp_rsm_ob_datain.ordern [8]);
tran (tlvp_rsm_ob_datain[101], \tlvp_rsm_ob_datain.ordern [9]);
tran (tlvp_rsm_ob_datain[102], \tlvp_rsm_ob_datain.ordern [10]);
tran (tlvp_rsm_ob_datain[103], \tlvp_rsm_ob_datain.ordern [11]);
tran (tlvp_rsm_ob_datain[104], \tlvp_rsm_ob_datain.ordern [12]);
tran (tlvp_rsm_ob_datain[105], \tlvp_rsm_ob_datain.insert );
tran (tlvp_rsm_pt_tlv[0], \tlvp_rsm_pt_tlv.tdata [0]);
tran (tlvp_rsm_pt_tlv[1], \tlvp_rsm_pt_tlv.tdata [1]);
tran (tlvp_rsm_pt_tlv[2], \tlvp_rsm_pt_tlv.tdata [2]);
tran (tlvp_rsm_pt_tlv[3], \tlvp_rsm_pt_tlv.tdata [3]);
tran (tlvp_rsm_pt_tlv[4], \tlvp_rsm_pt_tlv.tdata [4]);
tran (tlvp_rsm_pt_tlv[5], \tlvp_rsm_pt_tlv.tdata [5]);
tran (tlvp_rsm_pt_tlv[6], \tlvp_rsm_pt_tlv.tdata [6]);
tran (tlvp_rsm_pt_tlv[7], \tlvp_rsm_pt_tlv.tdata [7]);
tran (tlvp_rsm_pt_tlv[8], \tlvp_rsm_pt_tlv.tdata [8]);
tran (tlvp_rsm_pt_tlv[9], \tlvp_rsm_pt_tlv.tdata [9]);
tran (tlvp_rsm_pt_tlv[10], \tlvp_rsm_pt_tlv.tdata [10]);
tran (tlvp_rsm_pt_tlv[11], \tlvp_rsm_pt_tlv.tdata [11]);
tran (tlvp_rsm_pt_tlv[12], \tlvp_rsm_pt_tlv.tdata [12]);
tran (tlvp_rsm_pt_tlv[13], \tlvp_rsm_pt_tlv.tdata [13]);
tran (tlvp_rsm_pt_tlv[14], \tlvp_rsm_pt_tlv.tdata [14]);
tran (tlvp_rsm_pt_tlv[15], \tlvp_rsm_pt_tlv.tdata [15]);
tran (tlvp_rsm_pt_tlv[16], \tlvp_rsm_pt_tlv.tdata [16]);
tran (tlvp_rsm_pt_tlv[17], \tlvp_rsm_pt_tlv.tdata [17]);
tran (tlvp_rsm_pt_tlv[18], \tlvp_rsm_pt_tlv.tdata [18]);
tran (tlvp_rsm_pt_tlv[19], \tlvp_rsm_pt_tlv.tdata [19]);
tran (tlvp_rsm_pt_tlv[20], \tlvp_rsm_pt_tlv.tdata [20]);
tran (tlvp_rsm_pt_tlv[21], \tlvp_rsm_pt_tlv.tdata [21]);
tran (tlvp_rsm_pt_tlv[22], \tlvp_rsm_pt_tlv.tdata [22]);
tran (tlvp_rsm_pt_tlv[23], \tlvp_rsm_pt_tlv.tdata [23]);
tran (tlvp_rsm_pt_tlv[24], \tlvp_rsm_pt_tlv.tdata [24]);
tran (tlvp_rsm_pt_tlv[25], \tlvp_rsm_pt_tlv.tdata [25]);
tran (tlvp_rsm_pt_tlv[26], \tlvp_rsm_pt_tlv.tdata [26]);
tran (tlvp_rsm_pt_tlv[27], \tlvp_rsm_pt_tlv.tdata [27]);
tran (tlvp_rsm_pt_tlv[28], \tlvp_rsm_pt_tlv.tdata [28]);
tran (tlvp_rsm_pt_tlv[29], \tlvp_rsm_pt_tlv.tdata [29]);
tran (tlvp_rsm_pt_tlv[30], \tlvp_rsm_pt_tlv.tdata [30]);
tran (tlvp_rsm_pt_tlv[31], \tlvp_rsm_pt_tlv.tdata [31]);
tran (tlvp_rsm_pt_tlv[32], \tlvp_rsm_pt_tlv.tdata [32]);
tran (tlvp_rsm_pt_tlv[33], \tlvp_rsm_pt_tlv.tdata [33]);
tran (tlvp_rsm_pt_tlv[34], \tlvp_rsm_pt_tlv.tdata [34]);
tran (tlvp_rsm_pt_tlv[35], \tlvp_rsm_pt_tlv.tdata [35]);
tran (tlvp_rsm_pt_tlv[36], \tlvp_rsm_pt_tlv.tdata [36]);
tran (tlvp_rsm_pt_tlv[37], \tlvp_rsm_pt_tlv.tdata [37]);
tran (tlvp_rsm_pt_tlv[38], \tlvp_rsm_pt_tlv.tdata [38]);
tran (tlvp_rsm_pt_tlv[39], \tlvp_rsm_pt_tlv.tdata [39]);
tran (tlvp_rsm_pt_tlv[40], \tlvp_rsm_pt_tlv.tdata [40]);
tran (tlvp_rsm_pt_tlv[41], \tlvp_rsm_pt_tlv.tdata [41]);
tran (tlvp_rsm_pt_tlv[42], \tlvp_rsm_pt_tlv.tdata [42]);
tran (tlvp_rsm_pt_tlv[43], \tlvp_rsm_pt_tlv.tdata [43]);
tran (tlvp_rsm_pt_tlv[44], \tlvp_rsm_pt_tlv.tdata [44]);
tran (tlvp_rsm_pt_tlv[45], \tlvp_rsm_pt_tlv.tdata [45]);
tran (tlvp_rsm_pt_tlv[46], \tlvp_rsm_pt_tlv.tdata [46]);
tran (tlvp_rsm_pt_tlv[47], \tlvp_rsm_pt_tlv.tdata [47]);
tran (tlvp_rsm_pt_tlv[48], \tlvp_rsm_pt_tlv.tdata [48]);
tran (tlvp_rsm_pt_tlv[49], \tlvp_rsm_pt_tlv.tdata [49]);
tran (tlvp_rsm_pt_tlv[50], \tlvp_rsm_pt_tlv.tdata [50]);
tran (tlvp_rsm_pt_tlv[51], \tlvp_rsm_pt_tlv.tdata [51]);
tran (tlvp_rsm_pt_tlv[52], \tlvp_rsm_pt_tlv.tdata [52]);
tran (tlvp_rsm_pt_tlv[53], \tlvp_rsm_pt_tlv.tdata [53]);
tran (tlvp_rsm_pt_tlv[54], \tlvp_rsm_pt_tlv.tdata [54]);
tran (tlvp_rsm_pt_tlv[55], \tlvp_rsm_pt_tlv.tdata [55]);
tran (tlvp_rsm_pt_tlv[56], \tlvp_rsm_pt_tlv.tdata [56]);
tran (tlvp_rsm_pt_tlv[57], \tlvp_rsm_pt_tlv.tdata [57]);
tran (tlvp_rsm_pt_tlv[58], \tlvp_rsm_pt_tlv.tdata [58]);
tran (tlvp_rsm_pt_tlv[59], \tlvp_rsm_pt_tlv.tdata [59]);
tran (tlvp_rsm_pt_tlv[60], \tlvp_rsm_pt_tlv.tdata [60]);
tran (tlvp_rsm_pt_tlv[61], \tlvp_rsm_pt_tlv.tdata [61]);
tran (tlvp_rsm_pt_tlv[62], \tlvp_rsm_pt_tlv.tdata [62]);
tran (tlvp_rsm_pt_tlv[63], \tlvp_rsm_pt_tlv.tdata [63]);
tran (tlvp_rsm_pt_tlv[64], \tlvp_rsm_pt_tlv.tuser [0]);
tran (tlvp_rsm_pt_tlv[65], \tlvp_rsm_pt_tlv.tuser [1]);
tran (tlvp_rsm_pt_tlv[66], \tlvp_rsm_pt_tlv.tuser [2]);
tran (tlvp_rsm_pt_tlv[67], \tlvp_rsm_pt_tlv.tuser [3]);
tran (tlvp_rsm_pt_tlv[68], \tlvp_rsm_pt_tlv.tuser [4]);
tran (tlvp_rsm_pt_tlv[69], \tlvp_rsm_pt_tlv.tuser [5]);
tran (tlvp_rsm_pt_tlv[70], \tlvp_rsm_pt_tlv.tuser [6]);
tran (tlvp_rsm_pt_tlv[71], \tlvp_rsm_pt_tlv.tuser [7]);
tran (tlvp_rsm_pt_tlv[72], \tlvp_rsm_pt_tlv.tstrb [0]);
tran (tlvp_rsm_pt_tlv[73], \tlvp_rsm_pt_tlv.tstrb [1]);
tran (tlvp_rsm_pt_tlv[74], \tlvp_rsm_pt_tlv.tstrb [2]);
tran (tlvp_rsm_pt_tlv[75], \tlvp_rsm_pt_tlv.tstrb [3]);
tran (tlvp_rsm_pt_tlv[76], \tlvp_rsm_pt_tlv.tstrb [4]);
tran (tlvp_rsm_pt_tlv[77], \tlvp_rsm_pt_tlv.tstrb [5]);
tran (tlvp_rsm_pt_tlv[78], \tlvp_rsm_pt_tlv.tstrb [6]);
tran (tlvp_rsm_pt_tlv[79], \tlvp_rsm_pt_tlv.tstrb [7]);
tran (tlvp_rsm_pt_tlv[80], \tlvp_rsm_pt_tlv.tid [0]);
tran (tlvp_rsm_pt_tlv[81], \tlvp_rsm_pt_tlv.tlast );
tran (tlvp_rsm_pt_tlv[82], \tlvp_rsm_pt_tlv.eot );
tran (tlvp_rsm_pt_tlv[83], \tlvp_rsm_pt_tlv.sot );
tran (tlvp_rsm_pt_tlv[84], \tlvp_rsm_pt_tlv.typen [0]);
tran (tlvp_rsm_pt_tlv[85], \tlvp_rsm_pt_tlv.typen [1]);
tran (tlvp_rsm_pt_tlv[86], \tlvp_rsm_pt_tlv.typen [2]);
tran (tlvp_rsm_pt_tlv[87], \tlvp_rsm_pt_tlv.typen [3]);
tran (tlvp_rsm_pt_tlv[88], \tlvp_rsm_pt_tlv.typen [4]);
tran (tlvp_rsm_pt_tlv[89], \tlvp_rsm_pt_tlv.typen [5]);
tran (tlvp_rsm_pt_tlv[90], \tlvp_rsm_pt_tlv.typen [6]);
tran (tlvp_rsm_pt_tlv[91], \tlvp_rsm_pt_tlv.typen [7]);
tran (tlvp_rsm_pt_tlv[92], \tlvp_rsm_pt_tlv.ordern [0]);
tran (tlvp_rsm_pt_tlv[93], \tlvp_rsm_pt_tlv.ordern [1]);
tran (tlvp_rsm_pt_tlv[94], \tlvp_rsm_pt_tlv.ordern [2]);
tran (tlvp_rsm_pt_tlv[95], \tlvp_rsm_pt_tlv.ordern [3]);
tran (tlvp_rsm_pt_tlv[96], \tlvp_rsm_pt_tlv.ordern [4]);
tran (tlvp_rsm_pt_tlv[97], \tlvp_rsm_pt_tlv.ordern [5]);
tran (tlvp_rsm_pt_tlv[98], \tlvp_rsm_pt_tlv.ordern [6]);
tran (tlvp_rsm_pt_tlv[99], \tlvp_rsm_pt_tlv.ordern [7]);
tran (tlvp_rsm_pt_tlv[100], \tlvp_rsm_pt_tlv.ordern [8]);
tran (tlvp_rsm_pt_tlv[101], \tlvp_rsm_pt_tlv.ordern [9]);
tran (tlvp_rsm_pt_tlv[102], \tlvp_rsm_pt_tlv.ordern [10]);
tran (tlvp_rsm_pt_tlv[103], \tlvp_rsm_pt_tlv.ordern [11]);
tran (tlvp_rsm_pt_tlv[104], \tlvp_rsm_pt_tlv.ordern [12]);
tran (tlvp_rsm_pt_tlv[105], \tlvp_rsm_pt_tlv.insert );
tran (tlvp_rsm_usr_ob_tlv[0], \tlvp_rsm_usr_ob_tlv.tdata [0]);
tran (tlvp_rsm_usr_ob_tlv[1], \tlvp_rsm_usr_ob_tlv.tdata [1]);
tran (tlvp_rsm_usr_ob_tlv[2], \tlvp_rsm_usr_ob_tlv.tdata [2]);
tran (tlvp_rsm_usr_ob_tlv[3], \tlvp_rsm_usr_ob_tlv.tdata [3]);
tran (tlvp_rsm_usr_ob_tlv[4], \tlvp_rsm_usr_ob_tlv.tdata [4]);
tran (tlvp_rsm_usr_ob_tlv[5], \tlvp_rsm_usr_ob_tlv.tdata [5]);
tran (tlvp_rsm_usr_ob_tlv[6], \tlvp_rsm_usr_ob_tlv.tdata [6]);
tran (tlvp_rsm_usr_ob_tlv[7], \tlvp_rsm_usr_ob_tlv.tdata [7]);
tran (tlvp_rsm_usr_ob_tlv[8], \tlvp_rsm_usr_ob_tlv.tdata [8]);
tran (tlvp_rsm_usr_ob_tlv[9], \tlvp_rsm_usr_ob_tlv.tdata [9]);
tran (tlvp_rsm_usr_ob_tlv[10], \tlvp_rsm_usr_ob_tlv.tdata [10]);
tran (tlvp_rsm_usr_ob_tlv[11], \tlvp_rsm_usr_ob_tlv.tdata [11]);
tran (tlvp_rsm_usr_ob_tlv[12], \tlvp_rsm_usr_ob_tlv.tdata [12]);
tran (tlvp_rsm_usr_ob_tlv[13], \tlvp_rsm_usr_ob_tlv.tdata [13]);
tran (tlvp_rsm_usr_ob_tlv[14], \tlvp_rsm_usr_ob_tlv.tdata [14]);
tran (tlvp_rsm_usr_ob_tlv[15], \tlvp_rsm_usr_ob_tlv.tdata [15]);
tran (tlvp_rsm_usr_ob_tlv[16], \tlvp_rsm_usr_ob_tlv.tdata [16]);
tran (tlvp_rsm_usr_ob_tlv[17], \tlvp_rsm_usr_ob_tlv.tdata [17]);
tran (tlvp_rsm_usr_ob_tlv[18], \tlvp_rsm_usr_ob_tlv.tdata [18]);
tran (tlvp_rsm_usr_ob_tlv[19], \tlvp_rsm_usr_ob_tlv.tdata [19]);
tran (tlvp_rsm_usr_ob_tlv[20], \tlvp_rsm_usr_ob_tlv.tdata [20]);
tran (tlvp_rsm_usr_ob_tlv[21], \tlvp_rsm_usr_ob_tlv.tdata [21]);
tran (tlvp_rsm_usr_ob_tlv[22], \tlvp_rsm_usr_ob_tlv.tdata [22]);
tran (tlvp_rsm_usr_ob_tlv[23], \tlvp_rsm_usr_ob_tlv.tdata [23]);
tran (tlvp_rsm_usr_ob_tlv[24], \tlvp_rsm_usr_ob_tlv.tdata [24]);
tran (tlvp_rsm_usr_ob_tlv[25], \tlvp_rsm_usr_ob_tlv.tdata [25]);
tran (tlvp_rsm_usr_ob_tlv[26], \tlvp_rsm_usr_ob_tlv.tdata [26]);
tran (tlvp_rsm_usr_ob_tlv[27], \tlvp_rsm_usr_ob_tlv.tdata [27]);
tran (tlvp_rsm_usr_ob_tlv[28], \tlvp_rsm_usr_ob_tlv.tdata [28]);
tran (tlvp_rsm_usr_ob_tlv[29], \tlvp_rsm_usr_ob_tlv.tdata [29]);
tran (tlvp_rsm_usr_ob_tlv[30], \tlvp_rsm_usr_ob_tlv.tdata [30]);
tran (tlvp_rsm_usr_ob_tlv[31], \tlvp_rsm_usr_ob_tlv.tdata [31]);
tran (tlvp_rsm_usr_ob_tlv[32], \tlvp_rsm_usr_ob_tlv.tdata [32]);
tran (tlvp_rsm_usr_ob_tlv[33], \tlvp_rsm_usr_ob_tlv.tdata [33]);
tran (tlvp_rsm_usr_ob_tlv[34], \tlvp_rsm_usr_ob_tlv.tdata [34]);
tran (tlvp_rsm_usr_ob_tlv[35], \tlvp_rsm_usr_ob_tlv.tdata [35]);
tran (tlvp_rsm_usr_ob_tlv[36], \tlvp_rsm_usr_ob_tlv.tdata [36]);
tran (tlvp_rsm_usr_ob_tlv[37], \tlvp_rsm_usr_ob_tlv.tdata [37]);
tran (tlvp_rsm_usr_ob_tlv[38], \tlvp_rsm_usr_ob_tlv.tdata [38]);
tran (tlvp_rsm_usr_ob_tlv[39], \tlvp_rsm_usr_ob_tlv.tdata [39]);
tran (tlvp_rsm_usr_ob_tlv[40], \tlvp_rsm_usr_ob_tlv.tdata [40]);
tran (tlvp_rsm_usr_ob_tlv[41], \tlvp_rsm_usr_ob_tlv.tdata [41]);
tran (tlvp_rsm_usr_ob_tlv[42], \tlvp_rsm_usr_ob_tlv.tdata [42]);
tran (tlvp_rsm_usr_ob_tlv[43], \tlvp_rsm_usr_ob_tlv.tdata [43]);
tran (tlvp_rsm_usr_ob_tlv[44], \tlvp_rsm_usr_ob_tlv.tdata [44]);
tran (tlvp_rsm_usr_ob_tlv[45], \tlvp_rsm_usr_ob_tlv.tdata [45]);
tran (tlvp_rsm_usr_ob_tlv[46], \tlvp_rsm_usr_ob_tlv.tdata [46]);
tran (tlvp_rsm_usr_ob_tlv[47], \tlvp_rsm_usr_ob_tlv.tdata [47]);
tran (tlvp_rsm_usr_ob_tlv[48], \tlvp_rsm_usr_ob_tlv.tdata [48]);
tran (tlvp_rsm_usr_ob_tlv[49], \tlvp_rsm_usr_ob_tlv.tdata [49]);
tran (tlvp_rsm_usr_ob_tlv[50], \tlvp_rsm_usr_ob_tlv.tdata [50]);
tran (tlvp_rsm_usr_ob_tlv[51], \tlvp_rsm_usr_ob_tlv.tdata [51]);
tran (tlvp_rsm_usr_ob_tlv[52], \tlvp_rsm_usr_ob_tlv.tdata [52]);
tran (tlvp_rsm_usr_ob_tlv[53], \tlvp_rsm_usr_ob_tlv.tdata [53]);
tran (tlvp_rsm_usr_ob_tlv[54], \tlvp_rsm_usr_ob_tlv.tdata [54]);
tran (tlvp_rsm_usr_ob_tlv[55], \tlvp_rsm_usr_ob_tlv.tdata [55]);
tran (tlvp_rsm_usr_ob_tlv[56], \tlvp_rsm_usr_ob_tlv.tdata [56]);
tran (tlvp_rsm_usr_ob_tlv[57], \tlvp_rsm_usr_ob_tlv.tdata [57]);
tran (tlvp_rsm_usr_ob_tlv[58], \tlvp_rsm_usr_ob_tlv.tdata [58]);
tran (tlvp_rsm_usr_ob_tlv[59], \tlvp_rsm_usr_ob_tlv.tdata [59]);
tran (tlvp_rsm_usr_ob_tlv[60], \tlvp_rsm_usr_ob_tlv.tdata [60]);
tran (tlvp_rsm_usr_ob_tlv[61], \tlvp_rsm_usr_ob_tlv.tdata [61]);
tran (tlvp_rsm_usr_ob_tlv[62], \tlvp_rsm_usr_ob_tlv.tdata [62]);
tran (tlvp_rsm_usr_ob_tlv[63], \tlvp_rsm_usr_ob_tlv.tdata [63]);
tran (tlvp_rsm_usr_ob_tlv[64], \tlvp_rsm_usr_ob_tlv.tuser [0]);
tran (tlvp_rsm_usr_ob_tlv[65], \tlvp_rsm_usr_ob_tlv.tuser [1]);
tran (tlvp_rsm_usr_ob_tlv[66], \tlvp_rsm_usr_ob_tlv.tuser [2]);
tran (tlvp_rsm_usr_ob_tlv[67], \tlvp_rsm_usr_ob_tlv.tuser [3]);
tran (tlvp_rsm_usr_ob_tlv[68], \tlvp_rsm_usr_ob_tlv.tuser [4]);
tran (tlvp_rsm_usr_ob_tlv[69], \tlvp_rsm_usr_ob_tlv.tuser [5]);
tran (tlvp_rsm_usr_ob_tlv[70], \tlvp_rsm_usr_ob_tlv.tuser [6]);
tran (tlvp_rsm_usr_ob_tlv[71], \tlvp_rsm_usr_ob_tlv.tuser [7]);
tran (tlvp_rsm_usr_ob_tlv[72], \tlvp_rsm_usr_ob_tlv.tstrb [0]);
tran (tlvp_rsm_usr_ob_tlv[73], \tlvp_rsm_usr_ob_tlv.tstrb [1]);
tran (tlvp_rsm_usr_ob_tlv[74], \tlvp_rsm_usr_ob_tlv.tstrb [2]);
tran (tlvp_rsm_usr_ob_tlv[75], \tlvp_rsm_usr_ob_tlv.tstrb [3]);
tran (tlvp_rsm_usr_ob_tlv[76], \tlvp_rsm_usr_ob_tlv.tstrb [4]);
tran (tlvp_rsm_usr_ob_tlv[77], \tlvp_rsm_usr_ob_tlv.tstrb [5]);
tran (tlvp_rsm_usr_ob_tlv[78], \tlvp_rsm_usr_ob_tlv.tstrb [6]);
tran (tlvp_rsm_usr_ob_tlv[79], \tlvp_rsm_usr_ob_tlv.tstrb [7]);
tran (tlvp_rsm_usr_ob_tlv[80], \tlvp_rsm_usr_ob_tlv.tid [0]);
tran (tlvp_rsm_usr_ob_tlv[81], \tlvp_rsm_usr_ob_tlv.tlast );
tran (tlvp_rsm_usr_ob_tlv[82], \tlvp_rsm_usr_ob_tlv.eot );
tran (tlvp_rsm_usr_ob_tlv[83], \tlvp_rsm_usr_ob_tlv.sot );
tran (tlvp_rsm_usr_ob_tlv[84], \tlvp_rsm_usr_ob_tlv.typen [0]);
tran (tlvp_rsm_usr_ob_tlv[85], \tlvp_rsm_usr_ob_tlv.typen [1]);
tran (tlvp_rsm_usr_ob_tlv[86], \tlvp_rsm_usr_ob_tlv.typen [2]);
tran (tlvp_rsm_usr_ob_tlv[87], \tlvp_rsm_usr_ob_tlv.typen [3]);
tran (tlvp_rsm_usr_ob_tlv[88], \tlvp_rsm_usr_ob_tlv.typen [4]);
tran (tlvp_rsm_usr_ob_tlv[89], \tlvp_rsm_usr_ob_tlv.typen [5]);
tran (tlvp_rsm_usr_ob_tlv[90], \tlvp_rsm_usr_ob_tlv.typen [6]);
tran (tlvp_rsm_usr_ob_tlv[91], \tlvp_rsm_usr_ob_tlv.typen [7]);
tran (tlvp_rsm_usr_ob_tlv[92], \tlvp_rsm_usr_ob_tlv.ordern [0]);
tran (tlvp_rsm_usr_ob_tlv[93], \tlvp_rsm_usr_ob_tlv.ordern [1]);
tran (tlvp_rsm_usr_ob_tlv[94], \tlvp_rsm_usr_ob_tlv.ordern [2]);
tran (tlvp_rsm_usr_ob_tlv[95], \tlvp_rsm_usr_ob_tlv.ordern [3]);
tran (tlvp_rsm_usr_ob_tlv[96], \tlvp_rsm_usr_ob_tlv.ordern [4]);
tran (tlvp_rsm_usr_ob_tlv[97], \tlvp_rsm_usr_ob_tlv.ordern [5]);
tran (tlvp_rsm_usr_ob_tlv[98], \tlvp_rsm_usr_ob_tlv.ordern [6]);
tran (tlvp_rsm_usr_ob_tlv[99], \tlvp_rsm_usr_ob_tlv.ordern [7]);
tran (tlvp_rsm_usr_ob_tlv[100], \tlvp_rsm_usr_ob_tlv.ordern [8]);
tran (tlvp_rsm_usr_ob_tlv[101], \tlvp_rsm_usr_ob_tlv.ordern [9]);
tran (tlvp_rsm_usr_ob_tlv[102], \tlvp_rsm_usr_ob_tlv.ordern [10]);
tran (tlvp_rsm_usr_ob_tlv[103], \tlvp_rsm_usr_ob_tlv.ordern [11]);
tran (tlvp_rsm_usr_ob_tlv[104], \tlvp_rsm_usr_ob_tlv.ordern [12]);
tran (tlvp_rsm_usr_ob_tlv[105], \tlvp_rsm_usr_ob_tlv.insert );
tran (tlvp_rsm_usr_ob_rdata_dw0[0], \tlvp_rsm_usr_ob_rdata_dw0.tlv_type [0]);
tran (tlvp_rsm_usr_ob_rdata_dw0[1], \tlvp_rsm_usr_ob_rdata_dw0.tlv_type [1]);
tran (tlvp_rsm_usr_ob_rdata_dw0[2], \tlvp_rsm_usr_ob_rdata_dw0.tlv_type [2]);
tran (tlvp_rsm_usr_ob_rdata_dw0[3], \tlvp_rsm_usr_ob_rdata_dw0.tlv_type [3]);
tran (tlvp_rsm_usr_ob_rdata_dw0[4], \tlvp_rsm_usr_ob_rdata_dw0.tlv_type [4]);
tran (tlvp_rsm_usr_ob_rdata_dw0[5], \tlvp_rsm_usr_ob_rdata_dw0.tlv_type [5]);
tran (tlvp_rsm_usr_ob_rdata_dw0[6], \tlvp_rsm_usr_ob_rdata_dw0.tlv_type [6]);
tran (tlvp_rsm_usr_ob_rdata_dw0[7], \tlvp_rsm_usr_ob_rdata_dw0.tlv_type [7]);
tran (tlvp_rsm_usr_ob_rdata_dw0[8], \tlvp_rsm_usr_ob_rdata_dw0.tlv_len [0]);
tran (tlvp_rsm_usr_ob_rdata_dw0[9], \tlvp_rsm_usr_ob_rdata_dw0.tlv_len [1]);
tran (tlvp_rsm_usr_ob_rdata_dw0[10], \tlvp_rsm_usr_ob_rdata_dw0.tlv_len [2]);
tran (tlvp_rsm_usr_ob_rdata_dw0[11], \tlvp_rsm_usr_ob_rdata_dw0.tlv_len [3]);
tran (tlvp_rsm_usr_ob_rdata_dw0[12], \tlvp_rsm_usr_ob_rdata_dw0.tlv_len [4]);
tran (tlvp_rsm_usr_ob_rdata_dw0[13], \tlvp_rsm_usr_ob_rdata_dw0.tlv_len [5]);
tran (tlvp_rsm_usr_ob_rdata_dw0[14], \tlvp_rsm_usr_ob_rdata_dw0.tlv_len [6]);
tran (tlvp_rsm_usr_ob_rdata_dw0[15], \tlvp_rsm_usr_ob_rdata_dw0.tlv_len [7]);
tran (tlvp_rsm_usr_ob_rdata_dw0[16], \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num [0]);
tran (tlvp_rsm_usr_ob_rdata_dw0[17], \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num [1]);
tran (tlvp_rsm_usr_ob_rdata_dw0[18], \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num [2]);
tran (tlvp_rsm_usr_ob_rdata_dw0[19], \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num [3]);
tran (tlvp_rsm_usr_ob_rdata_dw0[20], \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num [4]);
tran (tlvp_rsm_usr_ob_rdata_dw0[21], \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num [5]);
tran (tlvp_rsm_usr_ob_rdata_dw0[22], \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num [6]);
tran (tlvp_rsm_usr_ob_rdata_dw0[23], \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num [7]);
tran (tlvp_rsm_usr_ob_rdata_dw0[24], \tlvp_rsm_usr_ob_rdata_dw0.tlv_eng_id [0]);
tran (tlvp_rsm_usr_ob_rdata_dw0[25], \tlvp_rsm_usr_ob_rdata_dw0.tlv_eng_id [1]);
tran (tlvp_rsm_usr_ob_rdata_dw0[26], \tlvp_rsm_usr_ob_rdata_dw0.tlv_eng_id [2]);
tran (tlvp_rsm_usr_ob_rdata_dw0[27], \tlvp_rsm_usr_ob_rdata_dw0.tlv_eng_id [3]);
tran (tlvp_rsm_usr_ob_rdata_dw0[28], \tlvp_rsm_usr_ob_rdata_dw0.resv1 [0]);
tran (tlvp_rsm_usr_ob_rdata_dw0[29], \tlvp_rsm_usr_ob_rdata_dw0.resv1 [1]);
tran (tlvp_rsm_usr_ob_rdata_dw0[30], \tlvp_rsm_usr_ob_rdata_dw0.resv1 [2]);
tran (tlvp_rsm_usr_ob_rdata_dw0[31], \tlvp_rsm_usr_ob_rdata_dw0.resv1 [3]);
tran (tlvp_rsm_usr_ob_rdata_dw0[32], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [0]);
tran (tlvp_rsm_usr_ob_rdata_dw0[33], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [1]);
tran (tlvp_rsm_usr_ob_rdata_dw0[34], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [2]);
tran (tlvp_rsm_usr_ob_rdata_dw0[35], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [3]);
tran (tlvp_rsm_usr_ob_rdata_dw0[36], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [4]);
tran (tlvp_rsm_usr_ob_rdata_dw0[37], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [5]);
tran (tlvp_rsm_usr_ob_rdata_dw0[38], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [6]);
tran (tlvp_rsm_usr_ob_rdata_dw0[39], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [7]);
tran (tlvp_rsm_usr_ob_rdata_dw0[40], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [8]);
tran (tlvp_rsm_usr_ob_rdata_dw0[41], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [9]);
tran (tlvp_rsm_usr_ob_rdata_dw0[42], \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num [10]);
tran (tlvp_rsm_usr_ob_rdata_dw0[43], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [0]);
tran (tlvp_rsm_usr_ob_rdata_dw0[44], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [1]);
tran (tlvp_rsm_usr_ob_rdata_dw0[45], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [2]);
tran (tlvp_rsm_usr_ob_rdata_dw0[46], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [3]);
tran (tlvp_rsm_usr_ob_rdata_dw0[47], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [4]);
tran (tlvp_rsm_usr_ob_rdata_dw0[48], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [5]);
tran (tlvp_rsm_usr_ob_rdata_dw0[49], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [6]);
tran (tlvp_rsm_usr_ob_rdata_dw0[50], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [7]);
tran (tlvp_rsm_usr_ob_rdata_dw0[51], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [8]);
tran (tlvp_rsm_usr_ob_rdata_dw0[52], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [9]);
tran (tlvp_rsm_usr_ob_rdata_dw0[53], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [10]);
tran (tlvp_rsm_usr_ob_rdata_dw0[54], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [11]);
tran (tlvp_rsm_usr_ob_rdata_dw0[55], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [12]);
tran (tlvp_rsm_usr_ob_rdata_dw0[56], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [13]);
tran (tlvp_rsm_usr_ob_rdata_dw0[57], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [14]);
tran (tlvp_rsm_usr_ob_rdata_dw0[58], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [15]);
tran (tlvp_rsm_usr_ob_rdata_dw0[59], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [16]);
tran (tlvp_rsm_usr_ob_rdata_dw0[60], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [17]);
tran (tlvp_rsm_usr_ob_rdata_dw0[61], \tlvp_rsm_usr_ob_rdata_dw0.resv0 [18]);
tran (tlvp_rsm_usr_ob_rdata_dw0[62], \tlvp_rsm_usr_ob_rdata_dw0.tlv_bip2 [0]);
tran (tlvp_rsm_usr_ob_rdata_dw0[63], \tlvp_rsm_usr_ob_rdata_dw0.tlv_bip2 [1]);
Q_BUF U0 ( .A(n1), .Z(next_state[2]));
Q_BUF U1 ( .A(n1), .Z(next_state[3]));
Q_BUF U2 ( .A(n1), .Z(next_state[4]));
Q_BUF U3 ( .A(n1), .Z(next_state[5]));
Q_BUF U4 ( .A(n1), .Z(next_state[6]));
Q_BUF U5 ( .A(n1), .Z(next_state[7]));
Q_BUF U6 ( .A(n1), .Z(next_state[8]));
Q_BUF U7 ( .A(n1), .Z(next_state[9]));
Q_BUF U8 ( .A(n1), .Z(next_state[10]));
Q_BUF U9 ( .A(n1), .Z(next_state[11]));
Q_BUF U10 ( .A(n1), .Z(next_state[12]));
Q_BUF U11 ( .A(n1), .Z(next_state[13]));
Q_BUF U12 ( .A(n1), .Z(next_state[14]));
Q_BUF U13 ( .A(n1), .Z(next_state[15]));
Q_BUF U14 ( .A(n1), .Z(next_state[16]));
Q_BUF U15 ( .A(n1), .Z(next_state[17]));
Q_BUF U16 ( .A(n1), .Z(next_state[18]));
Q_BUF U17 ( .A(n1), .Z(next_state[19]));
Q_BUF U18 ( .A(n1), .Z(next_state[20]));
Q_BUF U19 ( .A(n1), .Z(next_state[21]));
Q_BUF U20 ( .A(n1), .Z(next_state[22]));
Q_BUF U21 ( .A(n1), .Z(next_state[23]));
Q_BUF U22 ( .A(n1), .Z(next_state[24]));
Q_BUF U23 ( .A(n1), .Z(next_state[25]));
Q_BUF U24 ( .A(n1), .Z(next_state[26]));
Q_BUF U25 ( .A(n1), .Z(next_state[27]));
Q_BUF U26 ( .A(n1), .Z(next_state[28]));
Q_BUF U27 ( .A(n1), .Z(next_state[29]));
Q_BUF U28 ( .A(n1), .Z(next_state[30]));
Q_BUF U29 ( .A(n1), .Z(next_state[31]));
Q_XOR3 U30 ( .A0(tlvp_rsm_usr_ob_rdata[4]), .A1(tlvp_rsm_usr_ob_rdata[0]), .A2(tlvp_rsm_usr_ob_rdata[2]), .Z(n437));
Q_XOR3 U31 ( .A0(tlvp_rsm_usr_ob_rdata[10]), .A1(tlvp_rsm_usr_ob_rdata[6]), .A2(tlvp_rsm_usr_ob_rdata[8]), .Z(n436));
Q_XOR3 U32 ( .A0(tlvp_rsm_usr_ob_rdata[16]), .A1(tlvp_rsm_usr_ob_rdata[12]), .A2(tlvp_rsm_usr_ob_rdata[14]), .Z(n435));
Q_XOR3 U33 ( .A0(tlvp_rsm_usr_ob_rdata[22]), .A1(tlvp_rsm_usr_ob_rdata[18]), .A2(tlvp_rsm_usr_ob_rdata[20]), .Z(n434));
Q_XOR3 U34 ( .A0(tlvp_rsm_usr_ob_rdata[28]), .A1(tlvp_rsm_usr_ob_rdata[24]), .A2(tlvp_rsm_usr_ob_rdata[26]), .Z(n433));
Q_XOR3 U35 ( .A0(tlvp_rsm_usr_ob_rdata[34]), .A1(tlvp_rsm_usr_ob_rdata[30]), .A2(tlvp_rsm_usr_ob_rdata[32]), .Z(n432));
Q_XOR3 U36 ( .A0(tlvp_rsm_usr_ob_rdata[40]), .A1(tlvp_rsm_usr_ob_rdata[36]), .A2(tlvp_rsm_usr_ob_rdata[38]), .Z(n431));
Q_XOR3 U37 ( .A0(tlvp_rsm_usr_ob_rdata[46]), .A1(tlvp_rsm_usr_ob_rdata[42]), .A2(tlvp_rsm_usr_ob_rdata[44]), .Z(n430));
Q_XOR3 U38 ( .A0(tlvp_rsm_usr_ob_rdata[52]), .A1(tlvp_rsm_usr_ob_rdata[48]), .A2(tlvp_rsm_usr_ob_rdata[50]), .Z(n429));
Q_XOR3 U39 ( .A0(tlvp_rsm_usr_ob_rdata[58]), .A1(tlvp_rsm_usr_ob_rdata[54]), .A2(tlvp_rsm_usr_ob_rdata[56]), .Z(n428));
Q_XOR3 U40 ( .A0(n436), .A1(tlvp_rsm_usr_ob_rdata[60]), .A2(n437), .Z(n427));
Q_XOR3 U41 ( .A0(n433), .A1(n435), .A2(n434), .Z(n426));
Q_XOR3 U42 ( .A0(n430), .A1(n432), .A2(n431), .Z(n425));
Q_XOR3 U43 ( .A0(n427), .A1(n429), .A2(n428), .Z(n424));
Q_XOR3 U44 ( .A0(n424), .A1(n426), .A2(n425), .Z(tlvp_rsm_bip2[0]));
Q_XOR3 U45 ( .A0(tlvp_rsm_usr_ob_rdata[5]), .A1(tlvp_rsm_usr_ob_rdata[1]), .A2(tlvp_rsm_usr_ob_rdata[3]), .Z(n423));
Q_XOR3 U46 ( .A0(tlvp_rsm_usr_ob_rdata[11]), .A1(tlvp_rsm_usr_ob_rdata[7]), .A2(tlvp_rsm_usr_ob_rdata[9]), .Z(n422));
Q_XOR3 U47 ( .A0(tlvp_rsm_usr_ob_rdata[17]), .A1(tlvp_rsm_usr_ob_rdata[13]), .A2(tlvp_rsm_usr_ob_rdata[15]), .Z(n421));
Q_XOR3 U48 ( .A0(tlvp_rsm_usr_ob_rdata[23]), .A1(tlvp_rsm_usr_ob_rdata[19]), .A2(tlvp_rsm_usr_ob_rdata[21]), .Z(n420));
Q_XOR3 U49 ( .A0(tlvp_rsm_usr_ob_rdata[29]), .A1(tlvp_rsm_usr_ob_rdata[25]), .A2(tlvp_rsm_usr_ob_rdata[27]), .Z(n419));
Q_XOR3 U50 ( .A0(tlvp_rsm_usr_ob_rdata[35]), .A1(tlvp_rsm_usr_ob_rdata[31]), .A2(tlvp_rsm_usr_ob_rdata[33]), .Z(n418));
Q_XOR3 U51 ( .A0(tlvp_rsm_usr_ob_rdata[41]), .A1(tlvp_rsm_usr_ob_rdata[37]), .A2(tlvp_rsm_usr_ob_rdata[39]), .Z(n417));
Q_XOR3 U52 ( .A0(tlvp_rsm_usr_ob_rdata[47]), .A1(tlvp_rsm_usr_ob_rdata[43]), .A2(tlvp_rsm_usr_ob_rdata[45]), .Z(n416));
Q_XOR3 U53 ( .A0(tlvp_rsm_usr_ob_rdata[53]), .A1(tlvp_rsm_usr_ob_rdata[49]), .A2(tlvp_rsm_usr_ob_rdata[51]), .Z(n415));
Q_XOR3 U54 ( .A0(tlvp_rsm_usr_ob_rdata[59]), .A1(tlvp_rsm_usr_ob_rdata[55]), .A2(tlvp_rsm_usr_ob_rdata[57]), .Z(n414));
Q_XOR3 U55 ( .A0(n422), .A1(tlvp_rsm_usr_ob_rdata[61]), .A2(n423), .Z(n413));
Q_XOR3 U56 ( .A0(n419), .A1(n421), .A2(n420), .Z(n412));
Q_XOR3 U57 ( .A0(n416), .A1(n418), .A2(n417), .Z(n411));
Q_XOR3 U58 ( .A0(n413), .A1(n415), .A2(n414), .Z(n410));
Q_XOR3 U59 ( .A0(n410), .A1(n412), .A2(n411), .Z(tlvp_rsm_bip2[1]));
Q_INV U60 ( .A(next_state[1]), .Z(n13));
Q_INV U61 ( .A(next_state[0]), .Z(n5));
Q_NR02 U62 ( .A0(next_state[0]), .A1(tlvp_rsm_usr_ob_tlv[83]), .Z(n6));
Q_OR02 U63 ( .A0(n13), .A1(n6), .Z(n7));
Q_NR02 U64 ( .A0(next_state[1]), .A1(next_state[0]), .Z(n8));
Q_NR02 U65 ( .A0(tlvp_rsm_usr_ob_tlv[81]), .A1(tlvp_rsm_usr_ob_tlv[82]), .Z(n9));
Q_OA21 U66 ( .A0(n13), .A1(n9), .B0(n5), .Z(n11));
Q_NR02 U67 ( .A0(tlvp_rsm_pt_tlv[81]), .A1(tlvp_rsm_pt_tlv[82]), .Z(n10));
Q_AO21 U68 ( .A0(n13), .A1(n10), .B0(n11), .Z(n12));
Q_AN02 U69 ( .A0(n13), .A1(next_state[0]), .Z(n3));
Q_AN02 U70 ( .A0(next_state[1]), .A1(n5), .Z(n4));
Q_AN02 U71 ( .A0(n3), .A1(n14), .Z(n16));
Q_AO21 U72 ( .A0(n4), .A1(n15), .B0(n16), .Z(n2));
Q_MX02 U73 ( .S(n8), .A0(n266), .A1(tlvp_rsm_last_typen[0]), .Z(n17));
Q_FDP2 \tlvp_rsm_last_typen_REG[0] ( .CK(clk), .S(rst_n), .D(n17), .Q(tlvp_rsm_last_typen[0]), .QN( ));
Q_MX02 U75 ( .S(n8), .A0(n264), .A1(tlvp_rsm_last_typen[1]), .Z(n18));
Q_FDP2 \tlvp_rsm_last_typen_REG[1] ( .CK(clk), .S(rst_n), .D(n18), .Q(tlvp_rsm_last_typen[1]), .QN( ));
Q_MX02 U77 ( .S(n8), .A0(n262), .A1(tlvp_rsm_last_typen[2]), .Z(n19));
Q_FDP2 \tlvp_rsm_last_typen_REG[2] ( .CK(clk), .S(rst_n), .D(n19), .Q(tlvp_rsm_last_typen[2]), .QN( ));
Q_MX02 U79 ( .S(n8), .A0(n260), .A1(tlvp_rsm_last_typen[3]), .Z(n20));
Q_FDP2 \tlvp_rsm_last_typen_REG[3] ( .CK(clk), .S(rst_n), .D(n20), .Q(tlvp_rsm_last_typen[3]), .QN( ));
Q_MX02 U81 ( .S(n8), .A0(n258), .A1(tlvp_rsm_last_typen[4]), .Z(n21));
Q_FDP2 \tlvp_rsm_last_typen_REG[4] ( .CK(clk), .S(rst_n), .D(n21), .Q(tlvp_rsm_last_typen[4]), .QN( ));
Q_MX02 U83 ( .S(n8), .A0(n256), .A1(tlvp_rsm_last_typen[5]), .Z(n22));
Q_FDP2 \tlvp_rsm_last_typen_REG[5] ( .CK(clk), .S(rst_n), .D(n22), .Q(tlvp_rsm_last_typen[5]), .QN( ));
Q_MX02 U85 ( .S(n8), .A0(n254), .A1(tlvp_rsm_last_typen[6]), .Z(n23));
Q_FDP2 \tlvp_rsm_last_typen_REG[6] ( .CK(clk), .S(rst_n), .D(n23), .Q(tlvp_rsm_last_typen[6]), .QN( ));
Q_MX02 U87 ( .S(n8), .A0(n252), .A1(tlvp_rsm_last_typen[7]), .Z(n24));
Q_FDP2 \tlvp_rsm_last_typen_REG[7] ( .CK(clk), .S(rst_n), .D(n24), .Q(tlvp_rsm_last_typen[7]), .QN( ));
Q_MX02 U89 ( .S(n12), .A0(n251), .A1(tlvp_rsm_nxt_ordern[0]), .Z(n25));
Q_FDP2 \tlvp_rsm_nxt_ordern_REG[0] ( .CK(clk), .S(rst_n), .D(n25), .Q(tlvp_rsm_nxt_ordern[0]), .QN(n462));
Q_FDP1 \tlvp_rsm_ob_datain_REG[0] ( .CK(clk), .R(rst_n), .D(n237), .Q(tlvp_rsm_ob_datain[0]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[1] ( .CK(clk), .R(rst_n), .D(n235), .Q(tlvp_rsm_ob_datain[1]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[2] ( .CK(clk), .R(rst_n), .D(n233), .Q(tlvp_rsm_ob_datain[2]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[3] ( .CK(clk), .R(rst_n), .D(n231), .Q(tlvp_rsm_ob_datain[3]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[4] ( .CK(clk), .R(rst_n), .D(n229), .Q(tlvp_rsm_ob_datain[4]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[5] ( .CK(clk), .R(rst_n), .D(n227), .Q(tlvp_rsm_ob_datain[5]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[6] ( .CK(clk), .R(rst_n), .D(n225), .Q(tlvp_rsm_ob_datain[6]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[7] ( .CK(clk), .R(rst_n), .D(n223), .Q(tlvp_rsm_ob_datain[7]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[8] ( .CK(clk), .R(rst_n), .D(n221), .Q(tlvp_rsm_ob_datain[8]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[9] ( .CK(clk), .R(rst_n), .D(n219), .Q(tlvp_rsm_ob_datain[9]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[10] ( .CK(clk), .R(rst_n), .D(n217), .Q(tlvp_rsm_ob_datain[10]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[11] ( .CK(clk), .R(rst_n), .D(n215), .Q(tlvp_rsm_ob_datain[11]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[12] ( .CK(clk), .R(rst_n), .D(n213), .Q(tlvp_rsm_ob_datain[12]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[13] ( .CK(clk), .R(rst_n), .D(n211), .Q(tlvp_rsm_ob_datain[13]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[14] ( .CK(clk), .R(rst_n), .D(n209), .Q(tlvp_rsm_ob_datain[14]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[15] ( .CK(clk), .R(rst_n), .D(n207), .Q(tlvp_rsm_ob_datain[15]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[16] ( .CK(clk), .R(rst_n), .D(n205), .Q(tlvp_rsm_ob_datain[16]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[17] ( .CK(clk), .R(rst_n), .D(n203), .Q(tlvp_rsm_ob_datain[17]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[18] ( .CK(clk), .R(rst_n), .D(n201), .Q(tlvp_rsm_ob_datain[18]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[19] ( .CK(clk), .R(rst_n), .D(n199), .Q(tlvp_rsm_ob_datain[19]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[20] ( .CK(clk), .R(rst_n), .D(n197), .Q(tlvp_rsm_ob_datain[20]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[21] ( .CK(clk), .R(rst_n), .D(n195), .Q(tlvp_rsm_ob_datain[21]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[22] ( .CK(clk), .R(rst_n), .D(n193), .Q(tlvp_rsm_ob_datain[22]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[23] ( .CK(clk), .R(rst_n), .D(n191), .Q(tlvp_rsm_ob_datain[23]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[24] ( .CK(clk), .R(rst_n), .D(n189), .Q(tlvp_rsm_ob_datain[24]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[25] ( .CK(clk), .R(rst_n), .D(n187), .Q(tlvp_rsm_ob_datain[25]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[26] ( .CK(clk), .R(rst_n), .D(n185), .Q(tlvp_rsm_ob_datain[26]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[27] ( .CK(clk), .R(rst_n), .D(n183), .Q(tlvp_rsm_ob_datain[27]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[28] ( .CK(clk), .R(rst_n), .D(n181), .Q(tlvp_rsm_ob_datain[28]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[29] ( .CK(clk), .R(rst_n), .D(n179), .Q(tlvp_rsm_ob_datain[29]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[30] ( .CK(clk), .R(rst_n), .D(n177), .Q(tlvp_rsm_ob_datain[30]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[31] ( .CK(clk), .R(rst_n), .D(n175), .Q(tlvp_rsm_ob_datain[31]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[32] ( .CK(clk), .R(rst_n), .D(n173), .Q(tlvp_rsm_ob_datain[32]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[33] ( .CK(clk), .R(rst_n), .D(n171), .Q(tlvp_rsm_ob_datain[33]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[34] ( .CK(clk), .R(rst_n), .D(n169), .Q(tlvp_rsm_ob_datain[34]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[35] ( .CK(clk), .R(rst_n), .D(n167), .Q(tlvp_rsm_ob_datain[35]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[36] ( .CK(clk), .R(rst_n), .D(n165), .Q(tlvp_rsm_ob_datain[36]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[37] ( .CK(clk), .R(rst_n), .D(n163), .Q(tlvp_rsm_ob_datain[37]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[38] ( .CK(clk), .R(rst_n), .D(n161), .Q(tlvp_rsm_ob_datain[38]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[39] ( .CK(clk), .R(rst_n), .D(n159), .Q(tlvp_rsm_ob_datain[39]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[40] ( .CK(clk), .R(rst_n), .D(n157), .Q(tlvp_rsm_ob_datain[40]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[41] ( .CK(clk), .R(rst_n), .D(n155), .Q(tlvp_rsm_ob_datain[41]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[42] ( .CK(clk), .R(rst_n), .D(n153), .Q(tlvp_rsm_ob_datain[42]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[43] ( .CK(clk), .R(rst_n), .D(n151), .Q(tlvp_rsm_ob_datain[43]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[44] ( .CK(clk), .R(rst_n), .D(n149), .Q(tlvp_rsm_ob_datain[44]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[45] ( .CK(clk), .R(rst_n), .D(n147), .Q(tlvp_rsm_ob_datain[45]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[46] ( .CK(clk), .R(rst_n), .D(n145), .Q(tlvp_rsm_ob_datain[46]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[47] ( .CK(clk), .R(rst_n), .D(n143), .Q(tlvp_rsm_ob_datain[47]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[48] ( .CK(clk), .R(rst_n), .D(n141), .Q(tlvp_rsm_ob_datain[48]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[49] ( .CK(clk), .R(rst_n), .D(n139), .Q(tlvp_rsm_ob_datain[49]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[50] ( .CK(clk), .R(rst_n), .D(n137), .Q(tlvp_rsm_ob_datain[50]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[51] ( .CK(clk), .R(rst_n), .D(n135), .Q(tlvp_rsm_ob_datain[51]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[52] ( .CK(clk), .R(rst_n), .D(n133), .Q(tlvp_rsm_ob_datain[52]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[53] ( .CK(clk), .R(rst_n), .D(n131), .Q(tlvp_rsm_ob_datain[53]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[54] ( .CK(clk), .R(rst_n), .D(n129), .Q(tlvp_rsm_ob_datain[54]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[55] ( .CK(clk), .R(rst_n), .D(n127), .Q(tlvp_rsm_ob_datain[55]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[56] ( .CK(clk), .R(rst_n), .D(n125), .Q(tlvp_rsm_ob_datain[56]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[57] ( .CK(clk), .R(rst_n), .D(n123), .Q(tlvp_rsm_ob_datain[57]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[58] ( .CK(clk), .R(rst_n), .D(n121), .Q(tlvp_rsm_ob_datain[58]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[59] ( .CK(clk), .R(rst_n), .D(n119), .Q(tlvp_rsm_ob_datain[59]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[60] ( .CK(clk), .R(rst_n), .D(n117), .Q(tlvp_rsm_ob_datain[60]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[61] ( .CK(clk), .R(rst_n), .D(n115), .Q(tlvp_rsm_ob_datain[61]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[62] ( .CK(clk), .R(rst_n), .D(n113), .Q(tlvp_rsm_ob_datain[62]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[63] ( .CK(clk), .R(rst_n), .D(n111), .Q(tlvp_rsm_ob_datain[63]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[64] ( .CK(clk), .R(rst_n), .D(n109), .Q(tlvp_rsm_ob_datain[64]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[65] ( .CK(clk), .R(rst_n), .D(n107), .Q(tlvp_rsm_ob_datain[65]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[66] ( .CK(clk), .R(rst_n), .D(n105), .Q(tlvp_rsm_ob_datain[66]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[67] ( .CK(clk), .R(rst_n), .D(n103), .Q(tlvp_rsm_ob_datain[67]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[68] ( .CK(clk), .R(rst_n), .D(n101), .Q(tlvp_rsm_ob_datain[68]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[69] ( .CK(clk), .R(rst_n), .D(n99), .Q(tlvp_rsm_ob_datain[69]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[70] ( .CK(clk), .R(rst_n), .D(n97), .Q(tlvp_rsm_ob_datain[70]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[71] ( .CK(clk), .R(rst_n), .D(n95), .Q(tlvp_rsm_ob_datain[71]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[72] ( .CK(clk), .R(rst_n), .D(n93), .Q(tlvp_rsm_ob_datain[72]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[73] ( .CK(clk), .R(rst_n), .D(n91), .Q(tlvp_rsm_ob_datain[73]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[74] ( .CK(clk), .R(rst_n), .D(n89), .Q(tlvp_rsm_ob_datain[74]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[75] ( .CK(clk), .R(rst_n), .D(n87), .Q(tlvp_rsm_ob_datain[75]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[76] ( .CK(clk), .R(rst_n), .D(n85), .Q(tlvp_rsm_ob_datain[76]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[77] ( .CK(clk), .R(rst_n), .D(n83), .Q(tlvp_rsm_ob_datain[77]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[78] ( .CK(clk), .R(rst_n), .D(n81), .Q(tlvp_rsm_ob_datain[78]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[79] ( .CK(clk), .R(rst_n), .D(n79), .Q(tlvp_rsm_ob_datain[79]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[80] ( .CK(clk), .R(rst_n), .D(n77), .Q(tlvp_rsm_ob_datain[80]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[81] ( .CK(clk), .R(rst_n), .D(n75), .Q(tlvp_rsm_ob_datain[81]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[82] ( .CK(clk), .R(rst_n), .D(n73), .Q(tlvp_rsm_ob_datain[82]), .QN(n316));
Q_FDP1 \tlvp_rsm_ob_datain_REG[83] ( .CK(clk), .R(rst_n), .D(n71), .Q(tlvp_rsm_ob_datain[83]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[84] ( .CK(clk), .R(rst_n), .D(n69), .Q(tlvp_rsm_ob_datain[84]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[85] ( .CK(clk), .R(rst_n), .D(n67), .Q(tlvp_rsm_ob_datain[85]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[86] ( .CK(clk), .R(rst_n), .D(n65), .Q(tlvp_rsm_ob_datain[86]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[87] ( .CK(clk), .R(rst_n), .D(n63), .Q(tlvp_rsm_ob_datain[87]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[88] ( .CK(clk), .R(rst_n), .D(n61), .Q(tlvp_rsm_ob_datain[88]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[89] ( .CK(clk), .R(rst_n), .D(n59), .Q(tlvp_rsm_ob_datain[89]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[90] ( .CK(clk), .R(rst_n), .D(n57), .Q(tlvp_rsm_ob_datain[90]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[91] ( .CK(clk), .R(rst_n), .D(n55), .Q(tlvp_rsm_ob_datain[91]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[92] ( .CK(clk), .R(rst_n), .D(n53), .Q(tlvp_rsm_ob_datain[92]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[93] ( .CK(clk), .R(rst_n), .D(n51), .Q(tlvp_rsm_ob_datain[93]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[94] ( .CK(clk), .R(rst_n), .D(n49), .Q(tlvp_rsm_ob_datain[94]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[95] ( .CK(clk), .R(rst_n), .D(n47), .Q(tlvp_rsm_ob_datain[95]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[96] ( .CK(clk), .R(rst_n), .D(n45), .Q(tlvp_rsm_ob_datain[96]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[97] ( .CK(clk), .R(rst_n), .D(n43), .Q(tlvp_rsm_ob_datain[97]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[98] ( .CK(clk), .R(rst_n), .D(n41), .Q(tlvp_rsm_ob_datain[98]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[99] ( .CK(clk), .R(rst_n), .D(n39), .Q(tlvp_rsm_ob_datain[99]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[100] ( .CK(clk), .R(rst_n), .D(n37), .Q(tlvp_rsm_ob_datain[100]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[101] ( .CK(clk), .R(rst_n), .D(n35), .Q(tlvp_rsm_ob_datain[101]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[102] ( .CK(clk), .R(rst_n), .D(n33), .Q(tlvp_rsm_ob_datain[102]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[103] ( .CK(clk), .R(rst_n), .D(n31), .Q(tlvp_rsm_ob_datain[103]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[104] ( .CK(clk), .R(rst_n), .D(n29), .Q(tlvp_rsm_ob_datain[104]), .QN( ));
Q_FDP1 \tlvp_rsm_ob_datain_REG[105] ( .CK(clk), .R(rst_n), .D(n27), .Q(tlvp_rsm_ob_datain[105]), .QN( ));
Q_FDP1 tlvp_rsm_ob_wen_REG  ( .CK(clk), .R(rst_n), .D(n26), .Q(tlvp_rsm_ob_wen), .QN( ));
Q_MX02 U198 ( .S(n3), .A0(tlvp_rsm_usr_ob_wen), .A1(tlvp_rsm_pt_valid), .Z(n26));
Q_AN02 U199 ( .A0(n4), .A1(tlvp_rsm_usr_ob_valid), .Z(tlvp_rsm_usr_ob_wen));
Q_MX02 U200 ( .S(n3), .A0(n28), .A1(tlvp_rsm_pt_tlv[105]), .Z(n27));
Q_AN02 U201 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[105]), .Z(n28));
Q_MX02 U202 ( .S(n3), .A0(n30), .A1(tlvp_rsm_pt_tlv[104]), .Z(n29));
Q_AN02 U203 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[104]), .Z(n30));
Q_MX02 U204 ( .S(n3), .A0(n32), .A1(tlvp_rsm_pt_tlv[103]), .Z(n31));
Q_AN02 U205 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[103]), .Z(n32));
Q_MX02 U206 ( .S(n3), .A0(n34), .A1(tlvp_rsm_pt_tlv[102]), .Z(n33));
Q_AN02 U207 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[102]), .Z(n34));
Q_MX02 U208 ( .S(n3), .A0(n36), .A1(tlvp_rsm_pt_tlv[101]), .Z(n35));
Q_AN02 U209 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[101]), .Z(n36));
Q_MX02 U210 ( .S(n3), .A0(n38), .A1(tlvp_rsm_pt_tlv[100]), .Z(n37));
Q_AN02 U211 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[100]), .Z(n38));
Q_MX02 U212 ( .S(n3), .A0(n40), .A1(tlvp_rsm_pt_tlv[99]), .Z(n39));
Q_AN02 U213 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[99]), .Z(n40));
Q_MX02 U214 ( .S(n3), .A0(n42), .A1(tlvp_rsm_pt_tlv[98]), .Z(n41));
Q_AN02 U215 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[98]), .Z(n42));
Q_MX02 U216 ( .S(n3), .A0(n44), .A1(tlvp_rsm_pt_tlv[97]), .Z(n43));
Q_AN02 U217 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[97]), .Z(n44));
Q_MX02 U218 ( .S(n3), .A0(n46), .A1(tlvp_rsm_pt_tlv[96]), .Z(n45));
Q_AN02 U219 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[96]), .Z(n46));
Q_MX02 U220 ( .S(n3), .A0(n48), .A1(tlvp_rsm_pt_tlv[95]), .Z(n47));
Q_AN02 U221 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[95]), .Z(n48));
Q_MX02 U222 ( .S(n3), .A0(n50), .A1(tlvp_rsm_pt_tlv[94]), .Z(n49));
Q_AN02 U223 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[94]), .Z(n50));
Q_MX02 U224 ( .S(n3), .A0(n52), .A1(tlvp_rsm_pt_tlv[93]), .Z(n51));
Q_AN02 U225 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[93]), .Z(n52));
Q_MX02 U226 ( .S(n3), .A0(n54), .A1(tlvp_rsm_pt_tlv[92]), .Z(n53));
Q_AN02 U227 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[92]), .Z(n54));
Q_MX02 U228 ( .S(n3), .A0(n56), .A1(tlvp_rsm_pt_tlv[91]), .Z(n55));
Q_AN02 U229 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[91]), .Z(n56));
Q_MX02 U230 ( .S(n3), .A0(n58), .A1(tlvp_rsm_pt_tlv[90]), .Z(n57));
Q_AN02 U231 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[90]), .Z(n58));
Q_MX02 U232 ( .S(n3), .A0(n60), .A1(tlvp_rsm_pt_tlv[89]), .Z(n59));
Q_AN02 U233 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[89]), .Z(n60));
Q_MX02 U234 ( .S(n3), .A0(n62), .A1(tlvp_rsm_pt_tlv[88]), .Z(n61));
Q_AN02 U235 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[88]), .Z(n62));
Q_MX02 U236 ( .S(n3), .A0(n64), .A1(tlvp_rsm_pt_tlv[87]), .Z(n63));
Q_AN02 U237 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[87]), .Z(n64));
Q_MX02 U238 ( .S(n3), .A0(n66), .A1(tlvp_rsm_pt_tlv[86]), .Z(n65));
Q_AN02 U239 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[86]), .Z(n66));
Q_MX02 U240 ( .S(n3), .A0(n68), .A1(tlvp_rsm_pt_tlv[85]), .Z(n67));
Q_AN02 U241 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[85]), .Z(n68));
Q_MX02 U242 ( .S(n3), .A0(n70), .A1(tlvp_rsm_pt_tlv[84]), .Z(n69));
Q_AN02 U243 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[84]), .Z(n70));
Q_MX02 U244 ( .S(n3), .A0(n72), .A1(tlvp_rsm_pt_tlv[83]), .Z(n71));
Q_AN02 U245 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[83]), .Z(n72));
Q_MX02 U246 ( .S(n3), .A0(n74), .A1(tlvp_rsm_pt_tlv[82]), .Z(n73));
Q_AN02 U247 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[82]), .Z(n74));
Q_MX02 U248 ( .S(n3), .A0(n76), .A1(tlvp_rsm_pt_tlv[81]), .Z(n75));
Q_AN02 U249 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[81]), .Z(n76));
Q_MX02 U250 ( .S(n3), .A0(n78), .A1(tlvp_rsm_pt_tlv[80]), .Z(n77));
Q_AN02 U251 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[80]), .Z(n78));
Q_MX02 U252 ( .S(n3), .A0(n80), .A1(tlvp_rsm_pt_tlv[79]), .Z(n79));
Q_AN02 U253 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[79]), .Z(n80));
Q_MX02 U254 ( .S(n3), .A0(n82), .A1(tlvp_rsm_pt_tlv[78]), .Z(n81));
Q_AN02 U255 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[78]), .Z(n82));
Q_MX02 U256 ( .S(n3), .A0(n84), .A1(tlvp_rsm_pt_tlv[77]), .Z(n83));
Q_AN02 U257 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[77]), .Z(n84));
Q_MX02 U258 ( .S(n3), .A0(n86), .A1(tlvp_rsm_pt_tlv[76]), .Z(n85));
Q_AN02 U259 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[76]), .Z(n86));
Q_MX02 U260 ( .S(n3), .A0(n88), .A1(tlvp_rsm_pt_tlv[75]), .Z(n87));
Q_AN02 U261 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[75]), .Z(n88));
Q_MX02 U262 ( .S(n3), .A0(n90), .A1(tlvp_rsm_pt_tlv[74]), .Z(n89));
Q_AN02 U263 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[74]), .Z(n90));
Q_MX02 U264 ( .S(n3), .A0(n92), .A1(tlvp_rsm_pt_tlv[73]), .Z(n91));
Q_AN02 U265 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[73]), .Z(n92));
Q_MX02 U266 ( .S(n3), .A0(n94), .A1(tlvp_rsm_pt_tlv[72]), .Z(n93));
Q_AN02 U267 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[72]), .Z(n94));
Q_MX02 U268 ( .S(n3), .A0(n96), .A1(tlvp_rsm_pt_tlv[71]), .Z(n95));
Q_AN02 U269 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[71]), .Z(n96));
Q_MX02 U270 ( .S(n3), .A0(n98), .A1(tlvp_rsm_pt_tlv[70]), .Z(n97));
Q_AN02 U271 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[70]), .Z(n98));
Q_MX02 U272 ( .S(n3), .A0(n100), .A1(tlvp_rsm_pt_tlv[69]), .Z(n99));
Q_AN02 U273 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[69]), .Z(n100));
Q_MX02 U274 ( .S(n3), .A0(n102), .A1(tlvp_rsm_pt_tlv[68]), .Z(n101));
Q_AN02 U275 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[68]), .Z(n102));
Q_MX02 U276 ( .S(n3), .A0(n104), .A1(tlvp_rsm_pt_tlv[67]), .Z(n103));
Q_AN02 U277 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[67]), .Z(n104));
Q_MX02 U278 ( .S(n3), .A0(n106), .A1(tlvp_rsm_pt_tlv[66]), .Z(n105));
Q_AN02 U279 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[66]), .Z(n106));
Q_MX02 U280 ( .S(n3), .A0(n108), .A1(tlvp_rsm_pt_tlv[65]), .Z(n107));
Q_AN02 U281 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[65]), .Z(n108));
Q_MX02 U282 ( .S(n3), .A0(n110), .A1(tlvp_rsm_pt_tlv[64]), .Z(n109));
Q_AN02 U283 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[64]), .Z(n110));
Q_MX02 U284 ( .S(n3), .A0(n112), .A1(tlvp_rsm_pt_tlv[63]), .Z(n111));
Q_AN02 U285 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[63]), .Z(n112));
Q_MX02 U286 ( .S(n3), .A0(n114), .A1(tlvp_rsm_pt_tlv[62]), .Z(n113));
Q_AN02 U287 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[62]), .Z(n114));
Q_MX02 U288 ( .S(n3), .A0(n116), .A1(tlvp_rsm_pt_tlv[61]), .Z(n115));
Q_AN02 U289 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[61]), .Z(n116));
Q_MX02 U290 ( .S(n3), .A0(n118), .A1(tlvp_rsm_pt_tlv[60]), .Z(n117));
Q_AN02 U291 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[60]), .Z(n118));
Q_MX02 U292 ( .S(n3), .A0(n120), .A1(tlvp_rsm_pt_tlv[59]), .Z(n119));
Q_AN02 U293 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[59]), .Z(n120));
Q_MX02 U294 ( .S(n3), .A0(n122), .A1(tlvp_rsm_pt_tlv[58]), .Z(n121));
Q_AN02 U295 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[58]), .Z(n122));
Q_MX02 U296 ( .S(n3), .A0(n124), .A1(tlvp_rsm_pt_tlv[57]), .Z(n123));
Q_AN02 U297 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[57]), .Z(n124));
Q_MX02 U298 ( .S(n3), .A0(n126), .A1(tlvp_rsm_pt_tlv[56]), .Z(n125));
Q_AN02 U299 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[56]), .Z(n126));
Q_MX02 U300 ( .S(n3), .A0(n128), .A1(tlvp_rsm_pt_tlv[55]), .Z(n127));
Q_AN02 U301 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[55]), .Z(n128));
Q_MX02 U302 ( .S(n3), .A0(n130), .A1(tlvp_rsm_pt_tlv[54]), .Z(n129));
Q_AN02 U303 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[54]), .Z(n130));
Q_MX02 U304 ( .S(n3), .A0(n132), .A1(tlvp_rsm_pt_tlv[53]), .Z(n131));
Q_AN02 U305 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[53]), .Z(n132));
Q_MX02 U306 ( .S(n3), .A0(n134), .A1(tlvp_rsm_pt_tlv[52]), .Z(n133));
Q_AN02 U307 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[52]), .Z(n134));
Q_MX02 U308 ( .S(n3), .A0(n136), .A1(tlvp_rsm_pt_tlv[51]), .Z(n135));
Q_AN02 U309 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[51]), .Z(n136));
Q_MX02 U310 ( .S(n3), .A0(n138), .A1(tlvp_rsm_pt_tlv[50]), .Z(n137));
Q_AN02 U311 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[50]), .Z(n138));
Q_MX02 U312 ( .S(n3), .A0(n140), .A1(tlvp_rsm_pt_tlv[49]), .Z(n139));
Q_AN02 U313 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[49]), .Z(n140));
Q_MX02 U314 ( .S(n3), .A0(n142), .A1(tlvp_rsm_pt_tlv[48]), .Z(n141));
Q_AN02 U315 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[48]), .Z(n142));
Q_MX02 U316 ( .S(n3), .A0(n144), .A1(tlvp_rsm_pt_tlv[47]), .Z(n143));
Q_AN02 U317 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[47]), .Z(n144));
Q_MX02 U318 ( .S(n3), .A0(n146), .A1(tlvp_rsm_pt_tlv[46]), .Z(n145));
Q_AN02 U319 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[46]), .Z(n146));
Q_MX02 U320 ( .S(n3), .A0(n148), .A1(tlvp_rsm_pt_tlv[45]), .Z(n147));
Q_AN02 U321 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[45]), .Z(n148));
Q_MX02 U322 ( .S(n3), .A0(n150), .A1(tlvp_rsm_pt_tlv[44]), .Z(n149));
Q_AN02 U323 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[44]), .Z(n150));
Q_MX02 U324 ( .S(n3), .A0(n152), .A1(tlvp_rsm_pt_tlv[43]), .Z(n151));
Q_AN02 U325 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[43]), .Z(n152));
Q_MX02 U326 ( .S(n3), .A0(n154), .A1(tlvp_rsm_pt_tlv[42]), .Z(n153));
Q_AN02 U327 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[42]), .Z(n154));
Q_MX02 U328 ( .S(n3), .A0(n156), .A1(tlvp_rsm_pt_tlv[41]), .Z(n155));
Q_AN02 U329 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[41]), .Z(n156));
Q_MX02 U330 ( .S(n3), .A0(n158), .A1(tlvp_rsm_pt_tlv[40]), .Z(n157));
Q_AN02 U331 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[40]), .Z(n158));
Q_MX02 U332 ( .S(n3), .A0(n160), .A1(tlvp_rsm_pt_tlv[39]), .Z(n159));
Q_AN02 U333 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[39]), .Z(n160));
Q_MX02 U334 ( .S(n3), .A0(n162), .A1(tlvp_rsm_pt_tlv[38]), .Z(n161));
Q_AN02 U335 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[38]), .Z(n162));
Q_MX02 U336 ( .S(n3), .A0(n164), .A1(tlvp_rsm_pt_tlv[37]), .Z(n163));
Q_AN02 U337 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[37]), .Z(n164));
Q_MX02 U338 ( .S(n3), .A0(n166), .A1(tlvp_rsm_pt_tlv[36]), .Z(n165));
Q_AN02 U339 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[36]), .Z(n166));
Q_MX02 U340 ( .S(n3), .A0(n168), .A1(tlvp_rsm_pt_tlv[35]), .Z(n167));
Q_AN02 U341 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[35]), .Z(n168));
Q_MX02 U342 ( .S(n3), .A0(n170), .A1(tlvp_rsm_pt_tlv[34]), .Z(n169));
Q_AN02 U343 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[34]), .Z(n170));
Q_MX02 U344 ( .S(n3), .A0(n172), .A1(tlvp_rsm_pt_tlv[33]), .Z(n171));
Q_AN02 U345 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[33]), .Z(n172));
Q_MX02 U346 ( .S(n3), .A0(n174), .A1(tlvp_rsm_pt_tlv[32]), .Z(n173));
Q_AN02 U347 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[32]), .Z(n174));
Q_MX02 U348 ( .S(n3), .A0(n176), .A1(tlvp_rsm_pt_tlv[31]), .Z(n175));
Q_AN02 U349 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[31]), .Z(n176));
Q_MX02 U350 ( .S(n3), .A0(n178), .A1(tlvp_rsm_pt_tlv[30]), .Z(n177));
Q_AN02 U351 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[30]), .Z(n178));
Q_MX02 U352 ( .S(n3), .A0(n180), .A1(tlvp_rsm_pt_tlv[29]), .Z(n179));
Q_AN02 U353 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[29]), .Z(n180));
Q_MX02 U354 ( .S(n3), .A0(n182), .A1(tlvp_rsm_pt_tlv[28]), .Z(n181));
Q_AN02 U355 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[28]), .Z(n182));
Q_MX02 U356 ( .S(n3), .A0(n184), .A1(tlvp_rsm_pt_tlv[27]), .Z(n183));
Q_AN02 U357 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[27]), .Z(n184));
Q_MX02 U358 ( .S(n3), .A0(n186), .A1(tlvp_rsm_pt_tlv[26]), .Z(n185));
Q_AN02 U359 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[26]), .Z(n186));
Q_MX02 U360 ( .S(n3), .A0(n188), .A1(tlvp_rsm_pt_tlv[25]), .Z(n187));
Q_AN02 U361 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[25]), .Z(n188));
Q_MX02 U362 ( .S(n3), .A0(n190), .A1(tlvp_rsm_pt_tlv[24]), .Z(n189));
Q_AN02 U363 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[24]), .Z(n190));
Q_MX02 U364 ( .S(n3), .A0(n192), .A1(tlvp_rsm_pt_tlv[23]), .Z(n191));
Q_AN02 U365 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[23]), .Z(n192));
Q_MX02 U366 ( .S(n3), .A0(n194), .A1(tlvp_rsm_pt_tlv[22]), .Z(n193));
Q_AN02 U367 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[22]), .Z(n194));
Q_MX02 U368 ( .S(n3), .A0(n196), .A1(tlvp_rsm_pt_tlv[21]), .Z(n195));
Q_AN02 U369 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[21]), .Z(n196));
Q_MX02 U370 ( .S(n3), .A0(n198), .A1(tlvp_rsm_pt_tlv[20]), .Z(n197));
Q_AN02 U371 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[20]), .Z(n198));
Q_MX02 U372 ( .S(n3), .A0(n200), .A1(tlvp_rsm_pt_tlv[19]), .Z(n199));
Q_AN02 U373 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[19]), .Z(n200));
Q_MX02 U374 ( .S(n3), .A0(n202), .A1(tlvp_rsm_pt_tlv[18]), .Z(n201));
Q_AN02 U375 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[18]), .Z(n202));
Q_MX02 U376 ( .S(n3), .A0(n204), .A1(tlvp_rsm_pt_tlv[17]), .Z(n203));
Q_AN02 U377 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[17]), .Z(n204));
Q_MX02 U378 ( .S(n3), .A0(n206), .A1(tlvp_rsm_pt_tlv[16]), .Z(n205));
Q_AN02 U379 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[16]), .Z(n206));
Q_MX02 U380 ( .S(n3), .A0(n208), .A1(tlvp_rsm_pt_tlv[15]), .Z(n207));
Q_AN02 U381 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[15]), .Z(n208));
Q_MX02 U382 ( .S(n3), .A0(n210), .A1(tlvp_rsm_pt_tlv[14]), .Z(n209));
Q_AN02 U383 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[14]), .Z(n210));
Q_MX02 U384 ( .S(n3), .A0(n212), .A1(tlvp_rsm_pt_tlv[13]), .Z(n211));
Q_AN02 U385 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[13]), .Z(n212));
Q_MX02 U386 ( .S(n3), .A0(n214), .A1(tlvp_rsm_pt_tlv[12]), .Z(n213));
Q_AN02 U387 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[12]), .Z(n214));
Q_MX02 U388 ( .S(n3), .A0(n216), .A1(tlvp_rsm_pt_tlv[11]), .Z(n215));
Q_AN02 U389 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[11]), .Z(n216));
Q_MX02 U390 ( .S(n3), .A0(n218), .A1(tlvp_rsm_pt_tlv[10]), .Z(n217));
Q_AN02 U391 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[10]), .Z(n218));
Q_MX02 U392 ( .S(n3), .A0(n220), .A1(tlvp_rsm_pt_tlv[9]), .Z(n219));
Q_AN02 U393 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[9]), .Z(n220));
Q_MX02 U394 ( .S(n3), .A0(n222), .A1(tlvp_rsm_pt_tlv[8]), .Z(n221));
Q_AN02 U395 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[8]), .Z(n222));
Q_MX02 U396 ( .S(n3), .A0(n224), .A1(tlvp_rsm_pt_tlv[7]), .Z(n223));
Q_AN02 U397 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[7]), .Z(n224));
Q_MX02 U398 ( .S(n3), .A0(n226), .A1(tlvp_rsm_pt_tlv[6]), .Z(n225));
Q_AN02 U399 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[6]), .Z(n226));
Q_MX02 U400 ( .S(n3), .A0(n228), .A1(tlvp_rsm_pt_tlv[5]), .Z(n227));
Q_AN02 U401 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[5]), .Z(n228));
Q_MX02 U402 ( .S(n3), .A0(n230), .A1(tlvp_rsm_pt_tlv[4]), .Z(n229));
Q_AN02 U403 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[4]), .Z(n230));
Q_MX02 U404 ( .S(n3), .A0(n232), .A1(tlvp_rsm_pt_tlv[3]), .Z(n231));
Q_AN02 U405 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[3]), .Z(n232));
Q_MX02 U406 ( .S(n3), .A0(n234), .A1(tlvp_rsm_pt_tlv[2]), .Z(n233));
Q_AN02 U407 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[2]), .Z(n234));
Q_MX02 U408 ( .S(n3), .A0(n236), .A1(tlvp_rsm_pt_tlv[1]), .Z(n235));
Q_AN02 U409 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[1]), .Z(n236));
Q_MX02 U410 ( .S(n3), .A0(n238), .A1(tlvp_rsm_pt_tlv[0]), .Z(n237));
Q_AN02 U411 ( .A0(n4), .A1(tlvp_rsm_usr_ob_tlv[0]), .Z(n238));
Q_AN02 U412 ( .A0(n2), .A1(n270), .Z(n239));
Q_AN02 U413 ( .A0(n2), .A1(n272), .Z(n240));
Q_AN02 U414 ( .A0(n2), .A1(n274), .Z(n241));
Q_AN02 U415 ( .A0(n2), .A1(n276), .Z(n242));
Q_AN02 U416 ( .A0(n2), .A1(n278), .Z(n243));
Q_AN02 U417 ( .A0(n2), .A1(n280), .Z(n244));
Q_AN02 U418 ( .A0(n2), .A1(n282), .Z(n245));
Q_AN02 U419 ( .A0(n2), .A1(n284), .Z(n246));
Q_AN02 U420 ( .A0(n2), .A1(n286), .Z(n247));
Q_AN02 U421 ( .A0(n2), .A1(n288), .Z(n248));
Q_AN02 U422 ( .A0(n2), .A1(n290), .Z(n249));
Q_AN02 U423 ( .A0(n2), .A1(n292), .Z(n250));
Q_ND02 U424 ( .A0(n2), .A1(n305), .Z(n251));
Q_MX02 U425 ( .S(n3), .A0(n253), .A1(tlvp_rsm_pt_tlv[91]), .Z(n252));
Q_OR02 U426 ( .A0(n268), .A1(tlvp_rsm_usr_ob_tlv[91]), .Z(n253));
Q_MX02 U427 ( .S(n3), .A0(n255), .A1(tlvp_rsm_pt_tlv[90]), .Z(n254));
Q_OR02 U428 ( .A0(n268), .A1(tlvp_rsm_usr_ob_tlv[90]), .Z(n255));
Q_MX02 U429 ( .S(n3), .A0(n257), .A1(tlvp_rsm_pt_tlv[89]), .Z(n256));
Q_OR02 U430 ( .A0(n268), .A1(tlvp_rsm_usr_ob_tlv[89]), .Z(n257));
Q_MX02 U431 ( .S(n3), .A0(n259), .A1(tlvp_rsm_pt_tlv[88]), .Z(n258));
Q_OR02 U432 ( .A0(n268), .A1(tlvp_rsm_usr_ob_tlv[88]), .Z(n259));
Q_MX02 U433 ( .S(n3), .A0(n261), .A1(tlvp_rsm_pt_tlv[87]), .Z(n260));
Q_OR02 U434 ( .A0(n268), .A1(tlvp_rsm_usr_ob_tlv[87]), .Z(n261));
Q_MX02 U435 ( .S(n3), .A0(n263), .A1(tlvp_rsm_pt_tlv[86]), .Z(n262));
Q_OR02 U436 ( .A0(n268), .A1(tlvp_rsm_usr_ob_tlv[86]), .Z(n263));
Q_MX02 U437 ( .S(n3), .A0(n265), .A1(tlvp_rsm_pt_tlv[85]), .Z(n264));
Q_OR02 U438 ( .A0(n268), .A1(tlvp_rsm_usr_ob_tlv[85]), .Z(n265));
Q_MX02 U439 ( .S(n3), .A0(n267), .A1(tlvp_rsm_pt_tlv[84]), .Z(n266));
Q_OR02 U440 ( .A0(n268), .A1(tlvp_rsm_usr_ob_tlv[84]), .Z(n267));
Q_INV U441 ( .A(n4), .Z(n268));
Q_AN02 U442 ( .A0(n5), .A1(tlvp_rsm_usr_ob_tlv[105]), .Z(n269));
Q_XOR2 U443 ( .A0(n271), .A1(n293), .Z(n270));
Q_AD01HF U444 ( .A0(n273), .B0(n294), .S(n272), .CO(n271));
Q_AD01HF U445 ( .A0(n275), .B0(n295), .S(n274), .CO(n273));
Q_AD01HF U446 ( .A0(n277), .B0(n296), .S(n276), .CO(n275));
Q_AD01HF U447 ( .A0(n279), .B0(n297), .S(n278), .CO(n277));
Q_AD01HF U448 ( .A0(n281), .B0(n298), .S(n280), .CO(n279));
Q_AD01HF U449 ( .A0(n283), .B0(n299), .S(n282), .CO(n281));
Q_AD01HF U450 ( .A0(n285), .B0(n300), .S(n284), .CO(n283));
Q_AD01HF U451 ( .A0(n287), .B0(n301), .S(n286), .CO(n285));
Q_AD01HF U452 ( .A0(n289), .B0(n302), .S(n288), .CO(n287));
Q_AD01HF U453 ( .A0(n291), .B0(n303), .S(n290), .CO(n289));
Q_AD01HF U454 ( .A0(n304), .B0(n305), .S(n292), .CO(n291));
Q_MX02 U455 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[12]), .A1(tlvp_rsm_pt_tlv_ordern[12]), .Z(n293));
Q_MX02 U456 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[11]), .A1(tlvp_rsm_pt_tlv_ordern[11]), .Z(n294));
Q_MX02 U457 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[10]), .A1(tlvp_rsm_pt_tlv_ordern[10]), .Z(n295));
Q_MX02 U458 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[9]), .A1(tlvp_rsm_pt_tlv_ordern[9]), .Z(n296));
Q_MX02 U459 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[8]), .A1(tlvp_rsm_pt_tlv_ordern[8]), .Z(n297));
Q_MX02 U460 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[7]), .A1(tlvp_rsm_pt_tlv_ordern[7]), .Z(n298));
Q_MX02 U461 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[6]), .A1(tlvp_rsm_pt_tlv_ordern[6]), .Z(n299));
Q_MX02 U462 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[5]), .A1(tlvp_rsm_pt_tlv_ordern[5]), .Z(n300));
Q_MX02 U463 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[4]), .A1(tlvp_rsm_pt_tlv_ordern[4]), .Z(n301));
Q_MX02 U464 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[3]), .A1(tlvp_rsm_pt_tlv_ordern[3]), .Z(n302));
Q_MX02 U465 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[2]), .A1(tlvp_rsm_pt_tlv_ordern[2]), .Z(n303));
Q_MX02 U466 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[1]), .A1(tlvp_rsm_pt_tlv_ordern[1]), .Z(n304));
Q_MX02 U467 ( .S(n3), .A0(tlvp_rsm_usr_ob_tlv_ordern[0]), .A1(tlvp_rsm_pt_tlv_ordern[0]), .Z(n305));
Q_FDP1 \current_state_REG[31] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[31]), .QN( ));
Q_FDP1 \current_state_REG[30] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[30]), .QN( ));
Q_FDP1 \current_state_REG[29] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[29]), .QN( ));
Q_FDP1 \current_state_REG[28] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[28]), .QN( ));
Q_FDP1 \current_state_REG[27] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[27]), .QN( ));
Q_FDP1 \current_state_REG[26] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[26]), .QN( ));
Q_FDP1 \current_state_REG[25] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[25]), .QN( ));
Q_FDP1 \current_state_REG[24] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[24]), .QN( ));
Q_FDP1 \current_state_REG[23] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[23]), .QN( ));
Q_FDP1 \current_state_REG[22] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[22]), .QN( ));
Q_FDP1 \current_state_REG[21] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[21]), .QN( ));
Q_FDP1 \current_state_REG[20] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[20]), .QN( ));
Q_FDP1 \current_state_REG[19] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[19]), .QN( ));
Q_FDP1 \current_state_REG[18] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[18]), .QN( ));
Q_FDP1 \current_state_REG[17] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[17]), .QN( ));
Q_FDP1 \current_state_REG[16] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[16]), .QN( ));
Q_FDP1 \current_state_REG[15] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[15]), .QN( ));
Q_FDP1 \current_state_REG[14] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[14]), .QN( ));
Q_FDP1 \current_state_REG[13] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[13]), .QN( ));
Q_FDP1 \current_state_REG[12] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[12]), .QN( ));
Q_FDP1 \current_state_REG[11] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[11]), .QN( ));
Q_FDP1 \current_state_REG[10] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[10]), .QN( ));
Q_FDP1 \current_state_REG[9] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[9]), .QN( ));
Q_FDP1 \current_state_REG[8] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[8]), .QN( ));
Q_FDP1 \current_state_REG[7] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[7]), .QN( ));
Q_FDP1 \current_state_REG[6] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[6]), .QN( ));
Q_FDP1 \current_state_REG[5] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[5]), .QN( ));
Q_FDP1 \current_state_REG[4] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[4]), .QN( ));
Q_FDP1 \current_state_REG[3] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[3]), .QN( ));
Q_FDP1 \current_state_REG[2] ( .CK(clk), .R(rst_n), .D(next_state[2]), .Q(current_state[2]), .QN( ));
Q_FDP1 \current_state_REG[1] ( .CK(clk), .R(rst_n), .D(next_state[1]), .Q(current_state[1]), .QN(n310));
Q_FDP1 \current_state_REG[0] ( .CK(clk), .R(rst_n), .D(next_state[0]), .Q(current_state[0]), .QN(n342));
Q_OA21 U500 ( .A0(n307), .A1(n308), .B0(n306), .Z(next_state[0]));
Q_AN03 U501 ( .A0(n310), .A1(n311), .A2(n309), .Z(n307));
Q_AN03 U502 ( .A0(n313), .A1(tlvp_rsm_ob_datain[82]), .A2(n311), .Z(n312));
Q_AN02 U503 ( .A0(n314), .A1(tlvp_rsm_pt_sel), .Z(n311));
Q_INV U504 ( .A(tlvp_rsm_usr_ob_sel), .Z(n314));
Q_AO21 U505 ( .A0(n315), .A1(n316), .B0(n312), .Z(n308));
Q_AN02 U506 ( .A0(n310), .A1(current_state[0]), .Z(n315));
Q_AN02 U507 ( .A0(n319), .A1(n320), .Z(n318));
Q_NR02 U508 ( .A0(current_state[3]), .A1(current_state[2]), .Z(n320));
Q_NR02 U509 ( .A0(current_state[5]), .A1(current_state[4]), .Z(n319));
Q_AN03 U510 ( .A0(n321), .A1(n322), .A2(n318), .Z(n317));
Q_AN02 U511 ( .A0(n323), .A1(n324), .Z(n322));
Q_NR02 U512 ( .A0(current_state[7]), .A1(current_state[6]), .Z(n324));
Q_NR02 U513 ( .A0(current_state[9]), .A1(current_state[8]), .Z(n323));
Q_AN02 U514 ( .A0(n325), .A1(n326), .Z(n321));
Q_NR02 U515 ( .A0(current_state[11]), .A1(current_state[10]), .Z(n326));
Q_NR02 U516 ( .A0(current_state[13]), .A1(current_state[12]), .Z(n325));
Q_AN03 U517 ( .A0(n327), .A1(n328), .A2(n317), .Z(n306));
Q_AN02 U518 ( .A0(n330), .A1(n331), .Z(n329));
Q_NR02 U519 ( .A0(current_state[15]), .A1(current_state[14]), .Z(n331));
Q_NR02 U520 ( .A0(current_state[17]), .A1(current_state[16]), .Z(n330));
Q_AN03 U521 ( .A0(n332), .A1(n333), .A2(n329), .Z(n328));
Q_NR02 U522 ( .A0(current_state[19]), .A1(current_state[18]), .Z(n333));
Q_NR02 U523 ( .A0(current_state[21]), .A1(current_state[20]), .Z(n332));
Q_AN03 U524 ( .A0(n335), .A1(n336), .A2(n337), .Z(n334));
Q_NR02 U525 ( .A0(current_state[23]), .A1(current_state[22]), .Z(n336));
Q_NR02 U526 ( .A0(current_state[25]), .A1(current_state[24]), .Z(n335));
Q_NR02 U527 ( .A0(current_state[27]), .A1(current_state[26]), .Z(n337));
Q_AN03 U528 ( .A0(n338), .A1(n339), .A2(n334), .Z(n327));
Q_NR02 U529 ( .A0(current_state[29]), .A1(current_state[28]), .Z(n339));
Q_NR02 U530 ( .A0(current_state[31]), .A1(current_state[30]), .Z(n338));
Q_OA21 U531 ( .A0(n340), .A1(n341), .B0(n306), .Z(next_state[1]));
Q_AN02 U532 ( .A0(current_state[1]), .A1(n342), .Z(n313));
Q_AN03 U533 ( .A0(n310), .A1(tlvp_rsm_usr_ob_sel), .A2(n309), .Z(n340));
Q_OA21 U534 ( .A0(n343), .A1(n316), .B0(n313), .Z(n341));
Q_AN02 U535 ( .A0(tlvp_rsm_usr_ob_sel), .A1(tlvp_rsm_ob_datain[82]), .Z(n343));
Q_AO21 U536 ( .A0(current_state[0]), .A1(tlvp_rsm_ob_datain[82]), .B0(n342), .Z(n309));
Q_OR03 U537 ( .A0(tlvp_rsm_usr_ob_next), .A1(tlvp_rsm_usr_insert), .A2(n346), .Z(n347));
Q_AN03 U538 ( .A0(tlvp_rsm_selector[0]), .A1(n456), .A2(n345), .Z(n346));
Q_INV U539 ( .A(n344), .Z(n345));
Q_AN02 U540 ( .A0(tlvp_rsm_selector[1]), .A1(n347), .Z(tlvp_rsm_usr_ob_sel));
Q_AO21 U541 ( .A0(tlvp_rsm_selector[1]), .A1(n344), .B0(tlvp_rsm_pt_next), .Z(n349));
Q_NR02 U542 ( .A0(tlvp_rsm_selector[1]), .A1(n456), .Z(n350));
Q_INV U543 ( .A(tlvp_rsm_usr_ob_next), .Z(n348));
Q_AO21 U544 ( .A0(n349), .A1(n348), .B0(n350), .Z(n352));
Q_AN03 U545 ( .A0(tlvp_rsm_selector[0]), .A1(n351), .A2(n352), .Z(tlvp_rsm_pt_sel));
Q_OR03 U546 ( .A0(n388), .A1(n353), .A2(n354), .Z(n344));
Q_AO21 U547 ( .A0(n356), .A1(n360), .B0(n355), .Z(n354));
Q_AN03 U548 ( .A0(n356), .A1(n359), .A2(n357), .Z(n355));
Q_AN02 U549 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[0]), .A1(n358), .Z(n357));
Q_OR03 U550 ( .A0(n371), .A1(n361), .A2(n362), .Z(n360));
Q_AO21 U551 ( .A0(n365), .A1(n367), .B0(n363), .Z(n362));
Q_OA21 U552 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[1]), .A1(n366), .B0(n364), .Z(n359));
Q_AN03 U553 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[1]), .A1(n366), .A2(n364), .Z(n363));
Q_OA21 U554 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[2]), .A1(n368), .B0(n365), .Z(n364));
Q_AN02 U555 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[2]), .A1(n368), .Z(n367));
Q_OA21 U556 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[3]), .A1(n369), .B0(n370), .Z(n365));
Q_AN03 U557 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[3]), .A1(n369), .A2(n370), .Z(n361));
Q_OR02 U558 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[4]), .A1(n372), .Z(n370));
Q_AN02 U559 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[4]), .A1(n372), .Z(n371));
Q_AN03 U560 ( .A0(n376), .A1(n378), .A2(n387), .Z(n356));
Q_OA21 U561 ( .A0(n373), .A1(n374), .B0(n387), .Z(n353));
Q_AO21 U562 ( .A0(n384), .A1(n382), .B0(n385), .Z(n373));
Q_AO21 U563 ( .A0(n377), .A1(n380), .B0(n375), .Z(n374));
Q_OR02 U564 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[5]), .A1(n379), .Z(n378));
Q_AN03 U565 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[5]), .A1(n379), .A2(n376), .Z(n375));
Q_OA21 U566 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[6]), .A1(n381), .B0(n377), .Z(n376));
Q_AN02 U567 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[6]), .A1(n381), .Z(n380));
Q_OA21 U568 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[7]), .A1(n383), .B0(n384), .Z(n377));
Q_AN02 U569 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[7]), .A1(n383), .Z(n382));
Q_OR02 U570 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[8]), .A1(n386), .Z(n384));
Q_AN02 U571 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[8]), .A1(n386), .Z(n385));
Q_OR03 U572 ( .A0(n399), .A1(n389), .A2(n390), .Z(n388));
Q_AO21 U573 ( .A0(n393), .A1(n395), .B0(n391), .Z(n390));
Q_OA21 U574 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[9]), .A1(n394), .B0(n392), .Z(n387));
Q_AN03 U575 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[9]), .A1(n394), .A2(n392), .Z(n391));
Q_OA21 U576 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[10]), .A1(n396), .B0(n393), .Z(n392));
Q_AN02 U577 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[10]), .A1(n396), .Z(n395));
Q_OA21 U578 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[11]), .A1(n397), .B0(n398), .Z(n393));
Q_AN03 U579 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[11]), .A1(n397), .A2(n398), .Z(n389));
Q_OR02 U580 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[12]), .A1(n400), .Z(n398));
Q_AN02 U581 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[12]), .A1(n400), .Z(n399));
Q_AN02 U582 ( .A0(tlvp_rsm_usr_ob_ren), .A1(n404), .Z(n402));
Q_INV U583 ( .A(tlvp_rsm_pt_wen), .Z(n405));
Q_XOR2 U584 ( .A0(pt_ob_rd), .A1(n405), .Z(n406));
Q_INV U585 ( .A(tlvp_rsm_usr_ob_wen), .Z(n403));
Q_XOR2 U586 ( .A0(tlvp_rsm_usr_ob_ren), .A1(n403), .Z(n407));
Q_MX02 U587 ( .S(n404), .A0(tlvp_rsm_usr_ob_rdata[63]), .A1(tlvp_rsm_bip2[1]), .Z(n408));
Q_MX02 U588 ( .S(n404), .A0(tlvp_rsm_usr_ob_rdata[62]), .A1(tlvp_rsm_bip2[0]), .Z(n409));
Q_OA21 U589 ( .A0(pt_ob_tlv[83]), .A1(pt_ob_tlv[64]), .B0(pt_ob_rd), .Z(n401));
Q_OR02 U590 ( .A0(tlvp_rsm_usr_ob_rdata[83]), .A1(tlvp_rsm_usr_ob_rdata[64]), .Z(n404));
ixc_assign_64 _zz_strnp_0 ( tlvp_rsm_usr_ob_rdata_dw0[63:0], 
	tlvp_rsm_usr_ob_rdata[63:0]);
Q_AN02 U592 ( .A0(tlvp_rsm_pt_valid), .A1(n3), .Z(tlvp_rsm_pt_wen));
Q_INV U593 ( .A(usr_ob_empty), .Z(n511));
Q_INV U594 ( .A(tlvp_ob_afull), .Z(n510));
Q_OR02 U595 ( .A0(n509), .A1(tlvp_rsm_usr_ob_wen), .Z(n508));
Q_AN03 U596 ( .A0(n511), .A1(n510), .A2(n508), .Z(tlvp_rsm_usr_ob_ren));
Q_INV U597 ( .A(pt_ob_empty), .Z(n507));
Q_OR02 U598 ( .A0(n506), .A1(tlvp_rsm_pt_wen), .Z(n505));
Q_AN03 U599 ( .A0(n507), .A1(n510), .A2(n505), .Z(pt_ob_rd));
Q_AN02 U600 ( .A0(tlvp_rsm_pt_tlv_ordern[12]), .A1(n504), .Z(n503));
Q_OR02 U601 ( .A0(tlvp_rsm_pt_tlv_ordern[12]), .A1(n504), .Z(n502));
Q_AN03 U602 ( .A0(tlvp_rsm_pt_tlv_ordern[11]), .A1(n501), .A2(n502), .Z(n493));
Q_OA21 U603 ( .A0(tlvp_rsm_pt_tlv_ordern[11]), .A1(n501), .B0(n502), .Z(n497));
Q_AN02 U604 ( .A0(tlvp_rsm_pt_tlv_ordern[10]), .A1(n500), .Z(n499));
Q_OA21 U605 ( .A0(tlvp_rsm_pt_tlv_ordern[10]), .A1(n500), .B0(n497), .Z(n496));
Q_AN03 U606 ( .A0(tlvp_rsm_pt_tlv_ordern[9]), .A1(n498), .A2(n496), .Z(n495));
Q_OA21 U607 ( .A0(tlvp_rsm_pt_tlv_ordern[9]), .A1(n498), .B0(n496), .Z(n491));
Q_AO21 U608 ( .A0(n497), .A1(n499), .B0(n495), .Z(n494));
Q_OR03 U609 ( .A0(n503), .A1(n493), .A2(n494), .Z(n492));
Q_AN02 U610 ( .A0(tlvp_rsm_pt_tlv_ordern[8]), .A1(n490), .Z(n489));
Q_OR02 U611 ( .A0(tlvp_rsm_pt_tlv_ordern[8]), .A1(n490), .Z(n488));
Q_AN02 U612 ( .A0(tlvp_rsm_pt_tlv_ordern[7]), .A1(n487), .Z(n486));
Q_OA21 U613 ( .A0(tlvp_rsm_pt_tlv_ordern[7]), .A1(n487), .B0(n488), .Z(n481));
Q_AN02 U614 ( .A0(tlvp_rsm_pt_tlv_ordern[6]), .A1(n485), .Z(n484));
Q_OA21 U615 ( .A0(tlvp_rsm_pt_tlv_ordern[6]), .A1(n485), .B0(n481), .Z(n480));
Q_AN03 U616 ( .A0(tlvp_rsm_pt_tlv_ordern[5]), .A1(n483), .A2(n480), .Z(n479));
Q_OR02 U617 ( .A0(tlvp_rsm_pt_tlv_ordern[5]), .A1(n483), .Z(n482));
Q_AO21 U618 ( .A0(n481), .A1(n484), .B0(n479), .Z(n478));
Q_AO21 U619 ( .A0(n488), .A1(n486), .B0(n489), .Z(n477));
Q_OA21 U620 ( .A0(n477), .A1(n478), .B0(n491), .Z(n457));
Q_AN03 U621 ( .A0(n480), .A1(n482), .A2(n491), .Z(n460));
Q_AN02 U622 ( .A0(tlvp_rsm_pt_tlv_ordern[4]), .A1(n476), .Z(n475));
Q_OR02 U623 ( .A0(tlvp_rsm_pt_tlv_ordern[4]), .A1(n476), .Z(n474));
Q_AN03 U624 ( .A0(tlvp_rsm_pt_tlv_ordern[3]), .A1(n473), .A2(n474), .Z(n465));
Q_OA21 U625 ( .A0(tlvp_rsm_pt_tlv_ordern[3]), .A1(n473), .B0(n474), .Z(n469));
Q_AN02 U626 ( .A0(tlvp_rsm_pt_tlv_ordern[2]), .A1(n472), .Z(n471));
Q_OA21 U627 ( .A0(tlvp_rsm_pt_tlv_ordern[2]), .A1(n472), .B0(n469), .Z(n468));
Q_AN03 U628 ( .A0(tlvp_rsm_pt_tlv_ordern[1]), .A1(n470), .A2(n468), .Z(n467));
Q_OA21 U629 ( .A0(tlvp_rsm_pt_tlv_ordern[1]), .A1(n470), .B0(n468), .Z(n463));
Q_AO21 U630 ( .A0(n469), .A1(n471), .B0(n467), .Z(n466));
Q_OR03 U631 ( .A0(n475), .A1(n465), .A2(n466), .Z(n464));
Q_AN02 U632 ( .A0(tlvp_rsm_pt_tlv_ordern[0]), .A1(n462), .Z(n461));
Q_AN03 U633 ( .A0(n460), .A1(n463), .A2(n461), .Z(n459));
Q_AO21 U634 ( .A0(n460), .A1(n464), .B0(n459), .Z(n458));
Q_OR03 U635 ( .A0(n492), .A1(n457), .A2(n458), .Z(n456));
Q_INV U636 ( .A(n456), .Z(tlvp_rsm_pt_next));
Q_XNR2 U637 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[0]), .A1(tlvp_rsm_nxt_ordern[0]), .Z(n455));
Q_XNR2 U638 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[1]), .A1(tlvp_rsm_nxt_ordern[1]), .Z(n454));
Q_XNR2 U639 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[2]), .A1(tlvp_rsm_nxt_ordern[2]), .Z(n453));
Q_XNR2 U640 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[3]), .A1(tlvp_rsm_nxt_ordern[3]), .Z(n452));
Q_XNR2 U641 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[4]), .A1(tlvp_rsm_nxt_ordern[4]), .Z(n451));
Q_XNR2 U642 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[5]), .A1(tlvp_rsm_nxt_ordern[5]), .Z(n450));
Q_XNR2 U643 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[6]), .A1(tlvp_rsm_nxt_ordern[6]), .Z(n449));
Q_XNR2 U644 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[7]), .A1(tlvp_rsm_nxt_ordern[7]), .Z(n448));
Q_XNR2 U645 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[8]), .A1(tlvp_rsm_nxt_ordern[8]), .Z(n447));
Q_XNR2 U646 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[9]), .A1(tlvp_rsm_nxt_ordern[9]), .Z(n446));
Q_XNR2 U647 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[10]), .A1(tlvp_rsm_nxt_ordern[10]), .Z(n445));
Q_XNR2 U648 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[11]), .A1(tlvp_rsm_nxt_ordern[11]), .Z(n444));
Q_XNR2 U649 ( .A0(tlvp_rsm_usr_ob_tlv_ordern[12]), .A1(tlvp_rsm_nxt_ordern[12]), .Z(n443));
Q_AN03 U650 ( .A0(n443), .A1(n444), .A2(n445), .Z(n442));
Q_AN03 U651 ( .A0(n446), .A1(n447), .A2(n448), .Z(n441));
Q_AN03 U652 ( .A0(n449), .A1(n450), .A2(n451), .Z(n440));
Q_AN03 U653 ( .A0(n452), .A1(n453), .A2(n454), .Z(n439));
Q_AN03 U654 ( .A0(n455), .A1(n442), .A2(n441), .Z(n438));
Q_AN03 U655 ( .A0(n440), .A1(n439), .A2(n438), .Z(tlvp_rsm_usr_ob_next));
ixc_assign_2 _zz_strnp_1 ( tlvp_rsm_selector[1:0], { tlvp_rsm_usr_ob_valid, 
	tlvp_rsm_pt_valid});
ixc_assign _zz_strnp_2 ( tlvp_rsm_ob_wdata[82], tlvp_rsm_ob_wen);
ixc_assign _zz_strnp_4 ( tlvp_rsm_ob_wdata[80], tlvp_rsm_ob_datain[80]);
ixc_assign_8 _zz_strnp_5 ( tlvp_rsm_ob_wdata[79:72], 
	tlvp_rsm_ob_datain[79:72]);
ixc_assign_8 _zz_strnp_6 ( tlvp_rsm_ob_wdata[71:64], 
	tlvp_rsm_ob_datain[71:64]);
ixc_assign_64 _zz_strnp_7 ( tlvp_rsm_ob_wdata[63:0], 
	tlvp_rsm_ob_datain[63:0]);
ixc_assign _zz_strnp_8 ( _zy_simnet_pt_ob_rd_0_w$, pt_ob_rd);
ixc_assign _zz_strnp_9 ( _zy_simnet_tlvp_rsm_usr_ob_ren_1_w$, 
	tlvp_rsm_usr_ob_ren);
ixc_assign _zz_strnp_10 ( _zy_simnet_tlvp_rsm_ob_wen_2_w$, tlvp_rsm_ob_wen);
ixc_assign_83 _zz_strnp_11 ( _zy_simnet_tlvp_rsm_ob_wdata_3_w$[0:82], 
	tlvp_rsm_ob_wdata[82:0]);
ixc_assign _zz_strnp_3 ( tlvp_rsm_ob_wdata[81], tlvp_rsm_ob_datain[81]);
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[105] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[105]), .Q(tlvp_rsm_pt_tlv[105]));
Q_INV U668 ( .A(rst_n), .Z(n512));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[104] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[104]), .Q(tlvp_rsm_pt_tlv[104]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[103] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[103]), .Q(tlvp_rsm_pt_tlv[103]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[102] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[102]), .Q(tlvp_rsm_pt_tlv[102]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[101] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[101]), .Q(tlvp_rsm_pt_tlv[101]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[100] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[100]), .Q(tlvp_rsm_pt_tlv[100]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[99] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[99]), .Q(tlvp_rsm_pt_tlv[99]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[98] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[98]), .Q(tlvp_rsm_pt_tlv[98]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[97] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[97]), .Q(tlvp_rsm_pt_tlv[97]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[96] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[96]), .Q(tlvp_rsm_pt_tlv[96]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[95] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[95]), .Q(tlvp_rsm_pt_tlv[95]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[94] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[94]), .Q(tlvp_rsm_pt_tlv[94]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[93] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[93]), .Q(tlvp_rsm_pt_tlv[93]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[92] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[92]), .Q(tlvp_rsm_pt_tlv[92]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[91] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[91]), .Q(tlvp_rsm_pt_tlv[91]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[90] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[90]), .Q(tlvp_rsm_pt_tlv[90]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[89] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[89]), .Q(tlvp_rsm_pt_tlv[89]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[88] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[88]), .Q(tlvp_rsm_pt_tlv[88]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[87] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[87]), .Q(tlvp_rsm_pt_tlv[87]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[86] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[86]), .Q(tlvp_rsm_pt_tlv[86]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[85] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[85]), .Q(tlvp_rsm_pt_tlv[85]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[84] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[84]), .Q(tlvp_rsm_pt_tlv[84]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[83] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[83]), .Q(tlvp_rsm_pt_tlv[83]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[82] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[82]), .Q(tlvp_rsm_pt_tlv[82]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[81] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[81]), .Q(tlvp_rsm_pt_tlv[81]));
Q_INV U693 ( .A(tlvp_rsm_pt_tlv[81]), .Z(n14));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[80] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[80]), .Q(tlvp_rsm_pt_tlv[80]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[79] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[79]), .Q(tlvp_rsm_pt_tlv[79]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[78] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[78]), .Q(tlvp_rsm_pt_tlv[78]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[77] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[77]), .Q(tlvp_rsm_pt_tlv[77]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[76] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[76]), .Q(tlvp_rsm_pt_tlv[76]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[75] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[75]), .Q(tlvp_rsm_pt_tlv[75]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[74] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[74]), .Q(tlvp_rsm_pt_tlv[74]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[73] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[73]), .Q(tlvp_rsm_pt_tlv[73]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[72] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[72]), .Q(tlvp_rsm_pt_tlv[72]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[71] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[71]), .Q(tlvp_rsm_pt_tlv[71]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[70] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[70]), .Q(tlvp_rsm_pt_tlv[70]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[69] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[69]), .Q(tlvp_rsm_pt_tlv[69]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[68] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[68]), .Q(tlvp_rsm_pt_tlv[68]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[67] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[67]), .Q(tlvp_rsm_pt_tlv[67]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[66] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[66]), .Q(tlvp_rsm_pt_tlv[66]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[65] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[65]), .Q(tlvp_rsm_pt_tlv[65]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[64] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[64]), .Q(tlvp_rsm_pt_tlv[64]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[63] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[63]), .Q(tlvp_rsm_pt_tlv[63]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[62] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[62]), .Q(tlvp_rsm_pt_tlv[62]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[61] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[61]), .Q(tlvp_rsm_pt_tlv[61]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[60] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[60]), .Q(tlvp_rsm_pt_tlv[60]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[59] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[59]), .Q(tlvp_rsm_pt_tlv[59]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[58] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[58]), .Q(tlvp_rsm_pt_tlv[58]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[57] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[57]), .Q(tlvp_rsm_pt_tlv[57]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[56] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[56]), .Q(tlvp_rsm_pt_tlv[56]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[55] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[55]), .Q(tlvp_rsm_pt_tlv[55]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[54] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[54]), .Q(tlvp_rsm_pt_tlv[54]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[53] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[53]), .Q(tlvp_rsm_pt_tlv[53]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[52] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[52]), .Q(tlvp_rsm_pt_tlv[52]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[51] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[51]), .Q(tlvp_rsm_pt_tlv[51]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[50] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[50]), .Q(tlvp_rsm_pt_tlv[50]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[49] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[49]), .Q(tlvp_rsm_pt_tlv[49]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[48] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[48]), .Q(tlvp_rsm_pt_tlv[48]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[47] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[47]), .Q(tlvp_rsm_pt_tlv[47]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[46] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[46]), .Q(tlvp_rsm_pt_tlv[46]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[45] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[45]), .Q(tlvp_rsm_pt_tlv[45]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[44] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[44]), .Q(tlvp_rsm_pt_tlv[44]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[43] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[43]), .Q(tlvp_rsm_pt_tlv[43]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[42] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[42]), .Q(tlvp_rsm_pt_tlv[42]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[41] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[41]), .Q(tlvp_rsm_pt_tlv[41]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[40] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[40]), .Q(tlvp_rsm_pt_tlv[40]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[39] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[39]), .Q(tlvp_rsm_pt_tlv[39]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[38] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[38]), .Q(tlvp_rsm_pt_tlv[38]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[37] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[37]), .Q(tlvp_rsm_pt_tlv[37]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[36] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[36]), .Q(tlvp_rsm_pt_tlv[36]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[35] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[35]), .Q(tlvp_rsm_pt_tlv[35]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[34] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[34]), .Q(tlvp_rsm_pt_tlv[34]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[33] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[33]), .Q(tlvp_rsm_pt_tlv[33]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[32] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[32]), .Q(tlvp_rsm_pt_tlv[32]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[31] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[31]), .Q(tlvp_rsm_pt_tlv[31]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[30] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[30]), .Q(tlvp_rsm_pt_tlv[30]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[29] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[29]), .Q(tlvp_rsm_pt_tlv[29]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[28] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[28]), .Q(tlvp_rsm_pt_tlv[28]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[27] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[27]), .Q(tlvp_rsm_pt_tlv[27]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[26] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[26]), .Q(tlvp_rsm_pt_tlv[26]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[25] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[25]), .Q(tlvp_rsm_pt_tlv[25]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[24] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[24]), .Q(tlvp_rsm_pt_tlv[24]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[23] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[23]), .Q(tlvp_rsm_pt_tlv[23]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[22] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[22]), .Q(tlvp_rsm_pt_tlv[22]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[21] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[21]), .Q(tlvp_rsm_pt_tlv[21]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[20] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[20]), .Q(tlvp_rsm_pt_tlv[20]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[19] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[19]), .Q(tlvp_rsm_pt_tlv[19]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[18] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[18]), .Q(tlvp_rsm_pt_tlv[18]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[17] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[17]), .Q(tlvp_rsm_pt_tlv[17]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[16] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[16]), .Q(tlvp_rsm_pt_tlv[16]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[15] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[15]), .Q(tlvp_rsm_pt_tlv[15]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[14] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[14]), .Q(tlvp_rsm_pt_tlv[14]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[13] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[13]), .Q(tlvp_rsm_pt_tlv[13]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[12] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[12]), .Q(tlvp_rsm_pt_tlv[12]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[11] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[11]), .Q(tlvp_rsm_pt_tlv[11]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[10] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[10]), .Q(tlvp_rsm_pt_tlv[10]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[9] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[9]), .Q(tlvp_rsm_pt_tlv[9]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[8] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[8]), .Q(tlvp_rsm_pt_tlv[8]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[7] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[7]), .Q(tlvp_rsm_pt_tlv[7]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[6] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[6]), .Q(tlvp_rsm_pt_tlv[6]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[5] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[5]), .Q(tlvp_rsm_pt_tlv[5]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[4] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[4]), .Q(tlvp_rsm_pt_tlv[4]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[3] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[3]), .Q(tlvp_rsm_pt_tlv[3]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[2] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[2]), .Q(tlvp_rsm_pt_tlv[2]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[1] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[1]), .Q(tlvp_rsm_pt_tlv[1]));
Q_FDP4EP \tlvp_rsm_pt_tlv_REG[0] ( .CK(clk), .CE(pt_ob_rd), .R(n512), .D(pt_ob_tlv[0]), .Q(tlvp_rsm_pt_tlv[0]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[12] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[104]), .Q(tlvp_rsm_usr_ob_tlv_ordern[12]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[11] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[103]), .Q(tlvp_rsm_usr_ob_tlv_ordern[11]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[10] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[102]), .Q(tlvp_rsm_usr_ob_tlv_ordern[10]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[9] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[101]), .Q(tlvp_rsm_usr_ob_tlv_ordern[9]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[8] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[100]), .Q(tlvp_rsm_usr_ob_tlv_ordern[8]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[7] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[99]), .Q(tlvp_rsm_usr_ob_tlv_ordern[7]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[6] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[98]), .Q(tlvp_rsm_usr_ob_tlv_ordern[6]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[5] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[97]), .Q(tlvp_rsm_usr_ob_tlv_ordern[5]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[4] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[96]), .Q(tlvp_rsm_usr_ob_tlv_ordern[4]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[3] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[95]), .Q(tlvp_rsm_usr_ob_tlv_ordern[3]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[2] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[94]), .Q(tlvp_rsm_usr_ob_tlv_ordern[2]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[1] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[93]), .Q(tlvp_rsm_usr_ob_tlv_ordern[1]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_ordern_REG[0] ( .CK(clk), .CE(n402), .R(n512), .D(tlvp_rsm_usr_ob_rdata[92]), .Q(tlvp_rsm_usr_ob_tlv_ordern[0]));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[12] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[104]), .Q(tlvp_rsm_pt_tlv_ordern[12]));
Q_INV U789 ( .A(tlvp_rsm_pt_tlv_ordern[12]), .Z(n400));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[11] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[103]), .Q(tlvp_rsm_pt_tlv_ordern[11]));
Q_INV U791 ( .A(tlvp_rsm_pt_tlv_ordern[11]), .Z(n397));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[10] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[102]), .Q(tlvp_rsm_pt_tlv_ordern[10]));
Q_INV U793 ( .A(tlvp_rsm_pt_tlv_ordern[10]), .Z(n396));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[9] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[101]), .Q(tlvp_rsm_pt_tlv_ordern[9]));
Q_INV U795 ( .A(tlvp_rsm_pt_tlv_ordern[9]), .Z(n394));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[8] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[100]), .Q(tlvp_rsm_pt_tlv_ordern[8]));
Q_INV U797 ( .A(tlvp_rsm_pt_tlv_ordern[8]), .Z(n386));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[7] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[99]), .Q(tlvp_rsm_pt_tlv_ordern[7]));
Q_INV U799 ( .A(tlvp_rsm_pt_tlv_ordern[7]), .Z(n383));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[6] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[98]), .Q(tlvp_rsm_pt_tlv_ordern[6]));
Q_INV U801 ( .A(tlvp_rsm_pt_tlv_ordern[6]), .Z(n381));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[5] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[97]), .Q(tlvp_rsm_pt_tlv_ordern[5]));
Q_INV U803 ( .A(tlvp_rsm_pt_tlv_ordern[5]), .Z(n379));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[4] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[96]), .Q(tlvp_rsm_pt_tlv_ordern[4]));
Q_INV U805 ( .A(tlvp_rsm_pt_tlv_ordern[4]), .Z(n372));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[3] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[95]), .Q(tlvp_rsm_pt_tlv_ordern[3]));
Q_INV U807 ( .A(tlvp_rsm_pt_tlv_ordern[3]), .Z(n369));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[2] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[94]), .Q(tlvp_rsm_pt_tlv_ordern[2]));
Q_INV U809 ( .A(tlvp_rsm_pt_tlv_ordern[2]), .Z(n368));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[1] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[93]), .Q(tlvp_rsm_pt_tlv_ordern[1]));
Q_INV U811 ( .A(tlvp_rsm_pt_tlv_ordern[1]), .Z(n366));
Q_FDP4EP \tlvp_rsm_pt_tlv_ordern_REG[0] ( .CK(clk), .CE(n401), .R(n512), .D(pt_ob_tlv[92]), .Q(tlvp_rsm_pt_tlv_ordern[0]));
Q_INV U813 ( .A(tlvp_rsm_pt_tlv_ordern[0]), .Z(n358));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[105] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[105]), .Q(tlvp_rsm_usr_ob_tlv[105]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[104] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[104]), .Q(tlvp_rsm_usr_ob_tlv[104]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[103] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[103]), .Q(tlvp_rsm_usr_ob_tlv[103]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[102] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[102]), .Q(tlvp_rsm_usr_ob_tlv[102]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[101] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[101]), .Q(tlvp_rsm_usr_ob_tlv[101]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[100] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[100]), .Q(tlvp_rsm_usr_ob_tlv[100]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[99] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[99]), .Q(tlvp_rsm_usr_ob_tlv[99]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[98] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[98]), .Q(tlvp_rsm_usr_ob_tlv[98]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[97] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[97]), .Q(tlvp_rsm_usr_ob_tlv[97]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[96] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[96]), .Q(tlvp_rsm_usr_ob_tlv[96]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[95] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[95]), .Q(tlvp_rsm_usr_ob_tlv[95]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[94] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[94]), .Q(tlvp_rsm_usr_ob_tlv[94]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[93] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[93]), .Q(tlvp_rsm_usr_ob_tlv[93]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[92] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[92]), .Q(tlvp_rsm_usr_ob_tlv[92]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[91] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[91]), .Q(tlvp_rsm_usr_ob_tlv[91]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[90] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[90]), .Q(tlvp_rsm_usr_ob_tlv[90]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[89] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[89]), .Q(tlvp_rsm_usr_ob_tlv[89]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[88] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[88]), .Q(tlvp_rsm_usr_ob_tlv[88]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[87] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[87]), .Q(tlvp_rsm_usr_ob_tlv[87]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[86] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[86]), .Q(tlvp_rsm_usr_ob_tlv[86]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[85] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[85]), .Q(tlvp_rsm_usr_ob_tlv[85]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[84] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[84]), .Q(tlvp_rsm_usr_ob_tlv[84]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[83] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[83]), .Q(tlvp_rsm_usr_ob_tlv[83]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[82] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[82]), .Q(tlvp_rsm_usr_ob_tlv[82]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[81] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[81]), .Q(tlvp_rsm_usr_ob_tlv[81]));
Q_INV U839 ( .A(tlvp_rsm_usr_ob_tlv[81]), .Z(n15));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[80] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[80]), .Q(tlvp_rsm_usr_ob_tlv[80]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[79] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[79]), .Q(tlvp_rsm_usr_ob_tlv[79]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[78] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[78]), .Q(tlvp_rsm_usr_ob_tlv[78]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[77] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[77]), .Q(tlvp_rsm_usr_ob_tlv[77]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[76] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[76]), .Q(tlvp_rsm_usr_ob_tlv[76]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[75] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[75]), .Q(tlvp_rsm_usr_ob_tlv[75]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[74] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[74]), .Q(tlvp_rsm_usr_ob_tlv[74]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[73] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[73]), .Q(tlvp_rsm_usr_ob_tlv[73]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[72] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[72]), .Q(tlvp_rsm_usr_ob_tlv[72]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[71] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[71]), .Q(tlvp_rsm_usr_ob_tlv[71]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[70] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[70]), .Q(tlvp_rsm_usr_ob_tlv[70]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[69] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[69]), .Q(tlvp_rsm_usr_ob_tlv[69]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[68] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[68]), .Q(tlvp_rsm_usr_ob_tlv[68]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[67] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[67]), .Q(tlvp_rsm_usr_ob_tlv[67]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[66] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[66]), .Q(tlvp_rsm_usr_ob_tlv[66]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[65] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[65]), .Q(tlvp_rsm_usr_ob_tlv[65]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[64] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[64]), .Q(tlvp_rsm_usr_ob_tlv[64]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[63] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(n408), .Q(tlvp_rsm_usr_ob_tlv[63]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[62] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(n409), .Q(tlvp_rsm_usr_ob_tlv[62]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[61] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[61]), .Q(tlvp_rsm_usr_ob_tlv[61]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[60] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[60]), .Q(tlvp_rsm_usr_ob_tlv[60]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[59] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[59]), .Q(tlvp_rsm_usr_ob_tlv[59]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[58] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[58]), .Q(tlvp_rsm_usr_ob_tlv[58]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[57] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[57]), .Q(tlvp_rsm_usr_ob_tlv[57]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[56] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[56]), .Q(tlvp_rsm_usr_ob_tlv[56]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[55] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[55]), .Q(tlvp_rsm_usr_ob_tlv[55]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[54] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[54]), .Q(tlvp_rsm_usr_ob_tlv[54]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[53] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[53]), .Q(tlvp_rsm_usr_ob_tlv[53]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[52] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[52]), .Q(tlvp_rsm_usr_ob_tlv[52]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[51] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[51]), .Q(tlvp_rsm_usr_ob_tlv[51]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[50] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[50]), .Q(tlvp_rsm_usr_ob_tlv[50]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[49] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[49]), .Q(tlvp_rsm_usr_ob_tlv[49]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[48] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[48]), .Q(tlvp_rsm_usr_ob_tlv[48]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[47] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[47]), .Q(tlvp_rsm_usr_ob_tlv[47]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[46] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[46]), .Q(tlvp_rsm_usr_ob_tlv[46]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[45] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[45]), .Q(tlvp_rsm_usr_ob_tlv[45]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[44] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[44]), .Q(tlvp_rsm_usr_ob_tlv[44]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[43] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[43]), .Q(tlvp_rsm_usr_ob_tlv[43]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[42] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[42]), .Q(tlvp_rsm_usr_ob_tlv[42]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[41] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[41]), .Q(tlvp_rsm_usr_ob_tlv[41]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[40] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[40]), .Q(tlvp_rsm_usr_ob_tlv[40]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[39] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[39]), .Q(tlvp_rsm_usr_ob_tlv[39]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[38] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[38]), .Q(tlvp_rsm_usr_ob_tlv[38]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[37] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[37]), .Q(tlvp_rsm_usr_ob_tlv[37]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[36] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[36]), .Q(tlvp_rsm_usr_ob_tlv[36]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[35] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[35]), .Q(tlvp_rsm_usr_ob_tlv[35]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[34] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[34]), .Q(tlvp_rsm_usr_ob_tlv[34]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[33] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[33]), .Q(tlvp_rsm_usr_ob_tlv[33]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[32] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[32]), .Q(tlvp_rsm_usr_ob_tlv[32]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[31] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[31]), .Q(tlvp_rsm_usr_ob_tlv[31]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[30] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[30]), .Q(tlvp_rsm_usr_ob_tlv[30]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[29] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[29]), .Q(tlvp_rsm_usr_ob_tlv[29]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[28] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[28]), .Q(tlvp_rsm_usr_ob_tlv[28]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[27] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[27]), .Q(tlvp_rsm_usr_ob_tlv[27]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[26] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[26]), .Q(tlvp_rsm_usr_ob_tlv[26]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[25] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[25]), .Q(tlvp_rsm_usr_ob_tlv[25]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[24] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[24]), .Q(tlvp_rsm_usr_ob_tlv[24]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[23] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[23]), .Q(tlvp_rsm_usr_ob_tlv[23]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[22] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[22]), .Q(tlvp_rsm_usr_ob_tlv[22]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[21] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[21]), .Q(tlvp_rsm_usr_ob_tlv[21]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[20] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[20]), .Q(tlvp_rsm_usr_ob_tlv[20]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[19] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[19]), .Q(tlvp_rsm_usr_ob_tlv[19]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[18] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[18]), .Q(tlvp_rsm_usr_ob_tlv[18]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[17] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[17]), .Q(tlvp_rsm_usr_ob_tlv[17]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[16] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[16]), .Q(tlvp_rsm_usr_ob_tlv[16]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[15] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[15]), .Q(tlvp_rsm_usr_ob_tlv[15]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[14] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[14]), .Q(tlvp_rsm_usr_ob_tlv[14]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[13] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[13]), .Q(tlvp_rsm_usr_ob_tlv[13]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[12] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[12]), .Q(tlvp_rsm_usr_ob_tlv[12]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[11] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[11]), .Q(tlvp_rsm_usr_ob_tlv[11]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[10] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[10]), .Q(tlvp_rsm_usr_ob_tlv[10]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[9] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[9]), .Q(tlvp_rsm_usr_ob_tlv[9]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[8] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[8]), .Q(tlvp_rsm_usr_ob_tlv[8]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[7] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[7]), .Q(tlvp_rsm_usr_ob_tlv[7]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[6] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[6]), .Q(tlvp_rsm_usr_ob_tlv[6]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[5] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[5]), .Q(tlvp_rsm_usr_ob_tlv[5]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[4] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[4]), .Q(tlvp_rsm_usr_ob_tlv[4]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[3] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[3]), .Q(tlvp_rsm_usr_ob_tlv[3]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[2] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[2]), .Q(tlvp_rsm_usr_ob_tlv[2]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[1] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[1]), .Q(tlvp_rsm_usr_ob_tlv[1]));
Q_FDP4EP \tlvp_rsm_usr_ob_tlv_REG[0] ( .CK(clk), .CE(tlvp_rsm_usr_ob_ren), .R(n512), .D(tlvp_rsm_usr_ob_rdata[0]), .Q(tlvp_rsm_usr_ob_tlv[0]));
Q_INV U921 ( .A(n407), .Z(n513));
Q_FDP4EP tlvp_rsm_usr_ob_valid_REG  ( .CK(clk), .CE(n513), .R(n512), .D(n403), .Q(tlvp_rsm_usr_ob_valid));
Q_INV U923 ( .A(tlvp_rsm_usr_ob_valid), .Z(n509));
Q_INV U924 ( .A(n406), .Z(n514));
Q_FDP4EP tlvp_rsm_pt_valid_REG  ( .CK(clk), .CE(n514), .R(n512), .D(n405), .Q(tlvp_rsm_pt_valid));
Q_INV U926 ( .A(tlvp_rsm_pt_valid), .Z(n506));
Q_INV U927 ( .A(n12), .Z(n515));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[12] ( .CK(clk), .CE(n515), .R(n512), .D(n239), .Q(tlvp_rsm_nxt_ordern[12]));
Q_INV U929 ( .A(tlvp_rsm_nxt_ordern[12]), .Z(n504));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[11] ( .CK(clk), .CE(n515), .R(n512), .D(n240), .Q(tlvp_rsm_nxt_ordern[11]));
Q_INV U931 ( .A(tlvp_rsm_nxt_ordern[11]), .Z(n501));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[10] ( .CK(clk), .CE(n515), .R(n512), .D(n241), .Q(tlvp_rsm_nxt_ordern[10]));
Q_INV U933 ( .A(tlvp_rsm_nxt_ordern[10]), .Z(n500));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[9] ( .CK(clk), .CE(n515), .R(n512), .D(n242), .Q(tlvp_rsm_nxt_ordern[9]));
Q_INV U935 ( .A(tlvp_rsm_nxt_ordern[9]), .Z(n498));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[8] ( .CK(clk), .CE(n515), .R(n512), .D(n243), .Q(tlvp_rsm_nxt_ordern[8]));
Q_INV U937 ( .A(tlvp_rsm_nxt_ordern[8]), .Z(n490));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[7] ( .CK(clk), .CE(n515), .R(n512), .D(n244), .Q(tlvp_rsm_nxt_ordern[7]));
Q_INV U939 ( .A(tlvp_rsm_nxt_ordern[7]), .Z(n487));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[6] ( .CK(clk), .CE(n515), .R(n512), .D(n245), .Q(tlvp_rsm_nxt_ordern[6]));
Q_INV U941 ( .A(tlvp_rsm_nxt_ordern[6]), .Z(n485));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[5] ( .CK(clk), .CE(n515), .R(n512), .D(n246), .Q(tlvp_rsm_nxt_ordern[5]));
Q_INV U943 ( .A(tlvp_rsm_nxt_ordern[5]), .Z(n483));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[4] ( .CK(clk), .CE(n515), .R(n512), .D(n247), .Q(tlvp_rsm_nxt_ordern[4]));
Q_INV U945 ( .A(tlvp_rsm_nxt_ordern[4]), .Z(n476));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[3] ( .CK(clk), .CE(n515), .R(n512), .D(n248), .Q(tlvp_rsm_nxt_ordern[3]));
Q_INV U947 ( .A(tlvp_rsm_nxt_ordern[3]), .Z(n473));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[2] ( .CK(clk), .CE(n515), .R(n512), .D(n249), .Q(tlvp_rsm_nxt_ordern[2]));
Q_INV U949 ( .A(tlvp_rsm_nxt_ordern[2]), .Z(n472));
Q_FDP4EP \tlvp_rsm_nxt_ordern_REG[1] ( .CK(clk), .CE(n515), .R(n512), .D(n250), .Q(tlvp_rsm_nxt_ordern[1]));
Q_INV U951 ( .A(tlvp_rsm_nxt_ordern[1]), .Z(n470));
Q_INV U952 ( .A(n7), .Z(n516));
Q_FDP4EP tlvp_rsm_usr_insert_REG  ( .CK(clk), .CE(n516), .R(n512), .D(n269), .Q(tlvp_rsm_usr_insert));
Q_INV U954 ( .A(tlvp_rsm_usr_insert), .Z(n351));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\tlvp_rsm_ob_wdata.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\tlvp_rsm_ob_wdata.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\tlvp_rsm_ob_wdata.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\tlvp_rsm_ob_wdata.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\pt_ob_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\pt_ob_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\pt_ob_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\pt_ob_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\pt_ob_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\pt_ob_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\tlvp_rsm_usr_ob_rdata.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\tlvp_rsm_usr_ob_rdata.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\tlvp_rsm_usr_ob_rdata.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\tlvp_rsm_usr_ob_rdata.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\tlvp_rsm_usr_ob_rdata.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\tlvp_rsm_usr_ob_rdata.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\tlvp_rsm_usr_ob_rdata_dw0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\tlvp_rsm_usr_ob_rdata_dw0.resv0  (1,0) 1 18 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\tlvp_rsm_usr_ob_rdata_dw0.resv1  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\tlvp_rsm_usr_ob_rdata_dw0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\tlvp_rsm_usr_ob_rdata_dw0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\tlvp_rsm_usr_ob_rdata_dw0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\tlvp_rsm_usr_ob_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\tlvp_rsm_usr_ob_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\tlvp_rsm_usr_ob_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\tlvp_rsm_usr_ob_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\tlvp_rsm_usr_ob_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\tlvp_rsm_usr_ob_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\tlvp_rsm_pt_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\tlvp_rsm_pt_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\tlvp_rsm_pt_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\tlvp_rsm_pt_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\tlvp_rsm_pt_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\tlvp_rsm_pt_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\tlvp_rsm_ob_datain.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\tlvp_rsm_ob_datain.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m39 "\tlvp_rsm_ob_datain.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m40 "\tlvp_rsm_ob_datain.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m41 "\tlvp_rsm_ob_datain.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m42 "\tlvp_rsm_ob_datain.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "42"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "tlvp_rsm_ob_wdata 6 \tlvp_rsm_ob_wdata.tvalid  \tlvp_rsm_ob_wdata.tlast  \tlvp_rsm_ob_wdata.tid  \tlvp_rsm_ob_wdata.tstrb  \tlvp_rsm_ob_wdata.tuser  \tlvp_rsm_ob_wdata.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "pt_ob_tlv 10 \pt_ob_tlv.insert  \pt_ob_tlv.ordern  \pt_ob_tlv.typen  \pt_ob_tlv.sot  \pt_ob_tlv.eot  \pt_ob_tlv.tlast  \pt_ob_tlv.tid  \pt_ob_tlv.tstrb  \pt_ob_tlv.tuser  \pt_ob_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "tlvp_rsm_usr_ob_rdata 10 \tlvp_rsm_usr_ob_rdata.insert  \tlvp_rsm_usr_ob_rdata.ordern  \tlvp_rsm_usr_ob_rdata.typen  \tlvp_rsm_usr_ob_rdata.sot  \tlvp_rsm_usr_ob_rdata.eot  \tlvp_rsm_usr_ob_rdata.tlast  \tlvp_rsm_usr_ob_rdata.tid  \tlvp_rsm_usr_ob_rdata.tstrb  \tlvp_rsm_usr_ob_rdata.tuser  \tlvp_rsm_usr_ob_rdata.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "tlvp_rsm_usr_ob_rdata_dw0 8 \tlvp_rsm_usr_ob_rdata_dw0.tlv_bip2  \tlvp_rsm_usr_ob_rdata_dw0.resv0  \tlvp_rsm_usr_ob_rdata_dw0.tlv_frame_num  \tlvp_rsm_usr_ob_rdata_dw0.resv1  \tlvp_rsm_usr_ob_rdata_dw0.tlv_eng_id  \tlvp_rsm_usr_ob_rdata_dw0.tlv_seq_num  \tlvp_rsm_usr_ob_rdata_dw0.tlv_len  \tlvp_rsm_usr_ob_rdata_dw0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "tlvp_rsm_usr_ob_tlv 10 \tlvp_rsm_usr_ob_tlv.insert  \tlvp_rsm_usr_ob_tlv.ordern  \tlvp_rsm_usr_ob_tlv.typen  \tlvp_rsm_usr_ob_tlv.sot  \tlvp_rsm_usr_ob_tlv.eot  \tlvp_rsm_usr_ob_tlv.tlast  \tlvp_rsm_usr_ob_tlv.tid  \tlvp_rsm_usr_ob_tlv.tstrb  \tlvp_rsm_usr_ob_tlv.tuser  \tlvp_rsm_usr_ob_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "tlvp_rsm_pt_tlv 10 \tlvp_rsm_pt_tlv.insert  \tlvp_rsm_pt_tlv.ordern  \tlvp_rsm_pt_tlv.typen  \tlvp_rsm_pt_tlv.sot  \tlvp_rsm_pt_tlv.eot  \tlvp_rsm_pt_tlv.tlast  \tlvp_rsm_pt_tlv.tid  \tlvp_rsm_pt_tlv.tstrb  \tlvp_rsm_pt_tlv.tuser  \tlvp_rsm_pt_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "tlvp_rsm_ob_datain 10 \tlvp_rsm_ob_datain.insert  \tlvp_rsm_ob_datain.ordern  \tlvp_rsm_ob_datain.typen  \tlvp_rsm_ob_datain.sot  \tlvp_rsm_ob_datain.eot  \tlvp_rsm_ob_datain.tlast  \tlvp_rsm_ob_datain.tid  \tlvp_rsm_ob_datain.tstrb  \tlvp_rsm_ob_datain.tuser  \tlvp_rsm_ob_datain.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "7"
endmodule
