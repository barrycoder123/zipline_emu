architecture module of ixc_frequency_ptm is
  -- quickturn CVASTRPROP MODULE HDLICE IXCOM_FREQUENCY_CELL "1"
  -- quickturn CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE

begin
end module;
