architecture module of ixc_gfifo_bind_512_2 is

begin
end module;
