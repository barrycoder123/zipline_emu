
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_fifo_xcm26 ( empty, full, underflow, overflow, used_slots, free_slots, 
	rdata, clk, rst_n, wen, ren, clear, wdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output empty;
output full;
output underflow;
output overflow;
output [2:0] used_slots;
output [2:0] free_slots;
output [610:0] rdata;
input clk;
input rst_n;
input wen;
input ren;
input clear;
input [610:0] wdata;
wire _zy_simnet_underflow_0_w$;
wire _zy_simnet_overflow_1_w$;
wire \depth_n._zy_simnet_overflow_3_w$ ;
wire \depth_n._zy_simnet_underflow_2_w$ ;
wire [1:0] \depth_n.wptr ;
wire [1:0] \depth_n.rptr ;
supply0 n1235;
ixc_assign _zz_strnp_3 ( _zy_simnet_overflow_1_w$, overflow);
ixc_assign _zz_strnp_2 ( _zy_simnet_underflow_0_w$, underflow);
Q_FDP0 U2 ( .CK(clk), .D(wdata[610]), .Q(n1234), .QN( ));
Q_FDP0 U3 ( .CK(clk), .D(wdata[609]), .Q(n1233), .QN( ));
Q_FDP0 U4 ( .CK(clk), .D(wdata[608]), .Q(n1232), .QN( ));
Q_FDP0 U5 ( .CK(clk), .D(wdata[607]), .Q(n1231), .QN( ));
Q_FDP0 U6 ( .CK(clk), .D(wdata[606]), .Q(n1230), .QN( ));
Q_FDP0 U7 ( .CK(clk), .D(wdata[605]), .Q(n1229), .QN( ));
Q_FDP0 U8 ( .CK(clk), .D(wdata[604]), .Q(n1228), .QN( ));
Q_FDP0 U9 ( .CK(clk), .D(wdata[603]), .Q(n1227), .QN( ));
Q_FDP0 U10 ( .CK(clk), .D(wdata[602]), .Q(n1226), .QN( ));
Q_FDP0 U11 ( .CK(clk), .D(wdata[601]), .Q(n1225), .QN( ));
Q_FDP0 U12 ( .CK(clk), .D(wdata[600]), .Q(n1224), .QN( ));
Q_FDP0 U13 ( .CK(clk), .D(wdata[599]), .Q(n1223), .QN( ));
Q_FDP0 U14 ( .CK(clk), .D(wdata[598]), .Q(n1222), .QN( ));
Q_FDP0 U15 ( .CK(clk), .D(wdata[597]), .Q(n1221), .QN( ));
Q_FDP0 U16 ( .CK(clk), .D(wdata[596]), .Q(n1220), .QN( ));
Q_FDP0 U17 ( .CK(clk), .D(wdata[595]), .Q(n1219), .QN( ));
Q_FDP0 U18 ( .CK(clk), .D(wdata[594]), .Q(n1218), .QN( ));
Q_FDP0 U19 ( .CK(clk), .D(wdata[593]), .Q(n1217), .QN( ));
Q_FDP0 U20 ( .CK(clk), .D(wdata[592]), .Q(n1216), .QN( ));
Q_FDP0 U21 ( .CK(clk), .D(wdata[591]), .Q(n1215), .QN( ));
Q_FDP0 U22 ( .CK(clk), .D(wdata[590]), .Q(n1214), .QN( ));
Q_FDP0 U23 ( .CK(clk), .D(wdata[589]), .Q(n1213), .QN( ));
Q_FDP0 U24 ( .CK(clk), .D(wdata[588]), .Q(n1212), .QN( ));
Q_FDP0 U25 ( .CK(clk), .D(wdata[587]), .Q(n1211), .QN( ));
Q_FDP0 U26 ( .CK(clk), .D(wdata[586]), .Q(n1210), .QN( ));
Q_FDP0 U27 ( .CK(clk), .D(wdata[585]), .Q(n1209), .QN( ));
Q_FDP0 U28 ( .CK(clk), .D(wdata[584]), .Q(n1208), .QN( ));
Q_FDP0 U29 ( .CK(clk), .D(wdata[583]), .Q(n1207), .QN( ));
Q_FDP0 U30 ( .CK(clk), .D(wdata[582]), .Q(n1206), .QN( ));
Q_FDP0 U31 ( .CK(clk), .D(wdata[581]), .Q(n1205), .QN( ));
Q_FDP0 U32 ( .CK(clk), .D(wdata[580]), .Q(n1204), .QN( ));
Q_FDP0 U33 ( .CK(clk), .D(wdata[579]), .Q(n1203), .QN( ));
Q_FDP0 U34 ( .CK(clk), .D(wdata[578]), .Q(n1202), .QN( ));
Q_FDP0 U35 ( .CK(clk), .D(wdata[577]), .Q(n1201), .QN( ));
Q_FDP0 U36 ( .CK(clk), .D(wdata[576]), .Q(n1200), .QN( ));
Q_FDP0 U37 ( .CK(clk), .D(wdata[575]), .Q(n1199), .QN( ));
Q_FDP0 U38 ( .CK(clk), .D(wdata[574]), .Q(n1198), .QN( ));
Q_FDP0 U39 ( .CK(clk), .D(wdata[573]), .Q(n1197), .QN( ));
Q_FDP0 U40 ( .CK(clk), .D(wdata[572]), .Q(n1196), .QN( ));
Q_FDP0 U41 ( .CK(clk), .D(wdata[571]), .Q(n1195), .QN( ));
Q_FDP0 U42 ( .CK(clk), .D(wdata[570]), .Q(n1194), .QN( ));
Q_FDP0 U43 ( .CK(clk), .D(wdata[569]), .Q(n1193), .QN( ));
Q_FDP0 U44 ( .CK(clk), .D(wdata[568]), .Q(n1192), .QN( ));
Q_FDP0 U45 ( .CK(clk), .D(wdata[567]), .Q(n1191), .QN( ));
Q_FDP0 U46 ( .CK(clk), .D(wdata[566]), .Q(n1190), .QN( ));
Q_FDP0 U47 ( .CK(clk), .D(wdata[565]), .Q(n1189), .QN( ));
Q_FDP0 U48 ( .CK(clk), .D(wdata[564]), .Q(n1188), .QN( ));
Q_FDP0 U49 ( .CK(clk), .D(wdata[563]), .Q(n1187), .QN( ));
Q_FDP0 U50 ( .CK(clk), .D(wdata[562]), .Q(n1186), .QN( ));
Q_FDP0 U51 ( .CK(clk), .D(wdata[561]), .Q(n1185), .QN( ));
Q_FDP0 U52 ( .CK(clk), .D(wdata[560]), .Q(n1184), .QN( ));
Q_FDP0 U53 ( .CK(clk), .D(wdata[559]), .Q(n1183), .QN( ));
Q_FDP0 U54 ( .CK(clk), .D(wdata[558]), .Q(n1182), .QN( ));
Q_FDP0 U55 ( .CK(clk), .D(wdata[557]), .Q(n1181), .QN( ));
Q_FDP0 U56 ( .CK(clk), .D(wdata[556]), .Q(n1180), .QN( ));
Q_FDP0 U57 ( .CK(clk), .D(wdata[555]), .Q(n1179), .QN( ));
Q_FDP0 U58 ( .CK(clk), .D(wdata[554]), .Q(n1178), .QN( ));
Q_FDP0 U59 ( .CK(clk), .D(wdata[553]), .Q(n1177), .QN( ));
Q_FDP0 U60 ( .CK(clk), .D(wdata[552]), .Q(n1176), .QN( ));
Q_FDP0 U61 ( .CK(clk), .D(wdata[551]), .Q(n1175), .QN( ));
Q_FDP0 U62 ( .CK(clk), .D(wdata[550]), .Q(n1174), .QN( ));
Q_FDP0 U63 ( .CK(clk), .D(wdata[549]), .Q(n1173), .QN( ));
Q_FDP0 U64 ( .CK(clk), .D(wdata[548]), .Q(n1172), .QN( ));
Q_FDP0 U65 ( .CK(clk), .D(wdata[547]), .Q(n1171), .QN( ));
Q_FDP0 U66 ( .CK(clk), .D(wdata[546]), .Q(n1170), .QN( ));
Q_FDP0 U67 ( .CK(clk), .D(wdata[545]), .Q(n1169), .QN( ));
Q_FDP0 U68 ( .CK(clk), .D(wdata[544]), .Q(n1168), .QN( ));
Q_FDP0 U69 ( .CK(clk), .D(wdata[543]), .Q(n1167), .QN( ));
Q_FDP0 U70 ( .CK(clk), .D(wdata[542]), .Q(n1166), .QN( ));
Q_FDP0 U71 ( .CK(clk), .D(wdata[541]), .Q(n1165), .QN( ));
Q_FDP0 U72 ( .CK(clk), .D(wdata[540]), .Q(n1164), .QN( ));
Q_FDP0 U73 ( .CK(clk), .D(wdata[539]), .Q(n1163), .QN( ));
Q_FDP0 U74 ( .CK(clk), .D(wdata[538]), .Q(n1162), .QN( ));
Q_FDP0 U75 ( .CK(clk), .D(wdata[537]), .Q(n1161), .QN( ));
Q_FDP0 U76 ( .CK(clk), .D(wdata[536]), .Q(n1160), .QN( ));
Q_FDP0 U77 ( .CK(clk), .D(wdata[535]), .Q(n1159), .QN( ));
Q_FDP0 U78 ( .CK(clk), .D(wdata[534]), .Q(n1158), .QN( ));
Q_FDP0 U79 ( .CK(clk), .D(wdata[533]), .Q(n1157), .QN( ));
Q_FDP0 U80 ( .CK(clk), .D(wdata[532]), .Q(n1156), .QN( ));
Q_FDP0 U81 ( .CK(clk), .D(wdata[531]), .Q(n1155), .QN( ));
Q_FDP0 U82 ( .CK(clk), .D(wdata[530]), .Q(n1154), .QN( ));
Q_FDP0 U83 ( .CK(clk), .D(wdata[529]), .Q(n1153), .QN( ));
Q_FDP0 U84 ( .CK(clk), .D(wdata[528]), .Q(n1152), .QN( ));
Q_FDP0 U85 ( .CK(clk), .D(wdata[527]), .Q(n1151), .QN( ));
Q_FDP0 U86 ( .CK(clk), .D(wdata[526]), .Q(n1150), .QN( ));
Q_FDP0 U87 ( .CK(clk), .D(wdata[525]), .Q(n1149), .QN( ));
Q_FDP0 U88 ( .CK(clk), .D(wdata[524]), .Q(n1148), .QN( ));
Q_FDP0 U89 ( .CK(clk), .D(wdata[523]), .Q(n1147), .QN( ));
Q_FDP0 U90 ( .CK(clk), .D(wdata[522]), .Q(n1146), .QN( ));
Q_FDP0 U91 ( .CK(clk), .D(wdata[521]), .Q(n1145), .QN( ));
Q_FDP0 U92 ( .CK(clk), .D(wdata[520]), .Q(n1144), .QN( ));
Q_FDP0 U93 ( .CK(clk), .D(wdata[519]), .Q(n1143), .QN( ));
Q_FDP0 U94 ( .CK(clk), .D(wdata[518]), .Q(n1142), .QN( ));
Q_FDP0 U95 ( .CK(clk), .D(wdata[517]), .Q(n1141), .QN( ));
Q_FDP0 U96 ( .CK(clk), .D(wdata[516]), .Q(n1140), .QN( ));
Q_FDP0 U97 ( .CK(clk), .D(wdata[515]), .Q(n1139), .QN( ));
Q_FDP0 U98 ( .CK(clk), .D(wdata[514]), .Q(n1138), .QN( ));
Q_FDP0 U99 ( .CK(clk), .D(wdata[513]), .Q(n1137), .QN( ));
Q_FDP0 U100 ( .CK(clk), .D(wdata[512]), .Q(n1136), .QN( ));
Q_FDP0 U101 ( .CK(clk), .D(wdata[511]), .Q(n1135), .QN( ));
Q_FDP0 U102 ( .CK(clk), .D(wdata[510]), .Q(n1134), .QN( ));
Q_FDP0 U103 ( .CK(clk), .D(wdata[509]), .Q(n1133), .QN( ));
Q_FDP0 U104 ( .CK(clk), .D(wdata[508]), .Q(n1132), .QN( ));
Q_FDP0 U105 ( .CK(clk), .D(wdata[507]), .Q(n1131), .QN( ));
Q_FDP0 U106 ( .CK(clk), .D(wdata[506]), .Q(n1130), .QN( ));
Q_FDP0 U107 ( .CK(clk), .D(wdata[505]), .Q(n1129), .QN( ));
Q_FDP0 U108 ( .CK(clk), .D(wdata[504]), .Q(n1128), .QN( ));
Q_FDP0 U109 ( .CK(clk), .D(wdata[503]), .Q(n1127), .QN( ));
Q_FDP0 U110 ( .CK(clk), .D(wdata[502]), .Q(n1126), .QN( ));
Q_FDP0 U111 ( .CK(clk), .D(wdata[501]), .Q(n1125), .QN( ));
Q_FDP0 U112 ( .CK(clk), .D(wdata[500]), .Q(n1124), .QN( ));
Q_FDP0 U113 ( .CK(clk), .D(wdata[499]), .Q(n1123), .QN( ));
Q_FDP0 U114 ( .CK(clk), .D(wdata[498]), .Q(n1122), .QN( ));
Q_FDP0 U115 ( .CK(clk), .D(wdata[497]), .Q(n1121), .QN( ));
Q_FDP0 U116 ( .CK(clk), .D(wdata[496]), .Q(n1120), .QN( ));
Q_FDP0 U117 ( .CK(clk), .D(wdata[495]), .Q(n1119), .QN( ));
Q_FDP0 U118 ( .CK(clk), .D(wdata[494]), .Q(n1118), .QN( ));
Q_FDP0 U119 ( .CK(clk), .D(wdata[493]), .Q(n1117), .QN( ));
Q_FDP0 U120 ( .CK(clk), .D(wdata[492]), .Q(n1116), .QN( ));
Q_FDP0 U121 ( .CK(clk), .D(wdata[491]), .Q(n1115), .QN( ));
Q_FDP0 U122 ( .CK(clk), .D(wdata[490]), .Q(n1114), .QN( ));
Q_FDP0 U123 ( .CK(clk), .D(wdata[489]), .Q(n1113), .QN( ));
Q_FDP0 U124 ( .CK(clk), .D(wdata[488]), .Q(n1112), .QN( ));
Q_FDP0 U125 ( .CK(clk), .D(wdata[487]), .Q(n1111), .QN( ));
Q_FDP0 U126 ( .CK(clk), .D(wdata[486]), .Q(n1110), .QN( ));
Q_FDP0 U127 ( .CK(clk), .D(wdata[485]), .Q(n1109), .QN( ));
Q_FDP0 U128 ( .CK(clk), .D(wdata[484]), .Q(n1108), .QN( ));
Q_FDP0 U129 ( .CK(clk), .D(wdata[483]), .Q(n1107), .QN( ));
Q_FDP0 U130 ( .CK(clk), .D(wdata[482]), .Q(n1106), .QN( ));
Q_FDP0 U131 ( .CK(clk), .D(wdata[481]), .Q(n1105), .QN( ));
Q_FDP0 U132 ( .CK(clk), .D(wdata[480]), .Q(n1104), .QN( ));
Q_FDP0 U133 ( .CK(clk), .D(wdata[479]), .Q(n1103), .QN( ));
Q_FDP0 U134 ( .CK(clk), .D(wdata[478]), .Q(n1102), .QN( ));
Q_FDP0 U135 ( .CK(clk), .D(wdata[477]), .Q(n1101), .QN( ));
Q_FDP0 U136 ( .CK(clk), .D(wdata[476]), .Q(n1100), .QN( ));
Q_FDP0 U137 ( .CK(clk), .D(wdata[475]), .Q(n1099), .QN( ));
Q_FDP0 U138 ( .CK(clk), .D(wdata[474]), .Q(n1098), .QN( ));
Q_FDP0 U139 ( .CK(clk), .D(wdata[473]), .Q(n1097), .QN( ));
Q_FDP0 U140 ( .CK(clk), .D(wdata[472]), .Q(n1096), .QN( ));
Q_FDP0 U141 ( .CK(clk), .D(wdata[471]), .Q(n1095), .QN( ));
Q_FDP0 U142 ( .CK(clk), .D(wdata[470]), .Q(n1094), .QN( ));
Q_FDP0 U143 ( .CK(clk), .D(wdata[469]), .Q(n1093), .QN( ));
Q_FDP0 U144 ( .CK(clk), .D(wdata[468]), .Q(n1092), .QN( ));
Q_FDP0 U145 ( .CK(clk), .D(wdata[467]), .Q(n1091), .QN( ));
Q_FDP0 U146 ( .CK(clk), .D(wdata[466]), .Q(n1090), .QN( ));
Q_FDP0 U147 ( .CK(clk), .D(wdata[465]), .Q(n1089), .QN( ));
Q_FDP0 U148 ( .CK(clk), .D(wdata[464]), .Q(n1088), .QN( ));
Q_FDP0 U149 ( .CK(clk), .D(wdata[463]), .Q(n1087), .QN( ));
Q_FDP0 U150 ( .CK(clk), .D(wdata[462]), .Q(n1086), .QN( ));
Q_FDP0 U151 ( .CK(clk), .D(wdata[461]), .Q(n1085), .QN( ));
Q_FDP0 U152 ( .CK(clk), .D(wdata[460]), .Q(n1084), .QN( ));
Q_FDP0 U153 ( .CK(clk), .D(wdata[459]), .Q(n1083), .QN( ));
Q_FDP0 U154 ( .CK(clk), .D(wdata[458]), .Q(n1082), .QN( ));
Q_FDP0 U155 ( .CK(clk), .D(wdata[457]), .Q(n1081), .QN( ));
Q_FDP0 U156 ( .CK(clk), .D(wdata[456]), .Q(n1080), .QN( ));
Q_FDP0 U157 ( .CK(clk), .D(wdata[455]), .Q(n1079), .QN( ));
Q_FDP0 U158 ( .CK(clk), .D(wdata[454]), .Q(n1078), .QN( ));
Q_FDP0 U159 ( .CK(clk), .D(wdata[453]), .Q(n1077), .QN( ));
Q_FDP0 U160 ( .CK(clk), .D(wdata[452]), .Q(n1076), .QN( ));
Q_FDP0 U161 ( .CK(clk), .D(wdata[451]), .Q(n1075), .QN( ));
Q_FDP0 U162 ( .CK(clk), .D(wdata[450]), .Q(n1074), .QN( ));
Q_FDP0 U163 ( .CK(clk), .D(wdata[449]), .Q(n1073), .QN( ));
Q_FDP0 U164 ( .CK(clk), .D(wdata[448]), .Q(n1072), .QN( ));
Q_FDP0 U165 ( .CK(clk), .D(wdata[447]), .Q(n1071), .QN( ));
Q_FDP0 U166 ( .CK(clk), .D(wdata[446]), .Q(n1070), .QN( ));
Q_FDP0 U167 ( .CK(clk), .D(wdata[445]), .Q(n1069), .QN( ));
Q_FDP0 U168 ( .CK(clk), .D(wdata[444]), .Q(n1068), .QN( ));
Q_FDP0 U169 ( .CK(clk), .D(wdata[443]), .Q(n1067), .QN( ));
Q_FDP0 U170 ( .CK(clk), .D(wdata[442]), .Q(n1066), .QN( ));
Q_FDP0 U171 ( .CK(clk), .D(wdata[441]), .Q(n1065), .QN( ));
Q_FDP0 U172 ( .CK(clk), .D(wdata[440]), .Q(n1064), .QN( ));
Q_FDP0 U173 ( .CK(clk), .D(wdata[439]), .Q(n1063), .QN( ));
Q_FDP0 U174 ( .CK(clk), .D(wdata[438]), .Q(n1062), .QN( ));
Q_FDP0 U175 ( .CK(clk), .D(wdata[437]), .Q(n1061), .QN( ));
Q_FDP0 U176 ( .CK(clk), .D(wdata[436]), .Q(n1060), .QN( ));
Q_FDP0 U177 ( .CK(clk), .D(wdata[435]), .Q(n1059), .QN( ));
Q_FDP0 U178 ( .CK(clk), .D(wdata[434]), .Q(n1058), .QN( ));
Q_FDP0 U179 ( .CK(clk), .D(wdata[433]), .Q(n1057), .QN( ));
Q_FDP0 U180 ( .CK(clk), .D(wdata[432]), .Q(n1056), .QN( ));
Q_FDP0 U181 ( .CK(clk), .D(wdata[431]), .Q(n1055), .QN( ));
Q_FDP0 U182 ( .CK(clk), .D(wdata[430]), .Q(n1054), .QN( ));
Q_FDP0 U183 ( .CK(clk), .D(wdata[429]), .Q(n1053), .QN( ));
Q_FDP0 U184 ( .CK(clk), .D(wdata[428]), .Q(n1052), .QN( ));
Q_FDP0 U185 ( .CK(clk), .D(wdata[427]), .Q(n1051), .QN( ));
Q_FDP0 U186 ( .CK(clk), .D(wdata[426]), .Q(n1050), .QN( ));
Q_FDP0 U187 ( .CK(clk), .D(wdata[425]), .Q(n1049), .QN( ));
Q_FDP0 U188 ( .CK(clk), .D(wdata[424]), .Q(n1048), .QN( ));
Q_FDP0 U189 ( .CK(clk), .D(wdata[423]), .Q(n1047), .QN( ));
Q_FDP0 U190 ( .CK(clk), .D(wdata[422]), .Q(n1046), .QN( ));
Q_FDP0 U191 ( .CK(clk), .D(wdata[421]), .Q(n1045), .QN( ));
Q_FDP0 U192 ( .CK(clk), .D(wdata[420]), .Q(n1044), .QN( ));
Q_FDP0 U193 ( .CK(clk), .D(wdata[419]), .Q(n1043), .QN( ));
Q_FDP0 U194 ( .CK(clk), .D(wdata[418]), .Q(n1042), .QN( ));
Q_FDP0 U195 ( .CK(clk), .D(wdata[417]), .Q(n1041), .QN( ));
Q_FDP0 U196 ( .CK(clk), .D(wdata[416]), .Q(n1040), .QN( ));
Q_FDP0 U197 ( .CK(clk), .D(wdata[415]), .Q(n1039), .QN( ));
Q_FDP0 U198 ( .CK(clk), .D(wdata[414]), .Q(n1038), .QN( ));
Q_FDP0 U199 ( .CK(clk), .D(wdata[413]), .Q(n1037), .QN( ));
Q_FDP0 U200 ( .CK(clk), .D(wdata[412]), .Q(n1036), .QN( ));
Q_FDP0 U201 ( .CK(clk), .D(wdata[411]), .Q(n1035), .QN( ));
Q_FDP0 U202 ( .CK(clk), .D(wdata[410]), .Q(n1034), .QN( ));
Q_FDP0 U203 ( .CK(clk), .D(wdata[409]), .Q(n1033), .QN( ));
Q_FDP0 U204 ( .CK(clk), .D(wdata[408]), .Q(n1032), .QN( ));
Q_FDP0 U205 ( .CK(clk), .D(wdata[407]), .Q(n1031), .QN( ));
Q_FDP0 U206 ( .CK(clk), .D(wdata[406]), .Q(n1030), .QN( ));
Q_FDP0 U207 ( .CK(clk), .D(wdata[405]), .Q(n1029), .QN( ));
Q_FDP0 U208 ( .CK(clk), .D(wdata[404]), .Q(n1028), .QN( ));
Q_FDP0 U209 ( .CK(clk), .D(wdata[403]), .Q(n1027), .QN( ));
Q_FDP0 U210 ( .CK(clk), .D(wdata[402]), .Q(n1026), .QN( ));
Q_FDP0 U211 ( .CK(clk), .D(wdata[401]), .Q(n1025), .QN( ));
Q_FDP0 U212 ( .CK(clk), .D(wdata[400]), .Q(n1024), .QN( ));
Q_FDP0 U213 ( .CK(clk), .D(wdata[399]), .Q(n1023), .QN( ));
Q_FDP0 U214 ( .CK(clk), .D(wdata[398]), .Q(n1022), .QN( ));
Q_FDP0 U215 ( .CK(clk), .D(wdata[397]), .Q(n1021), .QN( ));
Q_FDP0 U216 ( .CK(clk), .D(wdata[396]), .Q(n1020), .QN( ));
Q_FDP0 U217 ( .CK(clk), .D(wdata[395]), .Q(n1019), .QN( ));
Q_FDP0 U218 ( .CK(clk), .D(wdata[394]), .Q(n1018), .QN( ));
Q_FDP0 U219 ( .CK(clk), .D(wdata[393]), .Q(n1017), .QN( ));
Q_FDP0 U220 ( .CK(clk), .D(wdata[392]), .Q(n1016), .QN( ));
Q_FDP0 U221 ( .CK(clk), .D(wdata[391]), .Q(n1015), .QN( ));
Q_FDP0 U222 ( .CK(clk), .D(wdata[390]), .Q(n1014), .QN( ));
Q_FDP0 U223 ( .CK(clk), .D(wdata[389]), .Q(n1013), .QN( ));
Q_FDP0 U224 ( .CK(clk), .D(wdata[388]), .Q(n1012), .QN( ));
Q_FDP0 U225 ( .CK(clk), .D(wdata[387]), .Q(n1011), .QN( ));
Q_FDP0 U226 ( .CK(clk), .D(wdata[386]), .Q(n1010), .QN( ));
Q_FDP0 U227 ( .CK(clk), .D(wdata[385]), .Q(n1009), .QN( ));
Q_FDP0 U228 ( .CK(clk), .D(wdata[384]), .Q(n1008), .QN( ));
Q_FDP0 U229 ( .CK(clk), .D(wdata[383]), .Q(n1007), .QN( ));
Q_FDP0 U230 ( .CK(clk), .D(wdata[382]), .Q(n1006), .QN( ));
Q_FDP0 U231 ( .CK(clk), .D(wdata[381]), .Q(n1005), .QN( ));
Q_FDP0 U232 ( .CK(clk), .D(wdata[380]), .Q(n1004), .QN( ));
Q_FDP0 U233 ( .CK(clk), .D(wdata[379]), .Q(n1003), .QN( ));
Q_FDP0 U234 ( .CK(clk), .D(wdata[378]), .Q(n1002), .QN( ));
Q_FDP0 U235 ( .CK(clk), .D(wdata[377]), .Q(n1001), .QN( ));
Q_FDP0 U236 ( .CK(clk), .D(wdata[376]), .Q(n1000), .QN( ));
Q_FDP0 U237 ( .CK(clk), .D(wdata[375]), .Q(n999), .QN( ));
Q_FDP0 U238 ( .CK(clk), .D(wdata[374]), .Q(n998), .QN( ));
Q_FDP0 U239 ( .CK(clk), .D(wdata[373]), .Q(n997), .QN( ));
Q_FDP0 U240 ( .CK(clk), .D(wdata[372]), .Q(n996), .QN( ));
Q_FDP0 U241 ( .CK(clk), .D(wdata[371]), .Q(n995), .QN( ));
Q_FDP0 U242 ( .CK(clk), .D(wdata[370]), .Q(n994), .QN( ));
Q_FDP0 U243 ( .CK(clk), .D(wdata[369]), .Q(n993), .QN( ));
Q_FDP0 U244 ( .CK(clk), .D(wdata[368]), .Q(n992), .QN( ));
Q_FDP0 U245 ( .CK(clk), .D(wdata[367]), .Q(n991), .QN( ));
Q_FDP0 U246 ( .CK(clk), .D(wdata[366]), .Q(n990), .QN( ));
Q_FDP0 U247 ( .CK(clk), .D(wdata[365]), .Q(n989), .QN( ));
Q_FDP0 U248 ( .CK(clk), .D(wdata[364]), .Q(n988), .QN( ));
Q_FDP0 U249 ( .CK(clk), .D(wdata[363]), .Q(n987), .QN( ));
Q_FDP0 U250 ( .CK(clk), .D(wdata[362]), .Q(n986), .QN( ));
Q_FDP0 U251 ( .CK(clk), .D(wdata[361]), .Q(n985), .QN( ));
Q_FDP0 U252 ( .CK(clk), .D(wdata[360]), .Q(n984), .QN( ));
Q_FDP0 U253 ( .CK(clk), .D(wdata[359]), .Q(n983), .QN( ));
Q_FDP0 U254 ( .CK(clk), .D(wdata[358]), .Q(n982), .QN( ));
Q_FDP0 U255 ( .CK(clk), .D(wdata[357]), .Q(n981), .QN( ));
Q_FDP0 U256 ( .CK(clk), .D(wdata[356]), .Q(n980), .QN( ));
Q_FDP0 U257 ( .CK(clk), .D(wdata[355]), .Q(n979), .QN( ));
Q_FDP0 U258 ( .CK(clk), .D(wdata[354]), .Q(n978), .QN( ));
Q_FDP0 U259 ( .CK(clk), .D(wdata[353]), .Q(n977), .QN( ));
Q_FDP0 U260 ( .CK(clk), .D(wdata[352]), .Q(n976), .QN( ));
Q_FDP0 U261 ( .CK(clk), .D(wdata[351]), .Q(n975), .QN( ));
Q_FDP0 U262 ( .CK(clk), .D(wdata[350]), .Q(n974), .QN( ));
Q_FDP0 U263 ( .CK(clk), .D(wdata[349]), .Q(n973), .QN( ));
Q_FDP0 U264 ( .CK(clk), .D(wdata[348]), .Q(n972), .QN( ));
Q_FDP0 U265 ( .CK(clk), .D(wdata[347]), .Q(n971), .QN( ));
Q_FDP0 U266 ( .CK(clk), .D(wdata[346]), .Q(n970), .QN( ));
Q_FDP0 U267 ( .CK(clk), .D(wdata[345]), .Q(n969), .QN( ));
Q_FDP0 U268 ( .CK(clk), .D(wdata[344]), .Q(n968), .QN( ));
Q_FDP0 U269 ( .CK(clk), .D(wdata[343]), .Q(n967), .QN( ));
Q_FDP0 U270 ( .CK(clk), .D(wdata[342]), .Q(n966), .QN( ));
Q_FDP0 U271 ( .CK(clk), .D(wdata[341]), .Q(n965), .QN( ));
Q_FDP0 U272 ( .CK(clk), .D(wdata[340]), .Q(n964), .QN( ));
Q_FDP0 U273 ( .CK(clk), .D(wdata[339]), .Q(n963), .QN( ));
Q_FDP0 U274 ( .CK(clk), .D(wdata[338]), .Q(n962), .QN( ));
Q_FDP0 U275 ( .CK(clk), .D(wdata[337]), .Q(n961), .QN( ));
Q_FDP0 U276 ( .CK(clk), .D(wdata[336]), .Q(n960), .QN( ));
Q_FDP0 U277 ( .CK(clk), .D(wdata[335]), .Q(n959), .QN( ));
Q_FDP0 U278 ( .CK(clk), .D(wdata[334]), .Q(n958), .QN( ));
Q_FDP0 U279 ( .CK(clk), .D(wdata[333]), .Q(n957), .QN( ));
Q_FDP0 U280 ( .CK(clk), .D(wdata[332]), .Q(n956), .QN( ));
Q_FDP0 U281 ( .CK(clk), .D(wdata[331]), .Q(n955), .QN( ));
Q_FDP0 U282 ( .CK(clk), .D(wdata[330]), .Q(n954), .QN( ));
Q_FDP0 U283 ( .CK(clk), .D(wdata[329]), .Q(n953), .QN( ));
Q_FDP0 U284 ( .CK(clk), .D(wdata[328]), .Q(n952), .QN( ));
Q_FDP0 U285 ( .CK(clk), .D(wdata[327]), .Q(n951), .QN( ));
Q_FDP0 U286 ( .CK(clk), .D(wdata[326]), .Q(n950), .QN( ));
Q_FDP0 U287 ( .CK(clk), .D(wdata[325]), .Q(n949), .QN( ));
Q_FDP0 U288 ( .CK(clk), .D(wdata[324]), .Q(n948), .QN( ));
Q_FDP0 U289 ( .CK(clk), .D(wdata[323]), .Q(n947), .QN( ));
Q_FDP0 U290 ( .CK(clk), .D(wdata[322]), .Q(n946), .QN( ));
Q_FDP0 U291 ( .CK(clk), .D(wdata[321]), .Q(n945), .QN( ));
Q_FDP0 U292 ( .CK(clk), .D(wdata[320]), .Q(n944), .QN( ));
Q_FDP0 U293 ( .CK(clk), .D(wdata[319]), .Q(n943), .QN( ));
Q_FDP0 U294 ( .CK(clk), .D(wdata[318]), .Q(n942), .QN( ));
Q_FDP0 U295 ( .CK(clk), .D(wdata[317]), .Q(n941), .QN( ));
Q_FDP0 U296 ( .CK(clk), .D(wdata[316]), .Q(n940), .QN( ));
Q_FDP0 U297 ( .CK(clk), .D(wdata[315]), .Q(n939), .QN( ));
Q_FDP0 U298 ( .CK(clk), .D(wdata[314]), .Q(n938), .QN( ));
Q_FDP0 U299 ( .CK(clk), .D(wdata[313]), .Q(n937), .QN( ));
Q_FDP0 U300 ( .CK(clk), .D(wdata[312]), .Q(n936), .QN( ));
Q_FDP0 U301 ( .CK(clk), .D(wdata[311]), .Q(n935), .QN( ));
Q_FDP0 U302 ( .CK(clk), .D(wdata[310]), .Q(n934), .QN( ));
Q_FDP0 U303 ( .CK(clk), .D(wdata[309]), .Q(n933), .QN( ));
Q_FDP0 U304 ( .CK(clk), .D(wdata[308]), .Q(n932), .QN( ));
Q_FDP0 U305 ( .CK(clk), .D(wdata[307]), .Q(n931), .QN( ));
Q_FDP0 U306 ( .CK(clk), .D(wdata[306]), .Q(n930), .QN( ));
Q_FDP0 U307 ( .CK(clk), .D(wdata[305]), .Q(n929), .QN( ));
Q_FDP0 U308 ( .CK(clk), .D(wdata[304]), .Q(n928), .QN( ));
Q_FDP0 U309 ( .CK(clk), .D(wdata[303]), .Q(n927), .QN( ));
Q_FDP0 U310 ( .CK(clk), .D(wdata[302]), .Q(n926), .QN( ));
Q_FDP0 U311 ( .CK(clk), .D(wdata[301]), .Q(n925), .QN( ));
Q_FDP0 U312 ( .CK(clk), .D(wdata[300]), .Q(n924), .QN( ));
Q_FDP0 U313 ( .CK(clk), .D(wdata[299]), .Q(n923), .QN( ));
Q_FDP0 U314 ( .CK(clk), .D(wdata[298]), .Q(n922), .QN( ));
Q_FDP0 U315 ( .CK(clk), .D(wdata[297]), .Q(n921), .QN( ));
Q_FDP0 U316 ( .CK(clk), .D(wdata[296]), .Q(n920), .QN( ));
Q_FDP0 U317 ( .CK(clk), .D(wdata[295]), .Q(n919), .QN( ));
Q_FDP0 U318 ( .CK(clk), .D(wdata[294]), .Q(n918), .QN( ));
Q_FDP0 U319 ( .CK(clk), .D(wdata[293]), .Q(n917), .QN( ));
Q_FDP0 U320 ( .CK(clk), .D(wdata[292]), .Q(n916), .QN( ));
Q_FDP0 U321 ( .CK(clk), .D(wdata[291]), .Q(n915), .QN( ));
Q_FDP0 U322 ( .CK(clk), .D(wdata[290]), .Q(n914), .QN( ));
Q_FDP0 U323 ( .CK(clk), .D(wdata[289]), .Q(n913), .QN( ));
Q_FDP0 U324 ( .CK(clk), .D(wdata[288]), .Q(n912), .QN( ));
Q_FDP0 U325 ( .CK(clk), .D(wdata[287]), .Q(n911), .QN( ));
Q_FDP0 U326 ( .CK(clk), .D(wdata[286]), .Q(n910), .QN( ));
Q_FDP0 U327 ( .CK(clk), .D(wdata[285]), .Q(n909), .QN( ));
Q_FDP0 U328 ( .CK(clk), .D(wdata[284]), .Q(n908), .QN( ));
Q_FDP0 U329 ( .CK(clk), .D(wdata[283]), .Q(n907), .QN( ));
Q_FDP0 U330 ( .CK(clk), .D(wdata[282]), .Q(n906), .QN( ));
Q_FDP0 U331 ( .CK(clk), .D(wdata[281]), .Q(n905), .QN( ));
Q_FDP0 U332 ( .CK(clk), .D(wdata[280]), .Q(n904), .QN( ));
Q_FDP0 U333 ( .CK(clk), .D(wdata[279]), .Q(n903), .QN( ));
Q_FDP0 U334 ( .CK(clk), .D(wdata[278]), .Q(n902), .QN( ));
Q_FDP0 U335 ( .CK(clk), .D(wdata[277]), .Q(n901), .QN( ));
Q_FDP0 U336 ( .CK(clk), .D(wdata[276]), .Q(n900), .QN( ));
Q_FDP0 U337 ( .CK(clk), .D(wdata[275]), .Q(n899), .QN( ));
Q_FDP0 U338 ( .CK(clk), .D(wdata[274]), .Q(n898), .QN( ));
Q_FDP0 U339 ( .CK(clk), .D(wdata[273]), .Q(n897), .QN( ));
Q_FDP0 U340 ( .CK(clk), .D(wdata[272]), .Q(n896), .QN( ));
Q_FDP0 U341 ( .CK(clk), .D(wdata[271]), .Q(n895), .QN( ));
Q_FDP0 U342 ( .CK(clk), .D(wdata[270]), .Q(n894), .QN( ));
Q_FDP0 U343 ( .CK(clk), .D(wdata[269]), .Q(n893), .QN( ));
Q_FDP0 U344 ( .CK(clk), .D(wdata[268]), .Q(n892), .QN( ));
Q_FDP0 U345 ( .CK(clk), .D(wdata[267]), .Q(n891), .QN( ));
Q_FDP0 U346 ( .CK(clk), .D(wdata[266]), .Q(n890), .QN( ));
Q_FDP0 U347 ( .CK(clk), .D(wdata[265]), .Q(n889), .QN( ));
Q_FDP0 U348 ( .CK(clk), .D(wdata[264]), .Q(n888), .QN( ));
Q_FDP0 U349 ( .CK(clk), .D(wdata[263]), .Q(n887), .QN( ));
Q_FDP0 U350 ( .CK(clk), .D(wdata[262]), .Q(n886), .QN( ));
Q_FDP0 U351 ( .CK(clk), .D(wdata[261]), .Q(n885), .QN( ));
Q_FDP0 U352 ( .CK(clk), .D(wdata[260]), .Q(n884), .QN( ));
Q_FDP0 U353 ( .CK(clk), .D(wdata[259]), .Q(n883), .QN( ));
Q_FDP0 U354 ( .CK(clk), .D(wdata[258]), .Q(n882), .QN( ));
Q_FDP0 U355 ( .CK(clk), .D(wdata[257]), .Q(n881), .QN( ));
Q_FDP0 U356 ( .CK(clk), .D(wdata[256]), .Q(n880), .QN( ));
Q_FDP0 U357 ( .CK(clk), .D(wdata[255]), .Q(n879), .QN( ));
Q_FDP0 U358 ( .CK(clk), .D(wdata[254]), .Q(n878), .QN( ));
Q_FDP0 U359 ( .CK(clk), .D(wdata[253]), .Q(n877), .QN( ));
Q_FDP0 U360 ( .CK(clk), .D(wdata[252]), .Q(n876), .QN( ));
Q_FDP0 U361 ( .CK(clk), .D(wdata[251]), .Q(n875), .QN( ));
Q_FDP0 U362 ( .CK(clk), .D(wdata[250]), .Q(n874), .QN( ));
Q_FDP0 U363 ( .CK(clk), .D(wdata[249]), .Q(n873), .QN( ));
Q_FDP0 U364 ( .CK(clk), .D(wdata[248]), .Q(n872), .QN( ));
Q_FDP0 U365 ( .CK(clk), .D(wdata[247]), .Q(n871), .QN( ));
Q_FDP0 U366 ( .CK(clk), .D(wdata[246]), .Q(n870), .QN( ));
Q_FDP0 U367 ( .CK(clk), .D(wdata[245]), .Q(n869), .QN( ));
Q_FDP0 U368 ( .CK(clk), .D(wdata[244]), .Q(n868), .QN( ));
Q_FDP0 U369 ( .CK(clk), .D(wdata[243]), .Q(n867), .QN( ));
Q_FDP0 U370 ( .CK(clk), .D(wdata[242]), .Q(n866), .QN( ));
Q_FDP0 U371 ( .CK(clk), .D(wdata[241]), .Q(n865), .QN( ));
Q_FDP0 U372 ( .CK(clk), .D(wdata[240]), .Q(n864), .QN( ));
Q_FDP0 U373 ( .CK(clk), .D(wdata[239]), .Q(n863), .QN( ));
Q_FDP0 U374 ( .CK(clk), .D(wdata[238]), .Q(n862), .QN( ));
Q_FDP0 U375 ( .CK(clk), .D(wdata[237]), .Q(n861), .QN( ));
Q_FDP0 U376 ( .CK(clk), .D(wdata[236]), .Q(n860), .QN( ));
Q_FDP0 U377 ( .CK(clk), .D(wdata[235]), .Q(n859), .QN( ));
Q_FDP0 U378 ( .CK(clk), .D(wdata[234]), .Q(n858), .QN( ));
Q_FDP0 U379 ( .CK(clk), .D(wdata[233]), .Q(n857), .QN( ));
Q_FDP0 U380 ( .CK(clk), .D(wdata[232]), .Q(n856), .QN( ));
Q_FDP0 U381 ( .CK(clk), .D(wdata[231]), .Q(n855), .QN( ));
Q_FDP0 U382 ( .CK(clk), .D(wdata[230]), .Q(n854), .QN( ));
Q_FDP0 U383 ( .CK(clk), .D(wdata[229]), .Q(n853), .QN( ));
Q_FDP0 U384 ( .CK(clk), .D(wdata[228]), .Q(n852), .QN( ));
Q_FDP0 U385 ( .CK(clk), .D(wdata[227]), .Q(n851), .QN( ));
Q_FDP0 U386 ( .CK(clk), .D(wdata[226]), .Q(n850), .QN( ));
Q_FDP0 U387 ( .CK(clk), .D(wdata[225]), .Q(n849), .QN( ));
Q_FDP0 U388 ( .CK(clk), .D(wdata[224]), .Q(n848), .QN( ));
Q_FDP0 U389 ( .CK(clk), .D(wdata[223]), .Q(n847), .QN( ));
Q_FDP0 U390 ( .CK(clk), .D(wdata[222]), .Q(n846), .QN( ));
Q_FDP0 U391 ( .CK(clk), .D(wdata[221]), .Q(n845), .QN( ));
Q_FDP0 U392 ( .CK(clk), .D(wdata[220]), .Q(n844), .QN( ));
Q_FDP0 U393 ( .CK(clk), .D(wdata[219]), .Q(n843), .QN( ));
Q_FDP0 U394 ( .CK(clk), .D(wdata[218]), .Q(n842), .QN( ));
Q_FDP0 U395 ( .CK(clk), .D(wdata[217]), .Q(n841), .QN( ));
Q_FDP0 U396 ( .CK(clk), .D(wdata[216]), .Q(n840), .QN( ));
Q_FDP0 U397 ( .CK(clk), .D(wdata[215]), .Q(n839), .QN( ));
Q_FDP0 U398 ( .CK(clk), .D(wdata[214]), .Q(n838), .QN( ));
Q_FDP0 U399 ( .CK(clk), .D(wdata[213]), .Q(n837), .QN( ));
Q_FDP0 U400 ( .CK(clk), .D(wdata[212]), .Q(n836), .QN( ));
Q_FDP0 U401 ( .CK(clk), .D(wdata[211]), .Q(n835), .QN( ));
Q_FDP0 U402 ( .CK(clk), .D(wdata[210]), .Q(n834), .QN( ));
Q_FDP0 U403 ( .CK(clk), .D(wdata[209]), .Q(n833), .QN( ));
Q_FDP0 U404 ( .CK(clk), .D(wdata[208]), .Q(n832), .QN( ));
Q_FDP0 U405 ( .CK(clk), .D(wdata[207]), .Q(n831), .QN( ));
Q_FDP0 U406 ( .CK(clk), .D(wdata[206]), .Q(n830), .QN( ));
Q_FDP0 U407 ( .CK(clk), .D(wdata[205]), .Q(n829), .QN( ));
Q_FDP0 U408 ( .CK(clk), .D(wdata[204]), .Q(n828), .QN( ));
Q_FDP0 U409 ( .CK(clk), .D(wdata[203]), .Q(n827), .QN( ));
Q_FDP0 U410 ( .CK(clk), .D(wdata[202]), .Q(n826), .QN( ));
Q_FDP0 U411 ( .CK(clk), .D(wdata[201]), .Q(n825), .QN( ));
Q_FDP0 U412 ( .CK(clk), .D(wdata[200]), .Q(n824), .QN( ));
Q_FDP0 U413 ( .CK(clk), .D(wdata[199]), .Q(n823), .QN( ));
Q_FDP0 U414 ( .CK(clk), .D(wdata[198]), .Q(n822), .QN( ));
Q_FDP0 U415 ( .CK(clk), .D(wdata[197]), .Q(n821), .QN( ));
Q_FDP0 U416 ( .CK(clk), .D(wdata[196]), .Q(n820), .QN( ));
Q_FDP0 U417 ( .CK(clk), .D(wdata[195]), .Q(n819), .QN( ));
Q_FDP0 U418 ( .CK(clk), .D(wdata[194]), .Q(n818), .QN( ));
Q_FDP0 U419 ( .CK(clk), .D(wdata[193]), .Q(n817), .QN( ));
Q_FDP0 U420 ( .CK(clk), .D(wdata[192]), .Q(n816), .QN( ));
Q_FDP0 U421 ( .CK(clk), .D(wdata[191]), .Q(n815), .QN( ));
Q_FDP0 U422 ( .CK(clk), .D(wdata[190]), .Q(n814), .QN( ));
Q_FDP0 U423 ( .CK(clk), .D(wdata[189]), .Q(n813), .QN( ));
Q_FDP0 U424 ( .CK(clk), .D(wdata[188]), .Q(n812), .QN( ));
Q_FDP0 U425 ( .CK(clk), .D(wdata[187]), .Q(n811), .QN( ));
Q_FDP0 U426 ( .CK(clk), .D(wdata[186]), .Q(n810), .QN( ));
Q_FDP0 U427 ( .CK(clk), .D(wdata[185]), .Q(n809), .QN( ));
Q_FDP0 U428 ( .CK(clk), .D(wdata[184]), .Q(n808), .QN( ));
Q_FDP0 U429 ( .CK(clk), .D(wdata[183]), .Q(n807), .QN( ));
Q_FDP0 U430 ( .CK(clk), .D(wdata[182]), .Q(n806), .QN( ));
Q_FDP0 U431 ( .CK(clk), .D(wdata[181]), .Q(n805), .QN( ));
Q_FDP0 U432 ( .CK(clk), .D(wdata[180]), .Q(n804), .QN( ));
Q_FDP0 U433 ( .CK(clk), .D(wdata[179]), .Q(n803), .QN( ));
Q_FDP0 U434 ( .CK(clk), .D(wdata[178]), .Q(n802), .QN( ));
Q_FDP0 U435 ( .CK(clk), .D(wdata[177]), .Q(n801), .QN( ));
Q_FDP0 U436 ( .CK(clk), .D(wdata[176]), .Q(n800), .QN( ));
Q_FDP0 U437 ( .CK(clk), .D(wdata[175]), .Q(n799), .QN( ));
Q_FDP0 U438 ( .CK(clk), .D(wdata[174]), .Q(n798), .QN( ));
Q_FDP0 U439 ( .CK(clk), .D(wdata[173]), .Q(n797), .QN( ));
Q_FDP0 U440 ( .CK(clk), .D(wdata[172]), .Q(n796), .QN( ));
Q_FDP0 U441 ( .CK(clk), .D(wdata[171]), .Q(n795), .QN( ));
Q_FDP0 U442 ( .CK(clk), .D(wdata[170]), .Q(n794), .QN( ));
Q_FDP0 U443 ( .CK(clk), .D(wdata[169]), .Q(n793), .QN( ));
Q_FDP0 U444 ( .CK(clk), .D(wdata[168]), .Q(n792), .QN( ));
Q_FDP0 U445 ( .CK(clk), .D(wdata[167]), .Q(n791), .QN( ));
Q_FDP0 U446 ( .CK(clk), .D(wdata[166]), .Q(n790), .QN( ));
Q_FDP0 U447 ( .CK(clk), .D(wdata[165]), .Q(n789), .QN( ));
Q_FDP0 U448 ( .CK(clk), .D(wdata[164]), .Q(n788), .QN( ));
Q_FDP0 U449 ( .CK(clk), .D(wdata[163]), .Q(n787), .QN( ));
Q_FDP0 U450 ( .CK(clk), .D(wdata[162]), .Q(n786), .QN( ));
Q_FDP0 U451 ( .CK(clk), .D(wdata[161]), .Q(n785), .QN( ));
Q_FDP0 U452 ( .CK(clk), .D(wdata[160]), .Q(n784), .QN( ));
Q_FDP0 U453 ( .CK(clk), .D(wdata[159]), .Q(n783), .QN( ));
Q_FDP0 U454 ( .CK(clk), .D(wdata[158]), .Q(n782), .QN( ));
Q_FDP0 U455 ( .CK(clk), .D(wdata[157]), .Q(n781), .QN( ));
Q_FDP0 U456 ( .CK(clk), .D(wdata[156]), .Q(n780), .QN( ));
Q_FDP0 U457 ( .CK(clk), .D(wdata[155]), .Q(n779), .QN( ));
Q_FDP0 U458 ( .CK(clk), .D(wdata[154]), .Q(n778), .QN( ));
Q_FDP0 U459 ( .CK(clk), .D(wdata[153]), .Q(n777), .QN( ));
Q_FDP0 U460 ( .CK(clk), .D(wdata[152]), .Q(n776), .QN( ));
Q_FDP0 U461 ( .CK(clk), .D(wdata[151]), .Q(n775), .QN( ));
Q_FDP0 U462 ( .CK(clk), .D(wdata[150]), .Q(n774), .QN( ));
Q_FDP0 U463 ( .CK(clk), .D(wdata[149]), .Q(n773), .QN( ));
Q_FDP0 U464 ( .CK(clk), .D(wdata[148]), .Q(n772), .QN( ));
Q_FDP0 U465 ( .CK(clk), .D(wdata[147]), .Q(n771), .QN( ));
Q_FDP0 U466 ( .CK(clk), .D(wdata[146]), .Q(n770), .QN( ));
Q_FDP0 U467 ( .CK(clk), .D(wdata[145]), .Q(n769), .QN( ));
Q_FDP0 U468 ( .CK(clk), .D(wdata[144]), .Q(n768), .QN( ));
Q_FDP0 U469 ( .CK(clk), .D(wdata[143]), .Q(n767), .QN( ));
Q_FDP0 U470 ( .CK(clk), .D(wdata[142]), .Q(n766), .QN( ));
Q_FDP0 U471 ( .CK(clk), .D(wdata[141]), .Q(n765), .QN( ));
Q_FDP0 U472 ( .CK(clk), .D(wdata[140]), .Q(n764), .QN( ));
Q_FDP0 U473 ( .CK(clk), .D(wdata[139]), .Q(n763), .QN( ));
Q_FDP0 U474 ( .CK(clk), .D(wdata[138]), .Q(n762), .QN( ));
Q_FDP0 U475 ( .CK(clk), .D(wdata[137]), .Q(n761), .QN( ));
Q_FDP0 U476 ( .CK(clk), .D(wdata[136]), .Q(n760), .QN( ));
Q_FDP0 U477 ( .CK(clk), .D(wdata[135]), .Q(n759), .QN( ));
Q_FDP0 U478 ( .CK(clk), .D(wdata[134]), .Q(n758), .QN( ));
Q_FDP0 U479 ( .CK(clk), .D(wdata[133]), .Q(n757), .QN( ));
Q_FDP0 U480 ( .CK(clk), .D(wdata[132]), .Q(n756), .QN( ));
Q_FDP0 U481 ( .CK(clk), .D(wdata[131]), .Q(n755), .QN( ));
Q_FDP0 U482 ( .CK(clk), .D(wdata[130]), .Q(n754), .QN( ));
Q_FDP0 U483 ( .CK(clk), .D(wdata[129]), .Q(n753), .QN( ));
Q_FDP0 U484 ( .CK(clk), .D(wdata[128]), .Q(n752), .QN( ));
Q_FDP0 U485 ( .CK(clk), .D(wdata[127]), .Q(n751), .QN( ));
Q_FDP0 U486 ( .CK(clk), .D(wdata[126]), .Q(n750), .QN( ));
Q_FDP0 U487 ( .CK(clk), .D(wdata[125]), .Q(n749), .QN( ));
Q_FDP0 U488 ( .CK(clk), .D(wdata[124]), .Q(n748), .QN( ));
Q_FDP0 U489 ( .CK(clk), .D(wdata[123]), .Q(n747), .QN( ));
Q_FDP0 U490 ( .CK(clk), .D(wdata[122]), .Q(n746), .QN( ));
Q_FDP0 U491 ( .CK(clk), .D(wdata[121]), .Q(n745), .QN( ));
Q_FDP0 U492 ( .CK(clk), .D(wdata[120]), .Q(n744), .QN( ));
Q_FDP0 U493 ( .CK(clk), .D(wdata[119]), .Q(n743), .QN( ));
Q_FDP0 U494 ( .CK(clk), .D(wdata[118]), .Q(n742), .QN( ));
Q_FDP0 U495 ( .CK(clk), .D(wdata[117]), .Q(n741), .QN( ));
Q_FDP0 U496 ( .CK(clk), .D(wdata[116]), .Q(n740), .QN( ));
Q_FDP0 U497 ( .CK(clk), .D(wdata[115]), .Q(n739), .QN( ));
Q_FDP0 U498 ( .CK(clk), .D(wdata[114]), .Q(n738), .QN( ));
Q_FDP0 U499 ( .CK(clk), .D(wdata[113]), .Q(n737), .QN( ));
Q_FDP0 U500 ( .CK(clk), .D(wdata[112]), .Q(n736), .QN( ));
Q_FDP0 U501 ( .CK(clk), .D(wdata[111]), .Q(n735), .QN( ));
Q_FDP0 U502 ( .CK(clk), .D(wdata[110]), .Q(n734), .QN( ));
Q_FDP0 U503 ( .CK(clk), .D(wdata[109]), .Q(n733), .QN( ));
Q_FDP0 U504 ( .CK(clk), .D(wdata[108]), .Q(n732), .QN( ));
Q_FDP0 U505 ( .CK(clk), .D(wdata[107]), .Q(n731), .QN( ));
Q_FDP0 U506 ( .CK(clk), .D(wdata[106]), .Q(n730), .QN( ));
Q_FDP0 U507 ( .CK(clk), .D(wdata[105]), .Q(n729), .QN( ));
Q_FDP0 U508 ( .CK(clk), .D(wdata[104]), .Q(n728), .QN( ));
Q_FDP0 U509 ( .CK(clk), .D(wdata[103]), .Q(n727), .QN( ));
Q_FDP0 U510 ( .CK(clk), .D(wdata[102]), .Q(n726), .QN( ));
Q_FDP0 U511 ( .CK(clk), .D(wdata[101]), .Q(n725), .QN( ));
Q_FDP0 U512 ( .CK(clk), .D(wdata[100]), .Q(n724), .QN( ));
Q_FDP0 U513 ( .CK(clk), .D(wdata[99]), .Q(n723), .QN( ));
Q_FDP0 U514 ( .CK(clk), .D(wdata[98]), .Q(n722), .QN( ));
Q_FDP0 U515 ( .CK(clk), .D(wdata[97]), .Q(n721), .QN( ));
Q_FDP0 U516 ( .CK(clk), .D(wdata[96]), .Q(n720), .QN( ));
Q_FDP0 U517 ( .CK(clk), .D(wdata[95]), .Q(n719), .QN( ));
Q_FDP0 U518 ( .CK(clk), .D(wdata[94]), .Q(n718), .QN( ));
Q_FDP0 U519 ( .CK(clk), .D(wdata[93]), .Q(n717), .QN( ));
Q_FDP0 U520 ( .CK(clk), .D(wdata[92]), .Q(n716), .QN( ));
Q_FDP0 U521 ( .CK(clk), .D(wdata[91]), .Q(n715), .QN( ));
Q_FDP0 U522 ( .CK(clk), .D(wdata[90]), .Q(n714), .QN( ));
Q_FDP0 U523 ( .CK(clk), .D(wdata[89]), .Q(n713), .QN( ));
Q_FDP0 U524 ( .CK(clk), .D(wdata[88]), .Q(n712), .QN( ));
Q_FDP0 U525 ( .CK(clk), .D(wdata[87]), .Q(n711), .QN( ));
Q_FDP0 U526 ( .CK(clk), .D(wdata[86]), .Q(n710), .QN( ));
Q_FDP0 U527 ( .CK(clk), .D(wdata[85]), .Q(n709), .QN( ));
Q_FDP0 U528 ( .CK(clk), .D(wdata[84]), .Q(n708), .QN( ));
Q_FDP0 U529 ( .CK(clk), .D(wdata[83]), .Q(n707), .QN( ));
Q_FDP0 U530 ( .CK(clk), .D(wdata[82]), .Q(n706), .QN( ));
Q_FDP0 U531 ( .CK(clk), .D(wdata[81]), .Q(n705), .QN( ));
Q_FDP0 U532 ( .CK(clk), .D(wdata[80]), .Q(n704), .QN( ));
Q_FDP0 U533 ( .CK(clk), .D(wdata[79]), .Q(n703), .QN( ));
Q_FDP0 U534 ( .CK(clk), .D(wdata[78]), .Q(n702), .QN( ));
Q_FDP0 U535 ( .CK(clk), .D(wdata[77]), .Q(n701), .QN( ));
Q_FDP0 U536 ( .CK(clk), .D(wdata[76]), .Q(n700), .QN( ));
Q_FDP0 U537 ( .CK(clk), .D(wdata[75]), .Q(n699), .QN( ));
Q_FDP0 U538 ( .CK(clk), .D(wdata[74]), .Q(n698), .QN( ));
Q_FDP0 U539 ( .CK(clk), .D(wdata[73]), .Q(n697), .QN( ));
Q_FDP0 U540 ( .CK(clk), .D(wdata[72]), .Q(n696), .QN( ));
Q_FDP0 U541 ( .CK(clk), .D(wdata[71]), .Q(n695), .QN( ));
Q_FDP0 U542 ( .CK(clk), .D(wdata[70]), .Q(n694), .QN( ));
Q_FDP0 U543 ( .CK(clk), .D(wdata[69]), .Q(n693), .QN( ));
Q_FDP0 U544 ( .CK(clk), .D(wdata[68]), .Q(n692), .QN( ));
Q_FDP0 U545 ( .CK(clk), .D(wdata[67]), .Q(n691), .QN( ));
Q_FDP0 U546 ( .CK(clk), .D(wdata[66]), .Q(n690), .QN( ));
Q_FDP0 U547 ( .CK(clk), .D(wdata[65]), .Q(n689), .QN( ));
Q_FDP0 U548 ( .CK(clk), .D(wdata[64]), .Q(n688), .QN( ));
Q_FDP0 U549 ( .CK(clk), .D(wdata[63]), .Q(n687), .QN( ));
Q_FDP0 U550 ( .CK(clk), .D(wdata[62]), .Q(n686), .QN( ));
Q_FDP0 U551 ( .CK(clk), .D(wdata[61]), .Q(n685), .QN( ));
Q_FDP0 U552 ( .CK(clk), .D(wdata[60]), .Q(n684), .QN( ));
Q_FDP0 U553 ( .CK(clk), .D(wdata[59]), .Q(n683), .QN( ));
Q_FDP0 U554 ( .CK(clk), .D(wdata[58]), .Q(n682), .QN( ));
Q_FDP0 U555 ( .CK(clk), .D(wdata[57]), .Q(n681), .QN( ));
Q_FDP0 U556 ( .CK(clk), .D(wdata[56]), .Q(n680), .QN( ));
Q_FDP0 U557 ( .CK(clk), .D(wdata[55]), .Q(n679), .QN( ));
Q_FDP0 U558 ( .CK(clk), .D(wdata[54]), .Q(n678), .QN( ));
Q_FDP0 U559 ( .CK(clk), .D(wdata[53]), .Q(n677), .QN( ));
Q_FDP0 U560 ( .CK(clk), .D(wdata[52]), .Q(n676), .QN( ));
Q_FDP0 U561 ( .CK(clk), .D(wdata[51]), .Q(n675), .QN( ));
Q_FDP0 U562 ( .CK(clk), .D(wdata[50]), .Q(n674), .QN( ));
Q_FDP0 U563 ( .CK(clk), .D(wdata[49]), .Q(n673), .QN( ));
Q_FDP0 U564 ( .CK(clk), .D(wdata[48]), .Q(n672), .QN( ));
Q_FDP0 U565 ( .CK(clk), .D(wdata[47]), .Q(n671), .QN( ));
Q_FDP0 U566 ( .CK(clk), .D(wdata[46]), .Q(n670), .QN( ));
Q_FDP0 U567 ( .CK(clk), .D(wdata[45]), .Q(n669), .QN( ));
Q_FDP0 U568 ( .CK(clk), .D(wdata[44]), .Q(n668), .QN( ));
Q_FDP0 U569 ( .CK(clk), .D(wdata[43]), .Q(n667), .QN( ));
Q_FDP0 U570 ( .CK(clk), .D(wdata[42]), .Q(n666), .QN( ));
Q_FDP0 U571 ( .CK(clk), .D(wdata[41]), .Q(n665), .QN( ));
Q_FDP0 U572 ( .CK(clk), .D(wdata[40]), .Q(n664), .QN( ));
Q_FDP0 U573 ( .CK(clk), .D(wdata[39]), .Q(n663), .QN( ));
Q_FDP0 U574 ( .CK(clk), .D(wdata[38]), .Q(n662), .QN( ));
Q_FDP0 U575 ( .CK(clk), .D(wdata[37]), .Q(n661), .QN( ));
Q_FDP0 U576 ( .CK(clk), .D(wdata[36]), .Q(n660), .QN( ));
Q_FDP0 U577 ( .CK(clk), .D(wdata[35]), .Q(n659), .QN( ));
Q_FDP0 U578 ( .CK(clk), .D(wdata[34]), .Q(n658), .QN( ));
Q_FDP0 U579 ( .CK(clk), .D(wdata[33]), .Q(n657), .QN( ));
Q_FDP0 U580 ( .CK(clk), .D(wdata[32]), .Q(n656), .QN( ));
Q_FDP0 U581 ( .CK(clk), .D(wdata[31]), .Q(n655), .QN( ));
Q_FDP0 U582 ( .CK(clk), .D(wdata[30]), .Q(n654), .QN( ));
Q_FDP0 U583 ( .CK(clk), .D(wdata[29]), .Q(n653), .QN( ));
Q_FDP0 U584 ( .CK(clk), .D(wdata[28]), .Q(n652), .QN( ));
Q_FDP0 U585 ( .CK(clk), .D(wdata[27]), .Q(n651), .QN( ));
Q_FDP0 U586 ( .CK(clk), .D(wdata[26]), .Q(n650), .QN( ));
Q_FDP0 U587 ( .CK(clk), .D(wdata[25]), .Q(n649), .QN( ));
Q_FDP0 U588 ( .CK(clk), .D(wdata[24]), .Q(n648), .QN( ));
Q_FDP0 U589 ( .CK(clk), .D(wdata[23]), .Q(n647), .QN( ));
Q_FDP0 U590 ( .CK(clk), .D(wdata[22]), .Q(n646), .QN( ));
Q_FDP0 U591 ( .CK(clk), .D(wdata[21]), .Q(n645), .QN( ));
Q_FDP0 U592 ( .CK(clk), .D(wdata[20]), .Q(n644), .QN( ));
Q_FDP0 U593 ( .CK(clk), .D(wdata[19]), .Q(n643), .QN( ));
Q_FDP0 U594 ( .CK(clk), .D(wdata[18]), .Q(n642), .QN( ));
Q_FDP0 U595 ( .CK(clk), .D(wdata[17]), .Q(n641), .QN( ));
Q_FDP0 U596 ( .CK(clk), .D(wdata[16]), .Q(n640), .QN( ));
Q_FDP0 U597 ( .CK(clk), .D(wdata[15]), .Q(n639), .QN( ));
Q_FDP0 U598 ( .CK(clk), .D(wdata[14]), .Q(n638), .QN( ));
Q_FDP0 U599 ( .CK(clk), .D(wdata[13]), .Q(n637), .QN( ));
Q_FDP0 U600 ( .CK(clk), .D(wdata[12]), .Q(n636), .QN( ));
Q_FDP0 U601 ( .CK(clk), .D(wdata[11]), .Q(n635), .QN( ));
Q_FDP0 U602 ( .CK(clk), .D(wdata[10]), .Q(n634), .QN( ));
Q_FDP0 U603 ( .CK(clk), .D(wdata[9]), .Q(n633), .QN( ));
Q_FDP0 U604 ( .CK(clk), .D(wdata[8]), .Q(n632), .QN( ));
Q_FDP0 U605 ( .CK(clk), .D(wdata[7]), .Q(n631), .QN( ));
Q_FDP0 U606 ( .CK(clk), .D(wdata[6]), .Q(n630), .QN( ));
Q_FDP0 U607 ( .CK(clk), .D(wdata[5]), .Q(n629), .QN( ));
Q_FDP0 U608 ( .CK(clk), .D(wdata[4]), .Q(n628), .QN( ));
Q_FDP0 U609 ( .CK(clk), .D(wdata[3]), .Q(n627), .QN( ));
Q_FDP0 U610 ( .CK(clk), .D(wdata[2]), .Q(n626), .QN( ));
Q_FDP0 U611 ( .CK(clk), .D(wdata[1]), .Q(n625), .QN( ));
Q_FDP0 U612 ( .CK(clk), .D(wdata[0]), .Q(n624), .QN( ));
Q_FDP0 U613 ( .CK(clk), .D(\depth_n.wptr [1]), .Q(n623), .QN( ));
Q_FDP0 U614 ( .CK(clk), .D(\depth_n.wptr [0]), .Q(n622), .QN( ));
Q_AN02 U615 ( .A0(n617), .A1(n620), .Z(n621));
Q_XOR2 U616 ( .A0(n616), .A1(n619), .Z(n620));
// pragma CVAINTPROP NET n616 _2_state_ 1
// pragma CVAINTPROP INSTANCE U616 NOBREAKS 1
Q_FDP0B U617 ( .D(n616), .QTFCLK( ), .Q(n619));
Q_FDP0 U618 ( .CK(clk), .D(n3), .Q(n617), .QN( ));
Q_FDP0 U619 ( .CK(clk), .D(n618), .Q(n616), .QN(n618));
Q_INV U620 ( .A(empty), .Z(n615));
Q_AN02 U621 ( .A0(n615), .A1(n4), .Z(rdata[610]));
Q_AN02 U622 ( .A0(n615), .A1(n5), .Z(rdata[609]));
Q_AN02 U623 ( .A0(n615), .A1(n6), .Z(rdata[608]));
Q_AN02 U624 ( .A0(n615), .A1(n7), .Z(rdata[607]));
Q_AN02 U625 ( .A0(n615), .A1(n8), .Z(rdata[606]));
Q_AN02 U626 ( .A0(n615), .A1(n9), .Z(rdata[605]));
Q_AN02 U627 ( .A0(n615), .A1(n10), .Z(rdata[604]));
Q_AN02 U628 ( .A0(n615), .A1(n11), .Z(rdata[603]));
Q_AN02 U629 ( .A0(n615), .A1(n12), .Z(rdata[602]));
Q_AN02 U630 ( .A0(n615), .A1(n13), .Z(rdata[601]));
Q_AN02 U631 ( .A0(n615), .A1(n14), .Z(rdata[600]));
Q_AN02 U632 ( .A0(n615), .A1(n15), .Z(rdata[599]));
Q_AN02 U633 ( .A0(n615), .A1(n16), .Z(rdata[598]));
Q_AN02 U634 ( .A0(n615), .A1(n17), .Z(rdata[597]));
Q_AN02 U635 ( .A0(n615), .A1(n18), .Z(rdata[596]));
Q_AN02 U636 ( .A0(n615), .A1(n19), .Z(rdata[595]));
Q_AN02 U637 ( .A0(n615), .A1(n20), .Z(rdata[594]));
Q_AN02 U638 ( .A0(n615), .A1(n21), .Z(rdata[593]));
Q_AN02 U639 ( .A0(n615), .A1(n22), .Z(rdata[592]));
Q_AN02 U640 ( .A0(n615), .A1(n23), .Z(rdata[591]));
Q_AN02 U641 ( .A0(n615), .A1(n24), .Z(rdata[590]));
Q_AN02 U642 ( .A0(n615), .A1(n25), .Z(rdata[589]));
Q_AN02 U643 ( .A0(n615), .A1(n26), .Z(rdata[588]));
Q_AN02 U644 ( .A0(n615), .A1(n27), .Z(rdata[587]));
Q_AN02 U645 ( .A0(n615), .A1(n28), .Z(rdata[586]));
Q_AN02 U646 ( .A0(n615), .A1(n29), .Z(rdata[585]));
Q_AN02 U647 ( .A0(n615), .A1(n30), .Z(rdata[584]));
Q_AN02 U648 ( .A0(n615), .A1(n31), .Z(rdata[583]));
Q_AN02 U649 ( .A0(n615), .A1(n32), .Z(rdata[582]));
Q_AN02 U650 ( .A0(n615), .A1(n33), .Z(rdata[581]));
Q_AN02 U651 ( .A0(n615), .A1(n34), .Z(rdata[580]));
Q_AN02 U652 ( .A0(n615), .A1(n35), .Z(rdata[579]));
Q_AN02 U653 ( .A0(n615), .A1(n36), .Z(rdata[578]));
Q_AN02 U654 ( .A0(n615), .A1(n37), .Z(rdata[577]));
Q_AN02 U655 ( .A0(n615), .A1(n38), .Z(rdata[576]));
Q_AN02 U656 ( .A0(n615), .A1(n39), .Z(rdata[575]));
Q_AN02 U657 ( .A0(n615), .A1(n40), .Z(rdata[574]));
Q_AN02 U658 ( .A0(n615), .A1(n41), .Z(rdata[573]));
Q_AN02 U659 ( .A0(n615), .A1(n42), .Z(rdata[572]));
Q_AN02 U660 ( .A0(n615), .A1(n43), .Z(rdata[571]));
Q_AN02 U661 ( .A0(n615), .A1(n44), .Z(rdata[570]));
Q_AN02 U662 ( .A0(n615), .A1(n45), .Z(rdata[569]));
Q_AN02 U663 ( .A0(n615), .A1(n46), .Z(rdata[568]));
Q_AN02 U664 ( .A0(n615), .A1(n47), .Z(rdata[567]));
Q_AN02 U665 ( .A0(n615), .A1(n48), .Z(rdata[566]));
Q_AN02 U666 ( .A0(n615), .A1(n49), .Z(rdata[565]));
Q_AN02 U667 ( .A0(n615), .A1(n50), .Z(rdata[564]));
Q_AN02 U668 ( .A0(n615), .A1(n51), .Z(rdata[563]));
Q_AN02 U669 ( .A0(n615), .A1(n52), .Z(rdata[562]));
Q_AN02 U670 ( .A0(n615), .A1(n53), .Z(rdata[561]));
Q_AN02 U671 ( .A0(n615), .A1(n54), .Z(rdata[560]));
Q_AN02 U672 ( .A0(n615), .A1(n55), .Z(rdata[559]));
Q_AN02 U673 ( .A0(n615), .A1(n56), .Z(rdata[558]));
Q_AN02 U674 ( .A0(n615), .A1(n57), .Z(rdata[557]));
Q_AN02 U675 ( .A0(n615), .A1(n58), .Z(rdata[556]));
Q_AN02 U676 ( .A0(n615), .A1(n59), .Z(rdata[555]));
Q_AN02 U677 ( .A0(n615), .A1(n60), .Z(rdata[554]));
Q_AN02 U678 ( .A0(n615), .A1(n61), .Z(rdata[553]));
Q_AN02 U679 ( .A0(n615), .A1(n62), .Z(rdata[552]));
Q_AN02 U680 ( .A0(n615), .A1(n63), .Z(rdata[551]));
Q_AN02 U681 ( .A0(n615), .A1(n64), .Z(rdata[550]));
Q_AN02 U682 ( .A0(n615), .A1(n65), .Z(rdata[549]));
Q_AN02 U683 ( .A0(n615), .A1(n66), .Z(rdata[548]));
Q_AN02 U684 ( .A0(n615), .A1(n67), .Z(rdata[547]));
Q_AN02 U685 ( .A0(n615), .A1(n68), .Z(rdata[546]));
Q_AN02 U686 ( .A0(n615), .A1(n69), .Z(rdata[545]));
Q_AN02 U687 ( .A0(n615), .A1(n70), .Z(rdata[544]));
Q_AN02 U688 ( .A0(n615), .A1(n71), .Z(rdata[543]));
Q_AN02 U689 ( .A0(n615), .A1(n72), .Z(rdata[542]));
Q_AN02 U690 ( .A0(n615), .A1(n73), .Z(rdata[541]));
Q_AN02 U691 ( .A0(n615), .A1(n74), .Z(rdata[540]));
Q_AN02 U692 ( .A0(n615), .A1(n75), .Z(rdata[539]));
Q_AN02 U693 ( .A0(n615), .A1(n76), .Z(rdata[538]));
Q_AN02 U694 ( .A0(n615), .A1(n77), .Z(rdata[537]));
Q_AN02 U695 ( .A0(n615), .A1(n78), .Z(rdata[536]));
Q_AN02 U696 ( .A0(n615), .A1(n79), .Z(rdata[535]));
Q_AN02 U697 ( .A0(n615), .A1(n80), .Z(rdata[534]));
Q_AN02 U698 ( .A0(n615), .A1(n81), .Z(rdata[533]));
Q_AN02 U699 ( .A0(n615), .A1(n82), .Z(rdata[532]));
Q_AN02 U700 ( .A0(n615), .A1(n83), .Z(rdata[531]));
Q_AN02 U701 ( .A0(n615), .A1(n84), .Z(rdata[530]));
Q_AN02 U702 ( .A0(n615), .A1(n85), .Z(rdata[529]));
Q_AN02 U703 ( .A0(n615), .A1(n86), .Z(rdata[528]));
Q_AN02 U704 ( .A0(n615), .A1(n87), .Z(rdata[527]));
Q_AN02 U705 ( .A0(n615), .A1(n88), .Z(rdata[526]));
Q_AN02 U706 ( .A0(n615), .A1(n89), .Z(rdata[525]));
Q_AN02 U707 ( .A0(n615), .A1(n90), .Z(rdata[524]));
Q_AN02 U708 ( .A0(n615), .A1(n91), .Z(rdata[523]));
Q_AN02 U709 ( .A0(n615), .A1(n92), .Z(rdata[522]));
Q_AN02 U710 ( .A0(n615), .A1(n93), .Z(rdata[521]));
Q_AN02 U711 ( .A0(n615), .A1(n94), .Z(rdata[520]));
Q_AN02 U712 ( .A0(n615), .A1(n95), .Z(rdata[519]));
Q_AN02 U713 ( .A0(n615), .A1(n96), .Z(rdata[518]));
Q_AN02 U714 ( .A0(n615), .A1(n97), .Z(rdata[517]));
Q_AN02 U715 ( .A0(n615), .A1(n98), .Z(rdata[516]));
Q_AN02 U716 ( .A0(n615), .A1(n99), .Z(rdata[515]));
Q_AN02 U717 ( .A0(n615), .A1(n100), .Z(rdata[514]));
Q_AN02 U718 ( .A0(n615), .A1(n101), .Z(rdata[513]));
Q_AN02 U719 ( .A0(n615), .A1(n102), .Z(rdata[512]));
Q_AN02 U720 ( .A0(n615), .A1(n103), .Z(rdata[511]));
Q_AN02 U721 ( .A0(n615), .A1(n104), .Z(rdata[510]));
Q_AN02 U722 ( .A0(n615), .A1(n105), .Z(rdata[509]));
Q_AN02 U723 ( .A0(n615), .A1(n106), .Z(rdata[508]));
Q_AN02 U724 ( .A0(n615), .A1(n107), .Z(rdata[507]));
Q_AN02 U725 ( .A0(n615), .A1(n108), .Z(rdata[506]));
Q_AN02 U726 ( .A0(n615), .A1(n109), .Z(rdata[505]));
Q_AN02 U727 ( .A0(n615), .A1(n110), .Z(rdata[504]));
Q_AN02 U728 ( .A0(n615), .A1(n111), .Z(rdata[503]));
Q_AN02 U729 ( .A0(n615), .A1(n112), .Z(rdata[502]));
Q_AN02 U730 ( .A0(n615), .A1(n113), .Z(rdata[501]));
Q_AN02 U731 ( .A0(n615), .A1(n114), .Z(rdata[500]));
Q_AN02 U732 ( .A0(n615), .A1(n115), .Z(rdata[499]));
Q_AN02 U733 ( .A0(n615), .A1(n116), .Z(rdata[498]));
Q_AN02 U734 ( .A0(n615), .A1(n117), .Z(rdata[497]));
Q_AN02 U735 ( .A0(n615), .A1(n118), .Z(rdata[496]));
Q_AN02 U736 ( .A0(n615), .A1(n119), .Z(rdata[495]));
Q_AN02 U737 ( .A0(n615), .A1(n120), .Z(rdata[494]));
Q_AN02 U738 ( .A0(n615), .A1(n121), .Z(rdata[493]));
Q_AN02 U739 ( .A0(n615), .A1(n122), .Z(rdata[492]));
Q_AN02 U740 ( .A0(n615), .A1(n123), .Z(rdata[491]));
Q_AN02 U741 ( .A0(n615), .A1(n124), .Z(rdata[490]));
Q_AN02 U742 ( .A0(n615), .A1(n125), .Z(rdata[489]));
Q_AN02 U743 ( .A0(n615), .A1(n126), .Z(rdata[488]));
Q_AN02 U744 ( .A0(n615), .A1(n127), .Z(rdata[487]));
Q_AN02 U745 ( .A0(n615), .A1(n128), .Z(rdata[486]));
Q_AN02 U746 ( .A0(n615), .A1(n129), .Z(rdata[485]));
Q_AN02 U747 ( .A0(n615), .A1(n130), .Z(rdata[484]));
Q_AN02 U748 ( .A0(n615), .A1(n131), .Z(rdata[483]));
Q_AN02 U749 ( .A0(n615), .A1(n132), .Z(rdata[482]));
Q_AN02 U750 ( .A0(n615), .A1(n133), .Z(rdata[481]));
Q_AN02 U751 ( .A0(n615), .A1(n134), .Z(rdata[480]));
Q_AN02 U752 ( .A0(n615), .A1(n135), .Z(rdata[479]));
Q_AN02 U753 ( .A0(n615), .A1(n136), .Z(rdata[478]));
Q_AN02 U754 ( .A0(n615), .A1(n137), .Z(rdata[477]));
Q_AN02 U755 ( .A0(n615), .A1(n138), .Z(rdata[476]));
Q_AN02 U756 ( .A0(n615), .A1(n139), .Z(rdata[475]));
Q_AN02 U757 ( .A0(n615), .A1(n140), .Z(rdata[474]));
Q_AN02 U758 ( .A0(n615), .A1(n141), .Z(rdata[473]));
Q_AN02 U759 ( .A0(n615), .A1(n142), .Z(rdata[472]));
Q_AN02 U760 ( .A0(n615), .A1(n143), .Z(rdata[471]));
Q_AN02 U761 ( .A0(n615), .A1(n144), .Z(rdata[470]));
Q_AN02 U762 ( .A0(n615), .A1(n145), .Z(rdata[469]));
Q_AN02 U763 ( .A0(n615), .A1(n146), .Z(rdata[468]));
Q_AN02 U764 ( .A0(n615), .A1(n147), .Z(rdata[467]));
Q_AN02 U765 ( .A0(n615), .A1(n148), .Z(rdata[466]));
Q_AN02 U766 ( .A0(n615), .A1(n149), .Z(rdata[465]));
Q_AN02 U767 ( .A0(n615), .A1(n150), .Z(rdata[464]));
Q_AN02 U768 ( .A0(n615), .A1(n151), .Z(rdata[463]));
Q_AN02 U769 ( .A0(n615), .A1(n152), .Z(rdata[462]));
Q_AN02 U770 ( .A0(n615), .A1(n153), .Z(rdata[461]));
Q_AN02 U771 ( .A0(n615), .A1(n154), .Z(rdata[460]));
Q_AN02 U772 ( .A0(n615), .A1(n155), .Z(rdata[459]));
Q_AN02 U773 ( .A0(n615), .A1(n156), .Z(rdata[458]));
Q_AN02 U774 ( .A0(n615), .A1(n157), .Z(rdata[457]));
Q_AN02 U775 ( .A0(n615), .A1(n158), .Z(rdata[456]));
Q_AN02 U776 ( .A0(n615), .A1(n159), .Z(rdata[455]));
Q_AN02 U777 ( .A0(n615), .A1(n160), .Z(rdata[454]));
Q_AN02 U778 ( .A0(n615), .A1(n161), .Z(rdata[453]));
Q_AN02 U779 ( .A0(n615), .A1(n162), .Z(rdata[452]));
Q_AN02 U780 ( .A0(n615), .A1(n163), .Z(rdata[451]));
Q_AN02 U781 ( .A0(n615), .A1(n164), .Z(rdata[450]));
Q_AN02 U782 ( .A0(n615), .A1(n165), .Z(rdata[449]));
Q_AN02 U783 ( .A0(n615), .A1(n166), .Z(rdata[448]));
Q_AN02 U784 ( .A0(n615), .A1(n167), .Z(rdata[447]));
Q_AN02 U785 ( .A0(n615), .A1(n168), .Z(rdata[446]));
Q_AN02 U786 ( .A0(n615), .A1(n169), .Z(rdata[445]));
Q_AN02 U787 ( .A0(n615), .A1(n170), .Z(rdata[444]));
Q_AN02 U788 ( .A0(n615), .A1(n171), .Z(rdata[443]));
Q_AN02 U789 ( .A0(n615), .A1(n172), .Z(rdata[442]));
Q_AN02 U790 ( .A0(n615), .A1(n173), .Z(rdata[441]));
Q_AN02 U791 ( .A0(n615), .A1(n174), .Z(rdata[440]));
Q_AN02 U792 ( .A0(n615), .A1(n175), .Z(rdata[439]));
Q_AN02 U793 ( .A0(n615), .A1(n176), .Z(rdata[438]));
Q_AN02 U794 ( .A0(n615), .A1(n177), .Z(rdata[437]));
Q_AN02 U795 ( .A0(n615), .A1(n178), .Z(rdata[436]));
Q_AN02 U796 ( .A0(n615), .A1(n179), .Z(rdata[435]));
Q_AN02 U797 ( .A0(n615), .A1(n180), .Z(rdata[434]));
Q_AN02 U798 ( .A0(n615), .A1(n181), .Z(rdata[433]));
Q_AN02 U799 ( .A0(n615), .A1(n182), .Z(rdata[432]));
Q_AN02 U800 ( .A0(n615), .A1(n183), .Z(rdata[431]));
Q_AN02 U801 ( .A0(n615), .A1(n184), .Z(rdata[430]));
Q_AN02 U802 ( .A0(n615), .A1(n185), .Z(rdata[429]));
Q_AN02 U803 ( .A0(n615), .A1(n186), .Z(rdata[428]));
Q_AN02 U804 ( .A0(n615), .A1(n187), .Z(rdata[427]));
Q_AN02 U805 ( .A0(n615), .A1(n188), .Z(rdata[426]));
Q_AN02 U806 ( .A0(n615), .A1(n189), .Z(rdata[425]));
Q_AN02 U807 ( .A0(n615), .A1(n190), .Z(rdata[424]));
Q_AN02 U808 ( .A0(n615), .A1(n191), .Z(rdata[423]));
Q_AN02 U809 ( .A0(n615), .A1(n192), .Z(rdata[422]));
Q_AN02 U810 ( .A0(n615), .A1(n193), .Z(rdata[421]));
Q_AN02 U811 ( .A0(n615), .A1(n194), .Z(rdata[420]));
Q_AN02 U812 ( .A0(n615), .A1(n195), .Z(rdata[419]));
Q_AN02 U813 ( .A0(n615), .A1(n196), .Z(rdata[418]));
Q_AN02 U814 ( .A0(n615), .A1(n197), .Z(rdata[417]));
Q_AN02 U815 ( .A0(n615), .A1(n198), .Z(rdata[416]));
Q_AN02 U816 ( .A0(n615), .A1(n199), .Z(rdata[415]));
Q_AN02 U817 ( .A0(n615), .A1(n200), .Z(rdata[414]));
Q_AN02 U818 ( .A0(n615), .A1(n201), .Z(rdata[413]));
Q_AN02 U819 ( .A0(n615), .A1(n202), .Z(rdata[412]));
Q_AN02 U820 ( .A0(n615), .A1(n203), .Z(rdata[411]));
Q_AN02 U821 ( .A0(n615), .A1(n204), .Z(rdata[410]));
Q_AN02 U822 ( .A0(n615), .A1(n205), .Z(rdata[409]));
Q_AN02 U823 ( .A0(n615), .A1(n206), .Z(rdata[408]));
Q_AN02 U824 ( .A0(n615), .A1(n207), .Z(rdata[407]));
Q_AN02 U825 ( .A0(n615), .A1(n208), .Z(rdata[406]));
Q_AN02 U826 ( .A0(n615), .A1(n209), .Z(rdata[405]));
Q_AN02 U827 ( .A0(n615), .A1(n210), .Z(rdata[404]));
Q_AN02 U828 ( .A0(n615), .A1(n211), .Z(rdata[403]));
Q_AN02 U829 ( .A0(n615), .A1(n212), .Z(rdata[402]));
Q_AN02 U830 ( .A0(n615), .A1(n213), .Z(rdata[401]));
Q_AN02 U831 ( .A0(n615), .A1(n214), .Z(rdata[400]));
Q_AN02 U832 ( .A0(n615), .A1(n215), .Z(rdata[399]));
Q_AN02 U833 ( .A0(n615), .A1(n216), .Z(rdata[398]));
Q_AN02 U834 ( .A0(n615), .A1(n217), .Z(rdata[397]));
Q_AN02 U835 ( .A0(n615), .A1(n218), .Z(rdata[396]));
Q_AN02 U836 ( .A0(n615), .A1(n219), .Z(rdata[395]));
Q_AN02 U837 ( .A0(n615), .A1(n220), .Z(rdata[394]));
Q_AN02 U838 ( .A0(n615), .A1(n221), .Z(rdata[393]));
Q_AN02 U839 ( .A0(n615), .A1(n222), .Z(rdata[392]));
Q_AN02 U840 ( .A0(n615), .A1(n223), .Z(rdata[391]));
Q_AN02 U841 ( .A0(n615), .A1(n224), .Z(rdata[390]));
Q_AN02 U842 ( .A0(n615), .A1(n225), .Z(rdata[389]));
Q_AN02 U843 ( .A0(n615), .A1(n226), .Z(rdata[388]));
Q_AN02 U844 ( .A0(n615), .A1(n227), .Z(rdata[387]));
Q_AN02 U845 ( .A0(n615), .A1(n228), .Z(rdata[386]));
Q_AN02 U846 ( .A0(n615), .A1(n229), .Z(rdata[385]));
Q_AN02 U847 ( .A0(n615), .A1(n230), .Z(rdata[384]));
Q_AN02 U848 ( .A0(n615), .A1(n231), .Z(rdata[383]));
Q_AN02 U849 ( .A0(n615), .A1(n232), .Z(rdata[382]));
Q_AN02 U850 ( .A0(n615), .A1(n233), .Z(rdata[381]));
Q_AN02 U851 ( .A0(n615), .A1(n234), .Z(rdata[380]));
Q_AN02 U852 ( .A0(n615), .A1(n235), .Z(rdata[379]));
Q_AN02 U853 ( .A0(n615), .A1(n236), .Z(rdata[378]));
Q_AN02 U854 ( .A0(n615), .A1(n237), .Z(rdata[377]));
Q_AN02 U855 ( .A0(n615), .A1(n238), .Z(rdata[376]));
Q_AN02 U856 ( .A0(n615), .A1(n239), .Z(rdata[375]));
Q_AN02 U857 ( .A0(n615), .A1(n240), .Z(rdata[374]));
Q_AN02 U858 ( .A0(n615), .A1(n241), .Z(rdata[373]));
Q_AN02 U859 ( .A0(n615), .A1(n242), .Z(rdata[372]));
Q_AN02 U860 ( .A0(n615), .A1(n243), .Z(rdata[371]));
Q_AN02 U861 ( .A0(n615), .A1(n244), .Z(rdata[370]));
Q_AN02 U862 ( .A0(n615), .A1(n245), .Z(rdata[369]));
Q_AN02 U863 ( .A0(n615), .A1(n246), .Z(rdata[368]));
Q_AN02 U864 ( .A0(n615), .A1(n247), .Z(rdata[367]));
Q_AN02 U865 ( .A0(n615), .A1(n248), .Z(rdata[366]));
Q_AN02 U866 ( .A0(n615), .A1(n249), .Z(rdata[365]));
Q_AN02 U867 ( .A0(n615), .A1(n250), .Z(rdata[364]));
Q_AN02 U868 ( .A0(n615), .A1(n251), .Z(rdata[363]));
Q_AN02 U869 ( .A0(n615), .A1(n252), .Z(rdata[362]));
Q_AN02 U870 ( .A0(n615), .A1(n253), .Z(rdata[361]));
Q_AN02 U871 ( .A0(n615), .A1(n254), .Z(rdata[360]));
Q_AN02 U872 ( .A0(n615), .A1(n255), .Z(rdata[359]));
Q_AN02 U873 ( .A0(n615), .A1(n256), .Z(rdata[358]));
Q_AN02 U874 ( .A0(n615), .A1(n257), .Z(rdata[357]));
Q_AN02 U875 ( .A0(n615), .A1(n258), .Z(rdata[356]));
Q_AN02 U876 ( .A0(n615), .A1(n259), .Z(rdata[355]));
Q_AN02 U877 ( .A0(n615), .A1(n260), .Z(rdata[354]));
Q_AN02 U878 ( .A0(n615), .A1(n261), .Z(rdata[353]));
Q_AN02 U879 ( .A0(n615), .A1(n262), .Z(rdata[352]));
Q_AN02 U880 ( .A0(n615), .A1(n263), .Z(rdata[351]));
Q_AN02 U881 ( .A0(n615), .A1(n264), .Z(rdata[350]));
Q_AN02 U882 ( .A0(n615), .A1(n265), .Z(rdata[349]));
Q_AN02 U883 ( .A0(n615), .A1(n266), .Z(rdata[348]));
Q_AN02 U884 ( .A0(n615), .A1(n267), .Z(rdata[347]));
Q_AN02 U885 ( .A0(n615), .A1(n268), .Z(rdata[346]));
Q_AN02 U886 ( .A0(n615), .A1(n269), .Z(rdata[345]));
Q_AN02 U887 ( .A0(n615), .A1(n270), .Z(rdata[344]));
Q_AN02 U888 ( .A0(n615), .A1(n271), .Z(rdata[343]));
Q_AN02 U889 ( .A0(n615), .A1(n272), .Z(rdata[342]));
Q_AN02 U890 ( .A0(n615), .A1(n273), .Z(rdata[341]));
Q_AN02 U891 ( .A0(n615), .A1(n274), .Z(rdata[340]));
Q_AN02 U892 ( .A0(n615), .A1(n275), .Z(rdata[339]));
Q_AN02 U893 ( .A0(n615), .A1(n276), .Z(rdata[338]));
Q_AN02 U894 ( .A0(n615), .A1(n277), .Z(rdata[337]));
Q_AN02 U895 ( .A0(n615), .A1(n278), .Z(rdata[336]));
Q_AN02 U896 ( .A0(n615), .A1(n279), .Z(rdata[335]));
Q_AN02 U897 ( .A0(n615), .A1(n280), .Z(rdata[334]));
Q_AN02 U898 ( .A0(n615), .A1(n281), .Z(rdata[333]));
Q_AN02 U899 ( .A0(n615), .A1(n282), .Z(rdata[332]));
Q_AN02 U900 ( .A0(n615), .A1(n283), .Z(rdata[331]));
Q_AN02 U901 ( .A0(n615), .A1(n284), .Z(rdata[330]));
Q_AN02 U902 ( .A0(n615), .A1(n285), .Z(rdata[329]));
Q_AN02 U903 ( .A0(n615), .A1(n286), .Z(rdata[328]));
Q_AN02 U904 ( .A0(n615), .A1(n287), .Z(rdata[327]));
Q_AN02 U905 ( .A0(n615), .A1(n288), .Z(rdata[326]));
Q_AN02 U906 ( .A0(n615), .A1(n289), .Z(rdata[325]));
Q_AN02 U907 ( .A0(n615), .A1(n290), .Z(rdata[324]));
Q_AN02 U908 ( .A0(n615), .A1(n291), .Z(rdata[323]));
Q_AN02 U909 ( .A0(n615), .A1(n292), .Z(rdata[322]));
Q_AN02 U910 ( .A0(n615), .A1(n293), .Z(rdata[321]));
Q_AN02 U911 ( .A0(n615), .A1(n294), .Z(rdata[320]));
Q_AN02 U912 ( .A0(n615), .A1(n295), .Z(rdata[319]));
Q_AN02 U913 ( .A0(n615), .A1(n296), .Z(rdata[318]));
Q_AN02 U914 ( .A0(n615), .A1(n297), .Z(rdata[317]));
Q_AN02 U915 ( .A0(n615), .A1(n298), .Z(rdata[316]));
Q_AN02 U916 ( .A0(n615), .A1(n299), .Z(rdata[315]));
Q_AN02 U917 ( .A0(n615), .A1(n300), .Z(rdata[314]));
Q_AN02 U918 ( .A0(n615), .A1(n301), .Z(rdata[313]));
Q_AN02 U919 ( .A0(n615), .A1(n302), .Z(rdata[312]));
Q_AN02 U920 ( .A0(n615), .A1(n303), .Z(rdata[311]));
Q_AN02 U921 ( .A0(n615), .A1(n304), .Z(rdata[310]));
Q_AN02 U922 ( .A0(n615), .A1(n305), .Z(rdata[309]));
Q_AN02 U923 ( .A0(n615), .A1(n306), .Z(rdata[308]));
Q_AN02 U924 ( .A0(n615), .A1(n307), .Z(rdata[307]));
Q_AN02 U925 ( .A0(n615), .A1(n308), .Z(rdata[306]));
Q_AN02 U926 ( .A0(n615), .A1(n309), .Z(rdata[305]));
Q_AN02 U927 ( .A0(n615), .A1(n310), .Z(rdata[304]));
Q_AN02 U928 ( .A0(n615), .A1(n311), .Z(rdata[303]));
Q_AN02 U929 ( .A0(n615), .A1(n312), .Z(rdata[302]));
Q_AN02 U930 ( .A0(n615), .A1(n313), .Z(rdata[301]));
Q_AN02 U931 ( .A0(n615), .A1(n314), .Z(rdata[300]));
Q_AN02 U932 ( .A0(n615), .A1(n315), .Z(rdata[299]));
Q_AN02 U933 ( .A0(n615), .A1(n316), .Z(rdata[298]));
Q_AN02 U934 ( .A0(n615), .A1(n317), .Z(rdata[297]));
Q_AN02 U935 ( .A0(n615), .A1(n318), .Z(rdata[296]));
Q_AN02 U936 ( .A0(n615), .A1(n319), .Z(rdata[295]));
Q_AN02 U937 ( .A0(n615), .A1(n320), .Z(rdata[294]));
Q_AN02 U938 ( .A0(n615), .A1(n321), .Z(rdata[293]));
Q_AN02 U939 ( .A0(n615), .A1(n322), .Z(rdata[292]));
Q_AN02 U940 ( .A0(n615), .A1(n323), .Z(rdata[291]));
Q_AN02 U941 ( .A0(n615), .A1(n324), .Z(rdata[290]));
Q_AN02 U942 ( .A0(n615), .A1(n325), .Z(rdata[289]));
Q_AN02 U943 ( .A0(n615), .A1(n326), .Z(rdata[288]));
Q_AN02 U944 ( .A0(n615), .A1(n327), .Z(rdata[287]));
Q_AN02 U945 ( .A0(n615), .A1(n328), .Z(rdata[286]));
Q_AN02 U946 ( .A0(n615), .A1(n329), .Z(rdata[285]));
Q_AN02 U947 ( .A0(n615), .A1(n330), .Z(rdata[284]));
Q_AN02 U948 ( .A0(n615), .A1(n331), .Z(rdata[283]));
Q_AN02 U949 ( .A0(n615), .A1(n332), .Z(rdata[282]));
Q_AN02 U950 ( .A0(n615), .A1(n333), .Z(rdata[281]));
Q_AN02 U951 ( .A0(n615), .A1(n334), .Z(rdata[280]));
Q_AN02 U952 ( .A0(n615), .A1(n335), .Z(rdata[279]));
Q_AN02 U953 ( .A0(n615), .A1(n336), .Z(rdata[278]));
Q_AN02 U954 ( .A0(n615), .A1(n337), .Z(rdata[277]));
Q_AN02 U955 ( .A0(n615), .A1(n338), .Z(rdata[276]));
Q_AN02 U956 ( .A0(n615), .A1(n339), .Z(rdata[275]));
Q_AN02 U957 ( .A0(n615), .A1(n340), .Z(rdata[274]));
Q_AN02 U958 ( .A0(n615), .A1(n341), .Z(rdata[273]));
Q_AN02 U959 ( .A0(n615), .A1(n342), .Z(rdata[272]));
Q_AN02 U960 ( .A0(n615), .A1(n343), .Z(rdata[271]));
Q_AN02 U961 ( .A0(n615), .A1(n344), .Z(rdata[270]));
Q_AN02 U962 ( .A0(n615), .A1(n345), .Z(rdata[269]));
Q_AN02 U963 ( .A0(n615), .A1(n346), .Z(rdata[268]));
Q_AN02 U964 ( .A0(n615), .A1(n347), .Z(rdata[267]));
Q_AN02 U965 ( .A0(n615), .A1(n348), .Z(rdata[266]));
Q_AN02 U966 ( .A0(n615), .A1(n349), .Z(rdata[265]));
Q_AN02 U967 ( .A0(n615), .A1(n350), .Z(rdata[264]));
Q_AN02 U968 ( .A0(n615), .A1(n351), .Z(rdata[263]));
Q_AN02 U969 ( .A0(n615), .A1(n352), .Z(rdata[262]));
Q_AN02 U970 ( .A0(n615), .A1(n353), .Z(rdata[261]));
Q_AN02 U971 ( .A0(n615), .A1(n354), .Z(rdata[260]));
Q_AN02 U972 ( .A0(n615), .A1(n355), .Z(rdata[259]));
Q_AN02 U973 ( .A0(n615), .A1(n356), .Z(rdata[258]));
Q_AN02 U974 ( .A0(n615), .A1(n357), .Z(rdata[257]));
Q_AN02 U975 ( .A0(n615), .A1(n358), .Z(rdata[256]));
Q_AN02 U976 ( .A0(n615), .A1(n359), .Z(rdata[255]));
Q_AN02 U977 ( .A0(n615), .A1(n360), .Z(rdata[254]));
Q_AN02 U978 ( .A0(n615), .A1(n361), .Z(rdata[253]));
Q_AN02 U979 ( .A0(n615), .A1(n362), .Z(rdata[252]));
Q_AN02 U980 ( .A0(n615), .A1(n363), .Z(rdata[251]));
Q_AN02 U981 ( .A0(n615), .A1(n364), .Z(rdata[250]));
Q_AN02 U982 ( .A0(n615), .A1(n365), .Z(rdata[249]));
Q_AN02 U983 ( .A0(n615), .A1(n366), .Z(rdata[248]));
Q_AN02 U984 ( .A0(n615), .A1(n367), .Z(rdata[247]));
Q_AN02 U985 ( .A0(n615), .A1(n368), .Z(rdata[246]));
Q_AN02 U986 ( .A0(n615), .A1(n369), .Z(rdata[245]));
Q_AN02 U987 ( .A0(n615), .A1(n370), .Z(rdata[244]));
Q_AN02 U988 ( .A0(n615), .A1(n371), .Z(rdata[243]));
Q_AN02 U989 ( .A0(n615), .A1(n372), .Z(rdata[242]));
Q_AN02 U990 ( .A0(n615), .A1(n373), .Z(rdata[241]));
Q_AN02 U991 ( .A0(n615), .A1(n374), .Z(rdata[240]));
Q_AN02 U992 ( .A0(n615), .A1(n375), .Z(rdata[239]));
Q_AN02 U993 ( .A0(n615), .A1(n376), .Z(rdata[238]));
Q_AN02 U994 ( .A0(n615), .A1(n377), .Z(rdata[237]));
Q_AN02 U995 ( .A0(n615), .A1(n378), .Z(rdata[236]));
Q_AN02 U996 ( .A0(n615), .A1(n379), .Z(rdata[235]));
Q_AN02 U997 ( .A0(n615), .A1(n380), .Z(rdata[234]));
Q_AN02 U998 ( .A0(n615), .A1(n381), .Z(rdata[233]));
Q_AN02 U999 ( .A0(n615), .A1(n382), .Z(rdata[232]));
Q_AN02 U1000 ( .A0(n615), .A1(n383), .Z(rdata[231]));
Q_AN02 U1001 ( .A0(n615), .A1(n384), .Z(rdata[230]));
Q_AN02 U1002 ( .A0(n615), .A1(n385), .Z(rdata[229]));
Q_AN02 U1003 ( .A0(n615), .A1(n386), .Z(rdata[228]));
Q_AN02 U1004 ( .A0(n615), .A1(n387), .Z(rdata[227]));
Q_AN02 U1005 ( .A0(n615), .A1(n388), .Z(rdata[226]));
Q_AN02 U1006 ( .A0(n615), .A1(n389), .Z(rdata[225]));
Q_AN02 U1007 ( .A0(n615), .A1(n390), .Z(rdata[224]));
Q_AN02 U1008 ( .A0(n615), .A1(n391), .Z(rdata[223]));
Q_AN02 U1009 ( .A0(n615), .A1(n392), .Z(rdata[222]));
Q_AN02 U1010 ( .A0(n615), .A1(n393), .Z(rdata[221]));
Q_AN02 U1011 ( .A0(n615), .A1(n394), .Z(rdata[220]));
Q_AN02 U1012 ( .A0(n615), .A1(n395), .Z(rdata[219]));
Q_AN02 U1013 ( .A0(n615), .A1(n396), .Z(rdata[218]));
Q_AN02 U1014 ( .A0(n615), .A1(n397), .Z(rdata[217]));
Q_AN02 U1015 ( .A0(n615), .A1(n398), .Z(rdata[216]));
Q_AN02 U1016 ( .A0(n615), .A1(n399), .Z(rdata[215]));
Q_AN02 U1017 ( .A0(n615), .A1(n400), .Z(rdata[214]));
Q_AN02 U1018 ( .A0(n615), .A1(n401), .Z(rdata[213]));
Q_AN02 U1019 ( .A0(n615), .A1(n402), .Z(rdata[212]));
Q_AN02 U1020 ( .A0(n615), .A1(n403), .Z(rdata[211]));
Q_AN02 U1021 ( .A0(n615), .A1(n404), .Z(rdata[210]));
Q_AN02 U1022 ( .A0(n615), .A1(n405), .Z(rdata[209]));
Q_AN02 U1023 ( .A0(n615), .A1(n406), .Z(rdata[208]));
Q_AN02 U1024 ( .A0(n615), .A1(n407), .Z(rdata[207]));
Q_AN02 U1025 ( .A0(n615), .A1(n408), .Z(rdata[206]));
Q_AN02 U1026 ( .A0(n615), .A1(n409), .Z(rdata[205]));
Q_AN02 U1027 ( .A0(n615), .A1(n410), .Z(rdata[204]));
Q_AN02 U1028 ( .A0(n615), .A1(n411), .Z(rdata[203]));
Q_AN02 U1029 ( .A0(n615), .A1(n412), .Z(rdata[202]));
Q_AN02 U1030 ( .A0(n615), .A1(n413), .Z(rdata[201]));
Q_AN02 U1031 ( .A0(n615), .A1(n414), .Z(rdata[200]));
Q_AN02 U1032 ( .A0(n615), .A1(n415), .Z(rdata[199]));
Q_AN02 U1033 ( .A0(n615), .A1(n416), .Z(rdata[198]));
Q_AN02 U1034 ( .A0(n615), .A1(n417), .Z(rdata[197]));
Q_AN02 U1035 ( .A0(n615), .A1(n418), .Z(rdata[196]));
Q_AN02 U1036 ( .A0(n615), .A1(n419), .Z(rdata[195]));
Q_AN02 U1037 ( .A0(n615), .A1(n420), .Z(rdata[194]));
Q_AN02 U1038 ( .A0(n615), .A1(n421), .Z(rdata[193]));
Q_AN02 U1039 ( .A0(n615), .A1(n422), .Z(rdata[192]));
Q_AN02 U1040 ( .A0(n615), .A1(n423), .Z(rdata[191]));
Q_AN02 U1041 ( .A0(n615), .A1(n424), .Z(rdata[190]));
Q_AN02 U1042 ( .A0(n615), .A1(n425), .Z(rdata[189]));
Q_AN02 U1043 ( .A0(n615), .A1(n426), .Z(rdata[188]));
Q_AN02 U1044 ( .A0(n615), .A1(n427), .Z(rdata[187]));
Q_AN02 U1045 ( .A0(n615), .A1(n428), .Z(rdata[186]));
Q_AN02 U1046 ( .A0(n615), .A1(n429), .Z(rdata[185]));
Q_AN02 U1047 ( .A0(n615), .A1(n430), .Z(rdata[184]));
Q_AN02 U1048 ( .A0(n615), .A1(n431), .Z(rdata[183]));
Q_AN02 U1049 ( .A0(n615), .A1(n432), .Z(rdata[182]));
Q_AN02 U1050 ( .A0(n615), .A1(n433), .Z(rdata[181]));
Q_AN02 U1051 ( .A0(n615), .A1(n434), .Z(rdata[180]));
Q_AN02 U1052 ( .A0(n615), .A1(n435), .Z(rdata[179]));
Q_AN02 U1053 ( .A0(n615), .A1(n436), .Z(rdata[178]));
Q_AN02 U1054 ( .A0(n615), .A1(n437), .Z(rdata[177]));
Q_AN02 U1055 ( .A0(n615), .A1(n438), .Z(rdata[176]));
Q_AN02 U1056 ( .A0(n615), .A1(n439), .Z(rdata[175]));
Q_AN02 U1057 ( .A0(n615), .A1(n440), .Z(rdata[174]));
Q_AN02 U1058 ( .A0(n615), .A1(n441), .Z(rdata[173]));
Q_AN02 U1059 ( .A0(n615), .A1(n442), .Z(rdata[172]));
Q_AN02 U1060 ( .A0(n615), .A1(n443), .Z(rdata[171]));
Q_AN02 U1061 ( .A0(n615), .A1(n444), .Z(rdata[170]));
Q_AN02 U1062 ( .A0(n615), .A1(n445), .Z(rdata[169]));
Q_AN02 U1063 ( .A0(n615), .A1(n446), .Z(rdata[168]));
Q_AN02 U1064 ( .A0(n615), .A1(n447), .Z(rdata[167]));
Q_AN02 U1065 ( .A0(n615), .A1(n448), .Z(rdata[166]));
Q_AN02 U1066 ( .A0(n615), .A1(n449), .Z(rdata[165]));
Q_AN02 U1067 ( .A0(n615), .A1(n450), .Z(rdata[164]));
Q_AN02 U1068 ( .A0(n615), .A1(n451), .Z(rdata[163]));
Q_AN02 U1069 ( .A0(n615), .A1(n452), .Z(rdata[162]));
Q_AN02 U1070 ( .A0(n615), .A1(n453), .Z(rdata[161]));
Q_AN02 U1071 ( .A0(n615), .A1(n454), .Z(rdata[160]));
Q_AN02 U1072 ( .A0(n615), .A1(n455), .Z(rdata[159]));
Q_AN02 U1073 ( .A0(n615), .A1(n456), .Z(rdata[158]));
Q_AN02 U1074 ( .A0(n615), .A1(n457), .Z(rdata[157]));
Q_AN02 U1075 ( .A0(n615), .A1(n458), .Z(rdata[156]));
Q_AN02 U1076 ( .A0(n615), .A1(n459), .Z(rdata[155]));
Q_AN02 U1077 ( .A0(n615), .A1(n460), .Z(rdata[154]));
Q_AN02 U1078 ( .A0(n615), .A1(n461), .Z(rdata[153]));
Q_AN02 U1079 ( .A0(n615), .A1(n462), .Z(rdata[152]));
Q_AN02 U1080 ( .A0(n615), .A1(n463), .Z(rdata[151]));
Q_AN02 U1081 ( .A0(n615), .A1(n464), .Z(rdata[150]));
Q_AN02 U1082 ( .A0(n615), .A1(n465), .Z(rdata[149]));
Q_AN02 U1083 ( .A0(n615), .A1(n466), .Z(rdata[148]));
Q_AN02 U1084 ( .A0(n615), .A1(n467), .Z(rdata[147]));
Q_AN02 U1085 ( .A0(n615), .A1(n468), .Z(rdata[146]));
Q_AN02 U1086 ( .A0(n615), .A1(n469), .Z(rdata[145]));
Q_AN02 U1087 ( .A0(n615), .A1(n470), .Z(rdata[144]));
Q_AN02 U1088 ( .A0(n615), .A1(n471), .Z(rdata[143]));
Q_AN02 U1089 ( .A0(n615), .A1(n472), .Z(rdata[142]));
Q_AN02 U1090 ( .A0(n615), .A1(n473), .Z(rdata[141]));
Q_AN02 U1091 ( .A0(n615), .A1(n474), .Z(rdata[140]));
Q_AN02 U1092 ( .A0(n615), .A1(n475), .Z(rdata[139]));
Q_AN02 U1093 ( .A0(n615), .A1(n476), .Z(rdata[138]));
Q_AN02 U1094 ( .A0(n615), .A1(n477), .Z(rdata[137]));
Q_AN02 U1095 ( .A0(n615), .A1(n478), .Z(rdata[136]));
Q_AN02 U1096 ( .A0(n615), .A1(n479), .Z(rdata[135]));
Q_AN02 U1097 ( .A0(n615), .A1(n480), .Z(rdata[134]));
Q_AN02 U1098 ( .A0(n615), .A1(n481), .Z(rdata[133]));
Q_AN02 U1099 ( .A0(n615), .A1(n482), .Z(rdata[132]));
Q_AN02 U1100 ( .A0(n615), .A1(n483), .Z(rdata[131]));
Q_AN02 U1101 ( .A0(n615), .A1(n484), .Z(rdata[130]));
Q_AN02 U1102 ( .A0(n615), .A1(n485), .Z(rdata[129]));
Q_AN02 U1103 ( .A0(n615), .A1(n486), .Z(rdata[128]));
Q_AN02 U1104 ( .A0(n615), .A1(n487), .Z(rdata[127]));
Q_AN02 U1105 ( .A0(n615), .A1(n488), .Z(rdata[126]));
Q_AN02 U1106 ( .A0(n615), .A1(n489), .Z(rdata[125]));
Q_AN02 U1107 ( .A0(n615), .A1(n490), .Z(rdata[124]));
Q_AN02 U1108 ( .A0(n615), .A1(n491), .Z(rdata[123]));
Q_AN02 U1109 ( .A0(n615), .A1(n492), .Z(rdata[122]));
Q_AN02 U1110 ( .A0(n615), .A1(n493), .Z(rdata[121]));
Q_AN02 U1111 ( .A0(n615), .A1(n494), .Z(rdata[120]));
Q_AN02 U1112 ( .A0(n615), .A1(n495), .Z(rdata[119]));
Q_AN02 U1113 ( .A0(n615), .A1(n496), .Z(rdata[118]));
Q_AN02 U1114 ( .A0(n615), .A1(n497), .Z(rdata[117]));
Q_AN02 U1115 ( .A0(n615), .A1(n498), .Z(rdata[116]));
Q_AN02 U1116 ( .A0(n615), .A1(n499), .Z(rdata[115]));
Q_AN02 U1117 ( .A0(n615), .A1(n500), .Z(rdata[114]));
Q_AN02 U1118 ( .A0(n615), .A1(n501), .Z(rdata[113]));
Q_AN02 U1119 ( .A0(n615), .A1(n502), .Z(rdata[112]));
Q_AN02 U1120 ( .A0(n615), .A1(n503), .Z(rdata[111]));
Q_AN02 U1121 ( .A0(n615), .A1(n504), .Z(rdata[110]));
Q_AN02 U1122 ( .A0(n615), .A1(n505), .Z(rdata[109]));
Q_AN02 U1123 ( .A0(n615), .A1(n506), .Z(rdata[108]));
Q_AN02 U1124 ( .A0(n615), .A1(n507), .Z(rdata[107]));
Q_AN02 U1125 ( .A0(n615), .A1(n508), .Z(rdata[106]));
Q_AN02 U1126 ( .A0(n615), .A1(n509), .Z(rdata[105]));
Q_AN02 U1127 ( .A0(n615), .A1(n510), .Z(rdata[104]));
Q_AN02 U1128 ( .A0(n615), .A1(n511), .Z(rdata[103]));
Q_AN02 U1129 ( .A0(n615), .A1(n512), .Z(rdata[102]));
Q_AN02 U1130 ( .A0(n615), .A1(n513), .Z(rdata[101]));
Q_AN02 U1131 ( .A0(n615), .A1(n514), .Z(rdata[100]));
Q_AN02 U1132 ( .A0(n615), .A1(n515), .Z(rdata[99]));
Q_AN02 U1133 ( .A0(n615), .A1(n516), .Z(rdata[98]));
Q_AN02 U1134 ( .A0(n615), .A1(n517), .Z(rdata[97]));
Q_AN02 U1135 ( .A0(n615), .A1(n518), .Z(rdata[96]));
Q_AN02 U1136 ( .A0(n615), .A1(n519), .Z(rdata[95]));
Q_AN02 U1137 ( .A0(n615), .A1(n520), .Z(rdata[94]));
Q_AN02 U1138 ( .A0(n615), .A1(n521), .Z(rdata[93]));
Q_AN02 U1139 ( .A0(n615), .A1(n522), .Z(rdata[92]));
Q_AN02 U1140 ( .A0(n615), .A1(n523), .Z(rdata[91]));
Q_AN02 U1141 ( .A0(n615), .A1(n524), .Z(rdata[90]));
Q_AN02 U1142 ( .A0(n615), .A1(n525), .Z(rdata[89]));
Q_AN02 U1143 ( .A0(n615), .A1(n526), .Z(rdata[88]));
Q_AN02 U1144 ( .A0(n615), .A1(n527), .Z(rdata[87]));
Q_AN02 U1145 ( .A0(n615), .A1(n528), .Z(rdata[86]));
Q_AN02 U1146 ( .A0(n615), .A1(n529), .Z(rdata[85]));
Q_AN02 U1147 ( .A0(n615), .A1(n530), .Z(rdata[84]));
Q_AN02 U1148 ( .A0(n615), .A1(n531), .Z(rdata[83]));
Q_AN02 U1149 ( .A0(n615), .A1(n532), .Z(rdata[82]));
Q_AN02 U1150 ( .A0(n615), .A1(n533), .Z(rdata[81]));
Q_AN02 U1151 ( .A0(n615), .A1(n534), .Z(rdata[80]));
Q_AN02 U1152 ( .A0(n615), .A1(n535), .Z(rdata[79]));
Q_AN02 U1153 ( .A0(n615), .A1(n536), .Z(rdata[78]));
Q_AN02 U1154 ( .A0(n615), .A1(n537), .Z(rdata[77]));
Q_AN02 U1155 ( .A0(n615), .A1(n538), .Z(rdata[76]));
Q_AN02 U1156 ( .A0(n615), .A1(n539), .Z(rdata[75]));
Q_AN02 U1157 ( .A0(n615), .A1(n540), .Z(rdata[74]));
Q_AN02 U1158 ( .A0(n615), .A1(n541), .Z(rdata[73]));
Q_AN02 U1159 ( .A0(n615), .A1(n542), .Z(rdata[72]));
Q_AN02 U1160 ( .A0(n615), .A1(n543), .Z(rdata[71]));
Q_AN02 U1161 ( .A0(n615), .A1(n544), .Z(rdata[70]));
Q_AN02 U1162 ( .A0(n615), .A1(n545), .Z(rdata[69]));
Q_AN02 U1163 ( .A0(n615), .A1(n546), .Z(rdata[68]));
Q_AN02 U1164 ( .A0(n615), .A1(n547), .Z(rdata[67]));
Q_AN02 U1165 ( .A0(n615), .A1(n548), .Z(rdata[66]));
Q_AN02 U1166 ( .A0(n615), .A1(n549), .Z(rdata[65]));
Q_AN02 U1167 ( .A0(n615), .A1(n550), .Z(rdata[64]));
Q_AN02 U1168 ( .A0(n615), .A1(n551), .Z(rdata[63]));
Q_AN02 U1169 ( .A0(n615), .A1(n552), .Z(rdata[62]));
Q_AN02 U1170 ( .A0(n615), .A1(n553), .Z(rdata[61]));
Q_AN02 U1171 ( .A0(n615), .A1(n554), .Z(rdata[60]));
Q_AN02 U1172 ( .A0(n615), .A1(n555), .Z(rdata[59]));
Q_AN02 U1173 ( .A0(n615), .A1(n556), .Z(rdata[58]));
Q_AN02 U1174 ( .A0(n615), .A1(n557), .Z(rdata[57]));
Q_AN02 U1175 ( .A0(n615), .A1(n558), .Z(rdata[56]));
Q_AN02 U1176 ( .A0(n615), .A1(n559), .Z(rdata[55]));
Q_AN02 U1177 ( .A0(n615), .A1(n560), .Z(rdata[54]));
Q_AN02 U1178 ( .A0(n615), .A1(n561), .Z(rdata[53]));
Q_AN02 U1179 ( .A0(n615), .A1(n562), .Z(rdata[52]));
Q_AN02 U1180 ( .A0(n615), .A1(n563), .Z(rdata[51]));
Q_AN02 U1181 ( .A0(n615), .A1(n564), .Z(rdata[50]));
Q_AN02 U1182 ( .A0(n615), .A1(n565), .Z(rdata[49]));
Q_AN02 U1183 ( .A0(n615), .A1(n566), .Z(rdata[48]));
Q_AN02 U1184 ( .A0(n615), .A1(n567), .Z(rdata[47]));
Q_AN02 U1185 ( .A0(n615), .A1(n568), .Z(rdata[46]));
Q_AN02 U1186 ( .A0(n615), .A1(n569), .Z(rdata[45]));
Q_AN02 U1187 ( .A0(n615), .A1(n570), .Z(rdata[44]));
Q_AN02 U1188 ( .A0(n615), .A1(n571), .Z(rdata[43]));
Q_AN02 U1189 ( .A0(n615), .A1(n572), .Z(rdata[42]));
Q_AN02 U1190 ( .A0(n615), .A1(n573), .Z(rdata[41]));
Q_AN02 U1191 ( .A0(n615), .A1(n574), .Z(rdata[40]));
Q_AN02 U1192 ( .A0(n615), .A1(n575), .Z(rdata[39]));
Q_AN02 U1193 ( .A0(n615), .A1(n576), .Z(rdata[38]));
Q_AN02 U1194 ( .A0(n615), .A1(n577), .Z(rdata[37]));
Q_AN02 U1195 ( .A0(n615), .A1(n578), .Z(rdata[36]));
Q_AN02 U1196 ( .A0(n615), .A1(n579), .Z(rdata[35]));
Q_AN02 U1197 ( .A0(n615), .A1(n580), .Z(rdata[34]));
Q_AN02 U1198 ( .A0(n615), .A1(n581), .Z(rdata[33]));
Q_AN02 U1199 ( .A0(n615), .A1(n582), .Z(rdata[32]));
Q_AN02 U1200 ( .A0(n615), .A1(n583), .Z(rdata[31]));
Q_AN02 U1201 ( .A0(n615), .A1(n584), .Z(rdata[30]));
Q_AN02 U1202 ( .A0(n615), .A1(n585), .Z(rdata[29]));
Q_AN02 U1203 ( .A0(n615), .A1(n586), .Z(rdata[28]));
Q_AN02 U1204 ( .A0(n615), .A1(n587), .Z(rdata[27]));
Q_AN02 U1205 ( .A0(n615), .A1(n588), .Z(rdata[26]));
Q_AN02 U1206 ( .A0(n615), .A1(n589), .Z(rdata[25]));
Q_AN02 U1207 ( .A0(n615), .A1(n590), .Z(rdata[24]));
Q_AN02 U1208 ( .A0(n615), .A1(n591), .Z(rdata[23]));
Q_AN02 U1209 ( .A0(n615), .A1(n592), .Z(rdata[22]));
Q_AN02 U1210 ( .A0(n615), .A1(n593), .Z(rdata[21]));
Q_AN02 U1211 ( .A0(n615), .A1(n594), .Z(rdata[20]));
Q_AN02 U1212 ( .A0(n615), .A1(n595), .Z(rdata[19]));
Q_AN02 U1213 ( .A0(n615), .A1(n596), .Z(rdata[18]));
Q_AN02 U1214 ( .A0(n615), .A1(n597), .Z(rdata[17]));
Q_AN02 U1215 ( .A0(n615), .A1(n598), .Z(rdata[16]));
Q_AN02 U1216 ( .A0(n615), .A1(n599), .Z(rdata[15]));
Q_AN02 U1217 ( .A0(n615), .A1(n600), .Z(rdata[14]));
Q_AN02 U1218 ( .A0(n615), .A1(n601), .Z(rdata[13]));
Q_AN02 U1219 ( .A0(n615), .A1(n602), .Z(rdata[12]));
Q_AN02 U1220 ( .A0(n615), .A1(n603), .Z(rdata[11]));
Q_AN02 U1221 ( .A0(n615), .A1(n604), .Z(rdata[10]));
Q_AN02 U1222 ( .A0(n615), .A1(n605), .Z(rdata[9]));
Q_AN02 U1223 ( .A0(n615), .A1(n606), .Z(rdata[8]));
Q_AN02 U1224 ( .A0(n615), .A1(n607), .Z(rdata[7]));
Q_AN02 U1225 ( .A0(n615), .A1(n608), .Z(rdata[6]));
Q_AN02 U1226 ( .A0(n615), .A1(n609), .Z(rdata[5]));
Q_AN02 U1227 ( .A0(n615), .A1(n610), .Z(rdata[4]));
Q_AN02 U1228 ( .A0(n615), .A1(n611), .Z(rdata[3]));
Q_AN02 U1229 ( .A0(n615), .A1(n612), .Z(rdata[2]));
Q_AN02 U1230 ( .A0(n615), .A1(n613), .Z(rdata[1]));
Q_AN02 U1231 ( .A0(n615), .A1(n614), .Z(rdata[0]));
Q_INV U1232 ( .A(full), .Z(n2));
Q_AN02 U1233 ( .A0(wen), .A1(n2), .Z(n3));
nx_fifo_ctrl_xcm37 \depth_n.fifo_ctrl ( .empty( empty), .full( full), 
	.used_slots( used_slots[2:0]), .free_slots( free_slots[2:0]), 
	.rptr( \depth_n.rptr [1:0]), .wptr( \depth_n.wptr [1:0]), 
	.underflow( \depth_n._zy_simnet_underflow_2_w$ ), .overflow( 
	\depth_n._zy_simnet_overflow_3_w$ ), .clk( clk), .rst_n( rst_n), 
	.wen( wen), .ren( ren), .clear( clear));
ixc_assign \depth_n._zz_strnp_1 ( overflow, 
	\depth_n._zy_simnet_overflow_3_w$ );
ixc_assign \depth_n._zz_strnp_0 ( underflow, 
	\depth_n._zy_simnet_underflow_2_w$ );
`ifdef CBV

reg [610:0] \depth_n.r_data  [3:0];
initial begin: U1237
  integer i;
  for (i=3; i>=0; i=i-1) \depth_n.r_data [i] =
`ifdef CBV_MEM_INIT1
  {611{1'b1}};
`else
  611'b0;
`endif
end
reg [610:0] n1236;
assign {n4, n5, n6, n7, n8, n9, n10,
n11, n12, n13, n14, n15, n16, n17, n18,
n19, n20, n21, n22, n23, n24, n25, n26,
n27, n28, n29, n30, n31, n32, n33, n34,
n35, n36, n37, n38, n39, n40, n41, n42,
n43, n44, n45, n46, n47, n48, n49, n50,
n51, n52, n53, n54, n55, n56, n57, n58,
n59, n60, n61, n62, n63, n64, n65, n66,
n67, n68, n69, n70, n71, n72, n73, n74,
n75, n76, n77, n78, n79, n80, n81, n82,
n83, n84, n85, n86, n87, n88, n89, n90,
n91, n92, n93, n94, n95, n96, n97, n98,
n99, n100, n101, n102, n103, n104, n105, n106,
n107, n108, n109, n110, n111, n112, n113, n114,
n115, n116, n117, n118, n119, n120, n121, n122,
n123, n124, n125, n126, n127, n128, n129, n130,
n131, n132, n133, n134, n135, n136, n137, n138,
n139, n140, n141, n142, n143, n144, n145, n146,
n147, n148, n149, n150, n151, n152, n153, n154,
n155, n156, n157, n158, n159, n160, n161, n162,
n163, n164, n165, n166, n167, n168, n169, n170,
n171, n172, n173, n174, n175, n176, n177, n178,
n179, n180, n181, n182, n183, n184, n185, n186,
n187, n188, n189, n190, n191, n192, n193, n194,
n195, n196, n197, n198, n199, n200, n201, n202,
n203, n204, n205, n206, n207, n208, n209, n210,
n211, n212, n213, n214, n215, n216, n217, n218,
n219, n220, n221, n222, n223, n224, n225, n226,
n227, n228, n229, n230, n231, n232, n233, n234,
n235, n236, n237, n238, n239, n240, n241, n242,
n243, n244, n245, n246, n247, n248, n249, n250,
n251, n252, n253, n254, n255, n256, n257, n258,
n259, n260, n261, n262, n263, n264, n265, n266,
n267, n268, n269, n270, n271, n272, n273, n274,
n275, n276, n277, n278, n279, n280, n281, n282,
n283, n284, n285, n286, n287, n288, n289, n290,
n291, n292, n293, n294, n295, n296, n297, n298,
n299, n300, n301, n302, n303, n304, n305, n306,
n307, n308, n309, n310, n311, n312, n313, n314,
n315, n316, n317, n318, n319, n320, n321, n322,
n323, n324, n325, n326, n327, n328, n329, n330,
n331, n332, n333, n334, n335, n336, n337, n338,
n339, n340, n341, n342, n343, n344, n345, n346,
n347, n348, n349, n350, n351, n352, n353, n354,
n355, n356, n357, n358, n359, n360, n361, n362,
n363, n364, n365, n366, n367, n368, n369, n370,
n371, n372, n373, n374, n375, n376, n377, n378,
n379, n380, n381, n382, n383, n384, n385, n386,
n387, n388, n389, n390, n391, n392, n393, n394,
n395, n396, n397, n398, n399, n400, n401, n402,
n403, n404, n405, n406, n407, n408, n409, n410,
n411, n412, n413, n414, n415, n416, n417, n418,
n419, n420, n421, n422, n423, n424, n425, n426,
n427, n428, n429, n430, n431, n432, n433, n434,
n435, n436, n437, n438, n439, n440, n441, n442,
n443, n444, n445, n446, n447, n448, n449, n450,
n451, n452, n453, n454, n455, n456, n457, n458,
n459, n460, n461, n462, n463, n464, n465, n466,
n467, n468, n469, n470, n471, n472, n473, n474,
n475, n476, n477, n478, n479, n480, n481, n482,
n483, n484, n485, n486, n487, n488, n489, n490,
n491, n492, n493, n494, n495, n496, n497, n498,
n499, n500, n501, n502, n503, n504, n505, n506,
n507, n508, n509, n510, n511, n512, n513, n514,
n515, n516, n517, n518, n519, n520, n521, n522,
n523, n524, n525, n526, n527, n528, n529, n530,
n531, n532, n533, n534, n535, n536, n537, n538,
n539, n540, n541, n542, n543, n544, n545, n546,
n547, n548, n549, n550, n551, n552, n553, n554,
n555, n556, n557, n558, n559, n560, n561, n562,
n563, n564, n565, n566, n567, n568, n569, n570,
n571, n572, n573, n574, n575, n576, n577, n578,
n579, n580, n581, n582, n583, n584, n585, n586,
n587, n588, n589, n590, n591, n592, n593, n594,
n595, n596, n597, n598, n599, n600, n601, n602,
n603, n604, n605, n606, n607, n608, n609, n610,
n611, n612, n613, n614} = n1236; 
always @(n623 or n622 or n1234 or n1233 or n1232
 or n1231 or n1230 or n1229 or n1228 or n1227 or n1226 or n1225 or n1224
 or n1223 or n1222 or n1221 or n1220 or n1219 or n1218 or n1217 or n1216
 or n1215 or n1214 or n1213 or n1212 or n1211 or n1210 or n1209 or n1208
 or n1207 or n1206 or n1205 or n1204 or n1203 or n1202 or n1201 or n1200
 or n1199 or n1198 or n1197 or n1196 or n1195 or n1194 or n1193 or n1192
 or n1191 or n1190 or n1189 or n1188 or n1187 or n1186 or n1185 or n1184
 or n1183 or n1182 or n1181 or n1180 or n1179 or n1178 or n1177 or n1176
 or n1175 or n1174 or n1173 or n1172 or n1171 or n1170 or n1169 or n1168
 or n1167 or n1166 or n1165 or n1164 or n1163 or n1162 or n1161 or n1160
 or n1159 or n1158 or n1157 or n1156 or n1155 or n1154 or n1153 or n1152
 or n1151 or n1150 or n1149 or n1148 or n1147 or n1146 or n1145 or n1144
 or n1143 or n1142 or n1141 or n1140 or n1139 or n1138 or n1137 or n1136
 or n1135 or n1134 or n1133 or n1132 or n1131 or n1130 or n1129 or n1128
 or n1127 or n1126 or n1125 or n1124 or n1123 or n1122 or n1121 or n1120
 or n1119 or n1118 or n1117 or n1116 or n1115 or n1114 or n1113 or n1112
 or n1111 or n1110 or n1109 or n1108 or n1107 or n1106 or n1105 or n1104
 or n1103 or n1102 or n1101 or n1100 or n1099 or n1098 or n1097 or n1096
 or n1095 or n1094 or n1093 or n1092 or n1091 or n1090 or n1089 or n1088
 or n1087 or n1086 or n1085 or n1084 or n1083 or n1082 or n1081 or n1080
 or n1079 or n1078 or n1077 or n1076 or n1075 or n1074 or n1073 or n1072
 or n1071 or n1070 or n1069 or n1068 or n1067 or n1066 or n1065 or n1064
 or n1063 or n1062 or n1061 or n1060 or n1059 or n1058 or n1057 or n1056
 or n1055 or n1054 or n1053 or n1052 or n1051 or n1050 or n1049 or n1048
 or n1047 or n1046 or n1045 or n1044 or n1043 or n1042 or n1041 or n1040
 or n1039 or n1038 or n1037 or n1036 or n1035 or n1034 or n1033 or n1032
 or n1031 or n1030 or n1029 or n1028 or n1027 or n1026 or n1025 or n1024
 or n1023 or n1022 or n1021 or n1020 or n1019 or n1018 or n1017 or n1016
 or n1015 or n1014 or n1013 or n1012 or n1011 or n1010 or n1009 or n1008
 or n1007 or n1006 or n1005 or n1004 or n1003 or n1002 or n1001 or n1000
 or n999 or n998 or n997 or n996 or n995 or n994 or n993 or n992
 or n991 or n990 or n989 or n988 or n987 or n986 or n985 or n984
 or n983 or n982 or n981 or n980 or n979 or n978 or n977 or n976
 or n975 or n974 or n973 or n972 or n971 or n970 or n969 or n968
 or n967 or n966 or n965 or n964 or n963 or n962 or n961 or n960
 or n959 or n958 or n957 or n956 or n955 or n954 or n953 or n952
 or n951 or n950 or n949 or n948 or n947 or n946 or n945 or n944
 or n943 or n942 or n941 or n940 or n939 or n938 or n937 or n936
 or n935 or n934 or n933 or n932 or n931 or n930 or n929 or n928
 or n927 or n926 or n925 or n924 or n923 or n922 or n921 or n920
 or n919 or n918 or n917 or n916 or n915 or n914 or n913 or n912
 or n911 or n910 or n909 or n908 or n907 or n906 or n905 or n904
 or n903 or n902 or n901 or n900 or n899 or n898 or n897 or n896
 or n895 or n894 or n893 or n892 or n891 or n890 or n889 or n888
 or n887 or n886 or n885 or n884 or n883 or n882 or n881 or n880
 or n879 or n878 or n877 or n876 or n875 or n874 or n873 or n872
 or n871 or n870 or n869 or n868 or n867 or n866 or n865 or n864
 or n863 or n862 or n861 or n860 or n859 or n858 or n857 or n856
 or n855 or n854 or n853 or n852 or n851 or n850 or n849 or n848
 or n847 or n846 or n845 or n844 or n843 or n842 or n841 or n840
 or n839 or n838 or n837 or n836 or n835 or n834 or n833 or n832
 or n831 or n830 or n829 or n828 or n827 or n826 or n825 or n824
 or n823 or n822 or n821 or n820 or n819 or n818 or n817 or n816
 or n815 or n814 or n813 or n812 or n811 or n810 or n809 or n808
 or n807 or n806 or n805 or n804 or n803 or n802 or n801 or n800
 or n799 or n798 or n797 or n796 or n795 or n794 or n793 or n792
 or n791 or n790 or n789 or n788 or n787 or n786 or n785 or n784
 or n783 or n782 or n781 or n780 or n779 or n778 or n777 or n776
 or n775 or n774 or n773 or n772 or n771 or n770 or n769 or n768
 or n767 or n766 or n765 or n764 or n763 or n762 or n761 or n760
 or n759 or n758 or n757 or n756 or n755 or n754 or n753 or n752
 or n751 or n750 or n749 or n748 or n747 or n746 or n745 or n744
 or n743 or n742 or n741 or n740 or n739 or n738 or n737 or n736
 or n735 or n734 or n733 or n732 or n731 or n730 or n729 or n728
 or n727 or n726 or n725 or n724 or n723 or n722 or n721 or n720
 or n719 or n718 or n717 or n716 or n715 or n714 or n713 or n712
 or n711 or n710 or n709 or n708 or n707 or n706 or n705 or n704
 or n703 or n702 or n701 or n700 or n699 or n698 or n697 or n696
 or n695 or n694 or n693 or n692 or n691 or n690 or n689 or n688
 or n687 or n686 or n685 or n684 or n683 or n682 or n681 or n680
 or n679 or n678 or n677 or n676 or n675 or n674 or n673 or n672
 or n671 or n670 or n669 or n668 or n667 or n666 or n665 or n664
 or n663 or n662 or n661 or n660 or n659 or n658 or n657 or n656
 or n655 or n654 or n653 or n652 or n651 or n650 or n649 or n648
 or n647 or n646 or n645 or n644 or n643 or n642 or n641 or n640
 or n639 or n638 or n637 or n636 or n635 or n634 or n633 or n632
 or n631 or n630 or n629 or n628 or n627 or n626 or n625 or n624
 or n621 or \depth_n.rptr [1] or \depth_n.rptr [0])
#0 begin
if (n621)
\depth_n.r_data [{n623, n622}] =
{n1234, n1233, n1232, n1231, n1230,
 n1229, n1228, n1227, n1226, n1225, n1224, n1223, n1222,
 n1221, n1220, n1219, n1218, n1217, n1216, n1215, n1214,
 n1213, n1212, n1211, n1210, n1209, n1208, n1207, n1206,
 n1205, n1204, n1203, n1202, n1201, n1200, n1199, n1198,
 n1197, n1196, n1195, n1194, n1193, n1192, n1191, n1190,
 n1189, n1188, n1187, n1186, n1185, n1184, n1183, n1182,
 n1181, n1180, n1179, n1178, n1177, n1176, n1175, n1174,
 n1173, n1172, n1171, n1170, n1169, n1168, n1167, n1166,
 n1165, n1164, n1163, n1162, n1161, n1160, n1159, n1158,
 n1157, n1156, n1155, n1154, n1153, n1152, n1151, n1150,
 n1149, n1148, n1147, n1146, n1145, n1144, n1143, n1142,
 n1141, n1140, n1139, n1138, n1137, n1136, n1135, n1134,
 n1133, n1132, n1131, n1130, n1129, n1128, n1127, n1126,
 n1125, n1124, n1123, n1122, n1121, n1120, n1119, n1118,
 n1117, n1116, n1115, n1114, n1113, n1112, n1111, n1110,
 n1109, n1108, n1107, n1106, n1105, n1104, n1103, n1102,
 n1101, n1100, n1099, n1098, n1097, n1096, n1095, n1094,
 n1093, n1092, n1091, n1090, n1089, n1088, n1087, n1086,
 n1085, n1084, n1083, n1082, n1081, n1080, n1079, n1078,
 n1077, n1076, n1075, n1074, n1073, n1072, n1071, n1070,
 n1069, n1068, n1067, n1066, n1065, n1064, n1063, n1062,
 n1061, n1060, n1059, n1058, n1057, n1056, n1055, n1054,
 n1053, n1052, n1051, n1050, n1049, n1048, n1047, n1046,
 n1045, n1044, n1043, n1042, n1041, n1040, n1039, n1038,
 n1037, n1036, n1035, n1034, n1033, n1032, n1031, n1030,
 n1029, n1028, n1027, n1026, n1025, n1024, n1023, n1022,
 n1021, n1020, n1019, n1018, n1017, n1016, n1015, n1014,
 n1013, n1012, n1011, n1010, n1009, n1008, n1007, n1006,
 n1005, n1004, n1003, n1002, n1001, n1000, n999, n998,
 n997, n996, n995, n994, n993, n992, n991, n990,
 n989, n988, n987, n986, n985, n984, n983, n982,
 n981, n980, n979, n978, n977, n976, n975, n974,
 n973, n972, n971, n970, n969, n968, n967, n966,
 n965, n964, n963, n962, n961, n960, n959, n958,
 n957, n956, n955, n954, n953, n952, n951, n950,
 n949, n948, n947, n946, n945, n944, n943, n942,
 n941, n940, n939, n938, n937, n936, n935, n934,
 n933, n932, n931, n930, n929, n928, n927, n926,
 n925, n924, n923, n922, n921, n920, n919, n918,
 n917, n916, n915, n914, n913, n912, n911, n910,
 n909, n908, n907, n906, n905, n904, n903, n902,
 n901, n900, n899, n898, n897, n896, n895, n894,
 n893, n892, n891, n890, n889, n888, n887, n886,
 n885, n884, n883, n882, n881, n880, n879, n878,
 n877, n876, n875, n874, n873, n872, n871, n870,
 n869, n868, n867, n866, n865, n864, n863, n862,
 n861, n860, n859, n858, n857, n856, n855, n854,
 n853, n852, n851, n850, n849, n848, n847, n846,
 n845, n844, n843, n842, n841, n840, n839, n838,
 n837, n836, n835, n834, n833, n832, n831, n830,
 n829, n828, n827, n826, n825, n824, n823, n822,
 n821, n820, n819, n818, n817, n816, n815, n814,
 n813, n812, n811, n810, n809, n808, n807, n806,
 n805, n804, n803, n802, n801, n800, n799, n798,
 n797, n796, n795, n794, n793, n792, n791, n790,
 n789, n788, n787, n786, n785, n784, n783, n782,
 n781, n780, n779, n778, n777, n776, n775, n774,
 n773, n772, n771, n770, n769, n768, n767, n766,
 n765, n764, n763, n762, n761, n760, n759, n758,
 n757, n756, n755, n754, n753, n752, n751, n750,
 n749, n748, n747, n746, n745, n744, n743, n742,
 n741, n740, n739, n738, n737, n736, n735, n734,
 n733, n732, n731, n730, n729, n728, n727, n726,
 n725, n724, n723, n722, n721, n720, n719, n718,
 n717, n716, n715, n714, n713, n712, n711, n710,
 n709, n708, n707, n706, n705, n704, n703, n702,
 n701, n700, n699, n698, n697, n696, n695, n694,
 n693, n692, n691, n690, n689, n688, n687, n686,
 n685, n684, n683, n682, n681, n680, n679, n678,
 n677, n676, n675, n674, n673, n672, n671, n670,
 n669, n668, n667, n666, n665, n664, n663, n662,
 n661, n660, n659, n658, n657, n656, n655, n654,
 n653, n652, n651, n650, n649, n648, n647, n646,
 n645, n644, n643, n642, n641, n640, n639, n638,
 n637, n636, n635, n634, n633, n632, n631, n630,
 n629, n628, n627, n626, n625, n624};
n1236 = \depth_n.r_data [{\depth_n.rptr [1], \depth_n.rptr [0]}];
end
`else

MPW4X611 \depth_n.r_data  ( .A1(n623), .A0(n622), .DI610(n1234), .DI609(n1233), .DI608(n1232), .DI607(n1231),
 .DI606(n1230), .DI605(n1229), .DI604(n1228), .DI603(n1227), .DI602(n1226), .DI601(n1225), .DI600(n1224), .DI599(n1223),
 .DI598(n1222), .DI597(n1221), .DI596(n1220), .DI595(n1219), .DI594(n1218), .DI593(n1217), .DI592(n1216), .DI591(n1215),
 .DI590(n1214), .DI589(n1213), .DI588(n1212), .DI587(n1211), .DI586(n1210), .DI585(n1209), .DI584(n1208), .DI583(n1207),
 .DI582(n1206), .DI581(n1205), .DI580(n1204), .DI579(n1203), .DI578(n1202), .DI577(n1201), .DI576(n1200), .DI575(n1199),
 .DI574(n1198), .DI573(n1197), .DI572(n1196), .DI571(n1195), .DI570(n1194), .DI569(n1193), .DI568(n1192), .DI567(n1191),
 .DI566(n1190), .DI565(n1189), .DI564(n1188), .DI563(n1187), .DI562(n1186), .DI561(n1185), .DI560(n1184), .DI559(n1183),
 .DI558(n1182), .DI557(n1181), .DI556(n1180), .DI555(n1179), .DI554(n1178), .DI553(n1177), .DI552(n1176), .DI551(n1175),
 .DI550(n1174), .DI549(n1173), .DI548(n1172), .DI547(n1171), .DI546(n1170), .DI545(n1169), .DI544(n1168), .DI543(n1167),
 .DI542(n1166), .DI541(n1165), .DI540(n1164), .DI539(n1163), .DI538(n1162), .DI537(n1161), .DI536(n1160), .DI535(n1159),
 .DI534(n1158), .DI533(n1157), .DI532(n1156), .DI531(n1155), .DI530(n1154), .DI529(n1153), .DI528(n1152), .DI527(n1151),
 .DI526(n1150), .DI525(n1149), .DI524(n1148), .DI523(n1147), .DI522(n1146), .DI521(n1145), .DI520(n1144), .DI519(n1143),
 .DI518(n1142), .DI517(n1141), .DI516(n1140), .DI515(n1139), .DI514(n1138), .DI513(n1137), .DI512(n1136), .DI511(n1135),
 .DI510(n1134), .DI509(n1133), .DI508(n1132), .DI507(n1131), .DI506(n1130), .DI505(n1129), .DI504(n1128), .DI503(n1127),
 .DI502(n1126), .DI501(n1125), .DI500(n1124), .DI499(n1123), .DI498(n1122), .DI497(n1121), .DI496(n1120), .DI495(n1119),
 .DI494(n1118), .DI493(n1117), .DI492(n1116), .DI491(n1115), .DI490(n1114), .DI489(n1113), .DI488(n1112), .DI487(n1111),
 .DI486(n1110), .DI485(n1109), .DI484(n1108), .DI483(n1107), .DI482(n1106), .DI481(n1105), .DI480(n1104), .DI479(n1103),
 .DI478(n1102), .DI477(n1101), .DI476(n1100), .DI475(n1099), .DI474(n1098), .DI473(n1097), .DI472(n1096), .DI471(n1095),
 .DI470(n1094), .DI469(n1093), .DI468(n1092), .DI467(n1091), .DI466(n1090), .DI465(n1089), .DI464(n1088), .DI463(n1087),
 .DI462(n1086), .DI461(n1085), .DI460(n1084), .DI459(n1083), .DI458(n1082), .DI457(n1081), .DI456(n1080), .DI455(n1079),
 .DI454(n1078), .DI453(n1077), .DI452(n1076), .DI451(n1075), .DI450(n1074), .DI449(n1073), .DI448(n1072), .DI447(n1071),
 .DI446(n1070), .DI445(n1069), .DI444(n1068), .DI443(n1067), .DI442(n1066), .DI441(n1065), .DI440(n1064), .DI439(n1063),
 .DI438(n1062), .DI437(n1061), .DI436(n1060), .DI435(n1059), .DI434(n1058), .DI433(n1057), .DI432(n1056), .DI431(n1055),
 .DI430(n1054), .DI429(n1053), .DI428(n1052), .DI427(n1051), .DI426(n1050), .DI425(n1049), .DI424(n1048), .DI423(n1047),
 .DI422(n1046), .DI421(n1045), .DI420(n1044), .DI419(n1043), .DI418(n1042), .DI417(n1041), .DI416(n1040), .DI415(n1039),
 .DI414(n1038), .DI413(n1037), .DI412(n1036), .DI411(n1035), .DI410(n1034), .DI409(n1033), .DI408(n1032), .DI407(n1031),
 .DI406(n1030), .DI405(n1029), .DI404(n1028), .DI403(n1027), .DI402(n1026), .DI401(n1025), .DI400(n1024), .DI399(n1023),
 .DI398(n1022), .DI397(n1021), .DI396(n1020), .DI395(n1019), .DI394(n1018), .DI393(n1017), .DI392(n1016), .DI391(n1015),
 .DI390(n1014), .DI389(n1013), .DI388(n1012), .DI387(n1011), .DI386(n1010), .DI385(n1009), .DI384(n1008), .DI383(n1007),
 .DI382(n1006), .DI381(n1005), .DI380(n1004), .DI379(n1003), .DI378(n1002), .DI377(n1001), .DI376(n1000), .DI375(n999),
 .DI374(n998), .DI373(n997), .DI372(n996), .DI371(n995), .DI370(n994), .DI369(n993), .DI368(n992), .DI367(n991),
 .DI366(n990), .DI365(n989), .DI364(n988), .DI363(n987), .DI362(n986), .DI361(n985), .DI360(n984), .DI359(n983),
 .DI358(n982), .DI357(n981), .DI356(n980), .DI355(n979), .DI354(n978), .DI353(n977), .DI352(n976), .DI351(n975),
 .DI350(n974), .DI349(n973), .DI348(n972), .DI347(n971), .DI346(n970), .DI345(n969), .DI344(n968), .DI343(n967),
 .DI342(n966), .DI341(n965), .DI340(n964), .DI339(n963), .DI338(n962), .DI337(n961), .DI336(n960), .DI335(n959),
 .DI334(n958), .DI333(n957), .DI332(n956), .DI331(n955), .DI330(n954), .DI329(n953), .DI328(n952), .DI327(n951),
 .DI326(n950), .DI325(n949), .DI324(n948), .DI323(n947), .DI322(n946), .DI321(n945), .DI320(n944), .DI319(n943),
 .DI318(n942), .DI317(n941), .DI316(n940), .DI315(n939), .DI314(n938), .DI313(n937), .DI312(n936), .DI311(n935),
 .DI310(n934), .DI309(n933), .DI308(n932), .DI307(n931), .DI306(n930), .DI305(n929), .DI304(n928), .DI303(n927),
 .DI302(n926), .DI301(n925), .DI300(n924), .DI299(n923), .DI298(n922), .DI297(n921), .DI296(n920), .DI295(n919),
 .DI294(n918), .DI293(n917), .DI292(n916), .DI291(n915), .DI290(n914), .DI289(n913), .DI288(n912), .DI287(n911),
 .DI286(n910), .DI285(n909), .DI284(n908), .DI283(n907), .DI282(n906), .DI281(n905), .DI280(n904), .DI279(n903),
 .DI278(n902), .DI277(n901), .DI276(n900), .DI275(n899), .DI274(n898), .DI273(n897), .DI272(n896), .DI271(n895),
 .DI270(n894), .DI269(n893), .DI268(n892), .DI267(n891), .DI266(n890), .DI265(n889), .DI264(n888), .DI263(n887),
 .DI262(n886), .DI261(n885), .DI260(n884), .DI259(n883), .DI258(n882), .DI257(n881), .DI256(n880), .DI255(n879),
 .DI254(n878), .DI253(n877), .DI252(n876), .DI251(n875), .DI250(n874), .DI249(n873), .DI248(n872), .DI247(n871),
 .DI246(n870), .DI245(n869), .DI244(n868), .DI243(n867), .DI242(n866), .DI241(n865), .DI240(n864), .DI239(n863),
 .DI238(n862), .DI237(n861), .DI236(n860), .DI235(n859), .DI234(n858), .DI233(n857), .DI232(n856), .DI231(n855),
 .DI230(n854), .DI229(n853), .DI228(n852), .DI227(n851), .DI226(n850), .DI225(n849), .DI224(n848), .DI223(n847),
 .DI222(n846), .DI221(n845), .DI220(n844), .DI219(n843), .DI218(n842), .DI217(n841), .DI216(n840), .DI215(n839),
 .DI214(n838), .DI213(n837), .DI212(n836), .DI211(n835), .DI210(n834), .DI209(n833), .DI208(n832), .DI207(n831),
 .DI206(n830), .DI205(n829), .DI204(n828), .DI203(n827), .DI202(n826), .DI201(n825), .DI200(n824), .DI199(n823),
 .DI198(n822), .DI197(n821), .DI196(n820), .DI195(n819), .DI194(n818), .DI193(n817), .DI192(n816), .DI191(n815),
 .DI190(n814), .DI189(n813), .DI188(n812), .DI187(n811), .DI186(n810), .DI185(n809), .DI184(n808), .DI183(n807),
 .DI182(n806), .DI181(n805), .DI180(n804), .DI179(n803), .DI178(n802), .DI177(n801), .DI176(n800), .DI175(n799),
 .DI174(n798), .DI173(n797), .DI172(n796), .DI171(n795), .DI170(n794), .DI169(n793), .DI168(n792), .DI167(n791),
 .DI166(n790), .DI165(n789), .DI164(n788), .DI163(n787), .DI162(n786), .DI161(n785), .DI160(n784), .DI159(n783),
 .DI158(n782), .DI157(n781), .DI156(n780), .DI155(n779), .DI154(n778), .DI153(n777), .DI152(n776), .DI151(n775),
 .DI150(n774), .DI149(n773), .DI148(n772), .DI147(n771), .DI146(n770), .DI145(n769), .DI144(n768), .DI143(n767),
 .DI142(n766), .DI141(n765), .DI140(n764), .DI139(n763), .DI138(n762), .DI137(n761), .DI136(n760), .DI135(n759),
 .DI134(n758), .DI133(n757), .DI132(n756), .DI131(n755), .DI130(n754), .DI129(n753), .DI128(n752), .DI127(n751),
 .DI126(n750), .DI125(n749), .DI124(n748), .DI123(n747), .DI122(n746), .DI121(n745), .DI120(n744), .DI119(n743),
 .DI118(n742), .DI117(n741), .DI116(n740), .DI115(n739), .DI114(n738), .DI113(n737), .DI112(n736), .DI111(n735),
 .DI110(n734), .DI109(n733), .DI108(n732), .DI107(n731), .DI106(n730), .DI105(n729), .DI104(n728), .DI103(n727),
 .DI102(n726), .DI101(n725), .DI100(n724), .DI99(n723), .DI98(n722), .DI97(n721), .DI96(n720), .DI95(n719),
 .DI94(n718), .DI93(n717), .DI92(n716), .DI91(n715), .DI90(n714), .DI89(n713), .DI88(n712), .DI87(n711),
 .DI86(n710), .DI85(n709), .DI84(n708), .DI83(n707), .DI82(n706), .DI81(n705), .DI80(n704), .DI79(n703),
 .DI78(n702), .DI77(n701), .DI76(n700), .DI75(n699), .DI74(n698), .DI73(n697), .DI72(n696), .DI71(n695),
 .DI70(n694), .DI69(n693), .DI68(n692), .DI67(n691), .DI66(n690), .DI65(n689), .DI64(n688), .DI63(n687),
 .DI62(n686), .DI61(n685), .DI60(n684), .DI59(n683), .DI58(n682), .DI57(n681), .DI56(n680), .DI55(n679),
 .DI54(n678), .DI53(n677), .DI52(n676), .DI51(n675), .DI50(n674), .DI49(n673), .DI48(n672), .DI47(n671),
 .DI46(n670), .DI45(n669), .DI44(n668), .DI43(n667), .DI42(n666), .DI41(n665), .DI40(n664), .DI39(n663),
 .DI38(n662), .DI37(n661), .DI36(n660), .DI35(n659), .DI34(n658), .DI33(n657), .DI32(n656), .DI31(n655),
 .DI30(n654), .DI29(n653), .DI28(n652), .DI27(n651), .DI26(n650), .DI25(n649), .DI24(n648), .DI23(n647),
 .DI22(n646), .DI21(n645), .DI20(n644), .DI19(n643), .DI18(n642), .DI17(n641), .DI16(n640), .DI15(n639),
 .DI14(n638), .DI13(n637), .DI12(n636), .DI11(n635), .DI10(n634), .DI9(n633), .DI8(n632), .DI7(n631),
 .DI6(n630), .DI5(n629), .DI4(n628), .DI3(n627), .DI2(n626), .DI1(n625), .DI0(n624), .WE(n621),
 .SYNC_IN(n1235), .SYNC_OUT(n1236));
// pragma CVASTRPROP INSTANCE "\depth_n.r_data " HDL_MEMORY_DECL "1 610 0 3 0"
MPR4X611 U1238 ( .A1(\depth_n.rptr [1]), .A0(\depth_n.rptr [0]), .SYNC_IN(n1236), .DO610(n4), .DO609(n5), .DO608(n6),
 .DO607(n7), .DO606(n8), .DO605(n9), .DO604(n10), .DO603(n11), .DO602(n12), .DO601(n13), .DO600(n14),
 .DO599(n15), .DO598(n16), .DO597(n17), .DO596(n18), .DO595(n19), .DO594(n20), .DO593(n21), .DO592(n22),
 .DO591(n23), .DO590(n24), .DO589(n25), .DO588(n26), .DO587(n27), .DO586(n28), .DO585(n29), .DO584(n30),
 .DO583(n31), .DO582(n32), .DO581(n33), .DO580(n34), .DO579(n35), .DO578(n36), .DO577(n37), .DO576(n38),
 .DO575(n39), .DO574(n40), .DO573(n41), .DO572(n42), .DO571(n43), .DO570(n44), .DO569(n45), .DO568(n46),
 .DO567(n47), .DO566(n48), .DO565(n49), .DO564(n50), .DO563(n51), .DO562(n52), .DO561(n53), .DO560(n54),
 .DO559(n55), .DO558(n56), .DO557(n57), .DO556(n58), .DO555(n59), .DO554(n60), .DO553(n61), .DO552(n62),
 .DO551(n63), .DO550(n64), .DO549(n65), .DO548(n66), .DO547(n67), .DO546(n68), .DO545(n69), .DO544(n70),
 .DO543(n71), .DO542(n72), .DO541(n73), .DO540(n74), .DO539(n75), .DO538(n76), .DO537(n77), .DO536(n78),
 .DO535(n79), .DO534(n80), .DO533(n81), .DO532(n82), .DO531(n83), .DO530(n84), .DO529(n85), .DO528(n86),
 .DO527(n87), .DO526(n88), .DO525(n89), .DO524(n90), .DO523(n91), .DO522(n92), .DO521(n93), .DO520(n94),
 .DO519(n95), .DO518(n96), .DO517(n97), .DO516(n98), .DO515(n99), .DO514(n100), .DO513(n101), .DO512(n102),
 .DO511(n103), .DO510(n104), .DO509(n105), .DO508(n106), .DO507(n107), .DO506(n108), .DO505(n109), .DO504(n110),
 .DO503(n111), .DO502(n112), .DO501(n113), .DO500(n114), .DO499(n115), .DO498(n116), .DO497(n117), .DO496(n118),
 .DO495(n119), .DO494(n120), .DO493(n121), .DO492(n122), .DO491(n123), .DO490(n124), .DO489(n125), .DO488(n126),
 .DO487(n127), .DO486(n128), .DO485(n129), .DO484(n130), .DO483(n131), .DO482(n132), .DO481(n133), .DO480(n134),
 .DO479(n135), .DO478(n136), .DO477(n137), .DO476(n138), .DO475(n139), .DO474(n140), .DO473(n141), .DO472(n142),
 .DO471(n143), .DO470(n144), .DO469(n145), .DO468(n146), .DO467(n147), .DO466(n148), .DO465(n149), .DO464(n150),
 .DO463(n151), .DO462(n152), .DO461(n153), .DO460(n154), .DO459(n155), .DO458(n156), .DO457(n157), .DO456(n158),
 .DO455(n159), .DO454(n160), .DO453(n161), .DO452(n162), .DO451(n163), .DO450(n164), .DO449(n165), .DO448(n166),
 .DO447(n167), .DO446(n168), .DO445(n169), .DO444(n170), .DO443(n171), .DO442(n172), .DO441(n173), .DO440(n174),
 .DO439(n175), .DO438(n176), .DO437(n177), .DO436(n178), .DO435(n179), .DO434(n180), .DO433(n181), .DO432(n182),
 .DO431(n183), .DO430(n184), .DO429(n185), .DO428(n186), .DO427(n187), .DO426(n188), .DO425(n189), .DO424(n190),
 .DO423(n191), .DO422(n192), .DO421(n193), .DO420(n194), .DO419(n195), .DO418(n196), .DO417(n197), .DO416(n198),
 .DO415(n199), .DO414(n200), .DO413(n201), .DO412(n202), .DO411(n203), .DO410(n204), .DO409(n205), .DO408(n206),
 .DO407(n207), .DO406(n208), .DO405(n209), .DO404(n210), .DO403(n211), .DO402(n212), .DO401(n213), .DO400(n214),
 .DO399(n215), .DO398(n216), .DO397(n217), .DO396(n218), .DO395(n219), .DO394(n220), .DO393(n221), .DO392(n222),
 .DO391(n223), .DO390(n224), .DO389(n225), .DO388(n226), .DO387(n227), .DO386(n228), .DO385(n229), .DO384(n230),
 .DO383(n231), .DO382(n232), .DO381(n233), .DO380(n234), .DO379(n235), .DO378(n236), .DO377(n237), .DO376(n238),
 .DO375(n239), .DO374(n240), .DO373(n241), .DO372(n242), .DO371(n243), .DO370(n244), .DO369(n245), .DO368(n246),
 .DO367(n247), .DO366(n248), .DO365(n249), .DO364(n250), .DO363(n251), .DO362(n252), .DO361(n253), .DO360(n254),
 .DO359(n255), .DO358(n256), .DO357(n257), .DO356(n258), .DO355(n259), .DO354(n260), .DO353(n261), .DO352(n262),
 .DO351(n263), .DO350(n264), .DO349(n265), .DO348(n266), .DO347(n267), .DO346(n268), .DO345(n269), .DO344(n270),
 .DO343(n271), .DO342(n272), .DO341(n273), .DO340(n274), .DO339(n275), .DO338(n276), .DO337(n277), .DO336(n278),
 .DO335(n279), .DO334(n280), .DO333(n281), .DO332(n282), .DO331(n283), .DO330(n284), .DO329(n285), .DO328(n286),
 .DO327(n287), .DO326(n288), .DO325(n289), .DO324(n290), .DO323(n291), .DO322(n292), .DO321(n293), .DO320(n294),
 .DO319(n295), .DO318(n296), .DO317(n297), .DO316(n298), .DO315(n299), .DO314(n300), .DO313(n301), .DO312(n302),
 .DO311(n303), .DO310(n304), .DO309(n305), .DO308(n306), .DO307(n307), .DO306(n308), .DO305(n309), .DO304(n310),
 .DO303(n311), .DO302(n312), .DO301(n313), .DO300(n314), .DO299(n315), .DO298(n316), .DO297(n317), .DO296(n318),
 .DO295(n319), .DO294(n320), .DO293(n321), .DO292(n322), .DO291(n323), .DO290(n324), .DO289(n325), .DO288(n326),
 .DO287(n327), .DO286(n328), .DO285(n329), .DO284(n330), .DO283(n331), .DO282(n332), .DO281(n333), .DO280(n334),
 .DO279(n335), .DO278(n336), .DO277(n337), .DO276(n338), .DO275(n339), .DO274(n340), .DO273(n341), .DO272(n342),
 .DO271(n343), .DO270(n344), .DO269(n345), .DO268(n346), .DO267(n347), .DO266(n348), .DO265(n349), .DO264(n350),
 .DO263(n351), .DO262(n352), .DO261(n353), .DO260(n354), .DO259(n355), .DO258(n356), .DO257(n357), .DO256(n358),
 .DO255(n359), .DO254(n360), .DO253(n361), .DO252(n362), .DO251(n363), .DO250(n364), .DO249(n365), .DO248(n366),
 .DO247(n367), .DO246(n368), .DO245(n369), .DO244(n370), .DO243(n371), .DO242(n372), .DO241(n373), .DO240(n374),
 .DO239(n375), .DO238(n376), .DO237(n377), .DO236(n378), .DO235(n379), .DO234(n380), .DO233(n381), .DO232(n382),
 .DO231(n383), .DO230(n384), .DO229(n385), .DO228(n386), .DO227(n387), .DO226(n388), .DO225(n389), .DO224(n390),
 .DO223(n391), .DO222(n392), .DO221(n393), .DO220(n394), .DO219(n395), .DO218(n396), .DO217(n397), .DO216(n398),
 .DO215(n399), .DO214(n400), .DO213(n401), .DO212(n402), .DO211(n403), .DO210(n404), .DO209(n405), .DO208(n406),
 .DO207(n407), .DO206(n408), .DO205(n409), .DO204(n410), .DO203(n411), .DO202(n412), .DO201(n413), .DO200(n414),
 .DO199(n415), .DO198(n416), .DO197(n417), .DO196(n418), .DO195(n419), .DO194(n420), .DO193(n421), .DO192(n422),
 .DO191(n423), .DO190(n424), .DO189(n425), .DO188(n426), .DO187(n427), .DO186(n428), .DO185(n429), .DO184(n430),
 .DO183(n431), .DO182(n432), .DO181(n433), .DO180(n434), .DO179(n435), .DO178(n436), .DO177(n437), .DO176(n438),
 .DO175(n439), .DO174(n440), .DO173(n441), .DO172(n442), .DO171(n443), .DO170(n444), .DO169(n445), .DO168(n446),
 .DO167(n447), .DO166(n448), .DO165(n449), .DO164(n450), .DO163(n451), .DO162(n452), .DO161(n453), .DO160(n454),
 .DO159(n455), .DO158(n456), .DO157(n457), .DO156(n458), .DO155(n459), .DO154(n460), .DO153(n461), .DO152(n462),
 .DO151(n463), .DO150(n464), .DO149(n465), .DO148(n466), .DO147(n467), .DO146(n468), .DO145(n469), .DO144(n470),
 .DO143(n471), .DO142(n472), .DO141(n473), .DO140(n474), .DO139(n475), .DO138(n476), .DO137(n477), .DO136(n478),
 .DO135(n479), .DO134(n480), .DO133(n481), .DO132(n482), .DO131(n483), .DO130(n484), .DO129(n485), .DO128(n486),
 .DO127(n487), .DO126(n488), .DO125(n489), .DO124(n490), .DO123(n491), .DO122(n492), .DO121(n493), .DO120(n494),
 .DO119(n495), .DO118(n496), .DO117(n497), .DO116(n498), .DO115(n499), .DO114(n500), .DO113(n501), .DO112(n502),
 .DO111(n503), .DO110(n504), .DO109(n505), .DO108(n506), .DO107(n507), .DO106(n508), .DO105(n509), .DO104(n510),
 .DO103(n511), .DO102(n512), .DO101(n513), .DO100(n514), .DO99(n515), .DO98(n516), .DO97(n517), .DO96(n518),
 .DO95(n519), .DO94(n520), .DO93(n521), .DO92(n522), .DO91(n523), .DO90(n524), .DO89(n525), .DO88(n526),
 .DO87(n527), .DO86(n528), .DO85(n529), .DO84(n530), .DO83(n531), .DO82(n532), .DO81(n533), .DO80(n534),
 .DO79(n535), .DO78(n536), .DO77(n537), .DO76(n538), .DO75(n539), .DO74(n540), .DO73(n541), .DO72(n542),
 .DO71(n543), .DO70(n544), .DO69(n545), .DO68(n546), .DO67(n547), .DO66(n548), .DO65(n549), .DO64(n550),
 .DO63(n551), .DO62(n552), .DO61(n553), .DO60(n554), .DO59(n555), .DO58(n556), .DO57(n557), .DO56(n558),
 .DO55(n559), .DO54(n560), .DO53(n561), .DO52(n562), .DO51(n563), .DO50(n564), .DO49(n565), .DO48(n566),
 .DO47(n567), .DO46(n568), .DO45(n569), .DO44(n570), .DO43(n571), .DO42(n572), .DO41(n573), .DO40(n574),
 .DO39(n575), .DO38(n576), .DO37(n577), .DO36(n578), .DO35(n579), .DO34(n580), .DO33(n581), .DO32(n582),
 .DO31(n583), .DO30(n584), .DO29(n585), .DO28(n586), .DO27(n587), .DO26(n588), .DO25(n589), .DO24(n590),
 .DO23(n591), .DO22(n592), .DO21(n593), .DO20(n594), .DO19(n595), .DO18(n596), .DO17(n597), .DO16(n598),
 .DO15(n599), .DO14(n600), .DO13(n601), .DO12(n602), .DO11(n603), .DO10(n604), .DO9(n605), .DO8(n606),
 .DO7(n607), .DO6(n608), .DO5(n609), .DO4(n610), .DO3(n611), .DO2(n612), .DO1(n613), .DO0(n614),
 .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "0 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 depth_n  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n.genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n"
endmodule
`ifdef CBV
`else
`ifdef MPW4X611_MPR4X611
`else
module MPW4X611( A1, A0, DI610, DI609, DI608, DI607, DI606,
 DI605, DI604, DI603, DI602, DI601, DI600, DI599, DI598,
 DI597, DI596, DI595, DI594, DI593, DI592, DI591, DI590,
 DI589, DI588, DI587, DI586, DI585, DI584, DI583, DI582,
 DI581, DI580, DI579, DI578, DI577, DI576, DI575, DI574,
 DI573, DI572, DI571, DI570, DI569, DI568, DI567, DI566,
 DI565, DI564, DI563, DI562, DI561, DI560, DI559, DI558,
 DI557, DI556, DI555, DI554, DI553, DI552, DI551, DI550,
 DI549, DI548, DI547, DI546, DI545, DI544, DI543, DI542,
 DI541, DI540, DI539, DI538, DI537, DI536, DI535, DI534,
 DI533, DI532, DI531, DI530, DI529, DI528, DI527, DI526,
 DI525, DI524, DI523, DI522, DI521, DI520, DI519, DI518,
 DI517, DI516, DI515, DI514, DI513, DI512, DI511, DI510,
 DI509, DI508, DI507, DI506, DI505, DI504, DI503, DI502,
 DI501, DI500, DI499, DI498, DI497, DI496, DI495, DI494,
 DI493, DI492, DI491, DI490, DI489, DI488, DI487, DI486,
 DI485, DI484, DI483, DI482, DI481, DI480, DI479, DI478,
 DI477, DI476, DI475, DI474, DI473, DI472, DI471, DI470,
 DI469, DI468, DI467, DI466, DI465, DI464, DI463, DI462,
 DI461, DI460, DI459, DI458, DI457, DI456, DI455, DI454,
 DI453, DI452, DI451, DI450, DI449, DI448, DI447, DI446,
 DI445, DI444, DI443, DI442, DI441, DI440, DI439, DI438,
 DI437, DI436, DI435, DI434, DI433, DI432, DI431, DI430,
 DI429, DI428, DI427, DI426, DI425, DI424, DI423, DI422,
 DI421, DI420, DI419, DI418, DI417, DI416, DI415, DI414,
 DI413, DI412, DI411, DI410, DI409, DI408, DI407, DI406,
 DI405, DI404, DI403, DI402, DI401, DI400, DI399, DI398,
 DI397, DI396, DI395, DI394, DI393, DI392, DI391, DI390,
 DI389, DI388, DI387, DI386, DI385, DI384, DI383, DI382,
 DI381, DI380, DI379, DI378, DI377, DI376, DI375, DI374,
 DI373, DI372, DI371, DI370, DI369, DI368, DI367, DI366,
 DI365, DI364, DI363, DI362, DI361, DI360, DI359, DI358,
 DI357, DI356, DI355, DI354, DI353, DI352, DI351, DI350,
 DI349, DI348, DI347, DI346, DI345, DI344, DI343, DI342,
 DI341, DI340, DI339, DI338, DI337, DI336, DI335, DI334,
 DI333, DI332, DI331, DI330, DI329, DI328, DI327, DI326,
 DI325, DI324, DI323, DI322, DI321, DI320, DI319, DI318,
 DI317, DI316, DI315, DI314, DI313, DI312, DI311, DI310,
 DI309, DI308, DI307, DI306, DI305, DI304, DI303, DI302,
 DI301, DI300, DI299, DI298, DI297, DI296, DI295, DI294,
 DI293, DI292, DI291, DI290, DI289, DI288, DI287, DI286,
 DI285, DI284, DI283, DI282, DI281, DI280, DI279, DI278,
 DI277, DI276, DI275, DI274, DI273, DI272, DI271, DI270,
 DI269, DI268, DI267, DI266, DI265, DI264, DI263, DI262,
 DI261, DI260, DI259, DI258, DI257, DI256, DI255, DI254,
 DI253, DI252, DI251, DI250, DI249, DI248, DI247, DI246,
 DI245, DI244, DI243, DI242, DI241, DI240, DI239, DI238,
 DI237, DI236, DI235, DI234, DI233, DI232, DI231, DI230,
 DI229, DI228, DI227, DI226, DI225, DI224, DI223, DI222,
 DI221, DI220, DI219, DI218, DI217, DI216, DI215, DI214,
 DI213, DI212, DI211, DI210, DI209, DI208, DI207, DI206,
 DI205, DI204, DI203, DI202, DI201, DI200, DI199, DI198,
 DI197, DI196, DI195, DI194, DI193, DI192, DI191, DI190,
 DI189, DI188, DI187, DI186, DI185, DI184, DI183, DI182,
 DI181, DI180, DI179, DI178, DI177, DI176, DI175, DI174,
 DI173, DI172, DI171, DI170, DI169, DI168, DI167, DI166,
 DI165, DI164, DI163, DI162, DI161, DI160, DI159, DI158,
 DI157, DI156, DI155, DI154, DI153, DI152, DI151, DI150,
 DI149, DI148, DI147, DI146, DI145, DI144, DI143, DI142,
 DI141, DI140, DI139, DI138, DI137, DI136, DI135, DI134,
 DI133, DI132, DI131, DI130, DI129, DI128, DI127, DI126,
 DI125, DI124, DI123, DI122, DI121, DI120, DI119, DI118,
 DI117, DI116, DI115, DI114, DI113, DI112, DI111, DI110,
 DI109, DI108, DI107, DI106, DI105, DI104, DI103, DI102,
 DI101, DI100, DI99, DI98, DI97, DI96, DI95, DI94,
 DI93, DI92, DI91, DI90, DI89, DI88, DI87, DI86,
 DI85, DI84, DI83, DI82, DI81, DI80, DI79, DI78,
 DI77, DI76, DI75, DI74, DI73, DI72, DI71, DI70,
 DI69, DI68, DI67, DI66, DI65, DI64, DI63, DI62,
 DI61, DI60, DI59, DI58, DI57, DI56, DI55, DI54,
 DI53, DI52, DI51, DI50, DI49, DI48, DI47, DI46,
 DI45, DI44, DI43, DI42, DI41, DI40, DI39, DI38,
 DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30,
 DI29, DI28, DI27, DI26, DI25, DI24, DI23, DI22,
 DI21, DI20, DI19, DI18, DI17, DI16, DI15, DI14,
 DI13, DI12, DI11, DI10, DI9, DI8, DI7, DI6,
 DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN,
 SYNC_OUT);
input  A1, A0, DI610, DI609, DI608, DI607, DI606, DI605,
 DI604, DI603, DI602, DI601, DI600, DI599, DI598, DI597, DI596, DI595,
 DI594, DI593, DI592, DI591, DI590, DI589, DI588, DI587, DI586, DI585,
 DI584, DI583, DI582, DI581, DI580, DI579, DI578, DI577, DI576, DI575,
 DI574, DI573, DI572, DI571, DI570, DI569, DI568, DI567, DI566, DI565,
 DI564, DI563, DI562, DI561, DI560, DI559, DI558, DI557, DI556, DI555,
 DI554, DI553, DI552, DI551, DI550, DI549, DI548, DI547, DI546, DI545,
 DI544, DI543, DI542, DI541, DI540, DI539, DI538, DI537, DI536, DI535,
 DI534, DI533, DI532, DI531, DI530, DI529, DI528, DI527, DI526, DI525,
 DI524, DI523, DI522, DI521, DI520, DI519, DI518, DI517, DI516, DI515,
 DI514, DI513, DI512, DI511, DI510, DI509, DI508, DI507, DI506, DI505,
 DI504, DI503, DI502, DI501, DI500, DI499, DI498, DI497, DI496, DI495,
 DI494, DI493, DI492, DI491, DI490, DI489, DI488, DI487, DI486, DI485,
 DI484, DI483, DI482, DI481, DI480, DI479, DI478, DI477, DI476, DI475,
 DI474, DI473, DI472, DI471, DI470, DI469, DI468, DI467, DI466, DI465,
 DI464, DI463, DI462, DI461, DI460, DI459, DI458, DI457, DI456, DI455,
 DI454, DI453, DI452, DI451, DI450, DI449, DI448, DI447, DI446, DI445,
 DI444, DI443, DI442, DI441, DI440, DI439, DI438, DI437, DI436, DI435,
 DI434, DI433, DI432, DI431, DI430, DI429, DI428, DI427, DI426, DI425,
 DI424, DI423, DI422, DI421, DI420, DI419, DI418, DI417, DI416, DI415,
 DI414, DI413, DI412, DI411, DI410, DI409, DI408, DI407, DI406, DI405,
 DI404, DI403, DI402, DI401, DI400, DI399, DI398, DI397, DI396, DI395,
 DI394, DI393, DI392, DI391, DI390, DI389, DI388, DI387, DI386, DI385,
 DI384, DI383, DI382, DI381, DI380, DI379, DI378, DI377, DI376, DI375,
 DI374, DI373, DI372, DI371, DI370, DI369, DI368, DI367, DI366, DI365,
 DI364, DI363, DI362, DI361, DI360, DI359, DI358, DI357, DI356, DI355,
 DI354, DI353, DI352, DI351, DI350, DI349, DI348, DI347, DI346, DI345,
 DI344, DI343, DI342, DI341, DI340, DI339, DI338, DI337, DI336, DI335,
 DI334, DI333, DI332, DI331, DI330, DI329, DI328, DI327, DI326, DI325,
 DI324, DI323, DI322, DI321, DI320, DI319, DI318, DI317, DI316, DI315,
 DI314, DI313, DI312, DI311, DI310, DI309, DI308, DI307, DI306, DI305,
 DI304, DI303, DI302, DI301, DI300, DI299, DI298, DI297, DI296, DI295,
 DI294, DI293, DI292, DI291, DI290, DI289, DI288, DI287, DI286, DI285,
 DI284, DI283, DI282, DI281, DI280, DI279, DI278, DI277, DI276, DI275,
 DI274, DI273, DI272, DI271, DI270, DI269, DI268, DI267, DI266, DI265,
 DI264, DI263, DI262, DI261, DI260, DI259, DI258, DI257, DI256, DI255,
 DI254, DI253, DI252, DI251, DI250, DI249, DI248, DI247, DI246, DI245,
 DI244, DI243, DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235,
 DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227, DI226, DI225,
 DI224, DI223, DI222, DI221, DI220, DI219, DI218, DI217, DI216, DI215,
 DI214, DI213, DI212, DI211, DI210, DI209, DI208, DI207, DI206, DI205,
 DI204, DI203, DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195,
 DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187, DI186, DI185,
 DI184, DI183, DI182, DI181, DI180, DI179, DI178, DI177, DI176, DI175,
 DI174, DI173, DI172, DI171, DI170, DI169, DI168, DI167, DI166, DI165,
 DI164, DI163, DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155,
 DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147, DI146, DI145,
 DI144, DI143, DI142, DI141, DI140, DI139, DI138, DI137, DI136, DI135,
 DI134, DI133, DI132, DI131, DI130, DI129, DI128, DI127, DI126, DI125,
 DI124, DI123, DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115,
 DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107, DI106, DI105,
 DI104, DI103, DI102, DI101, DI100, DI99, DI98, DI97, DI96, DI95,
 DI94, DI93, DI92, DI91, DI90, DI89, DI88, DI87, DI86, DI85,
 DI84, DI83, DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75,
 DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67, DI66, DI65,
 DI64, DI63, DI62, DI61, DI60, DI59, DI58, DI57, DI56, DI55,
 DI54, DI53, DI52, DI51, DI50, DI49, DI48, DI47, DI46, DI45,
 DI44, DI43, DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35,
 DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26, DI25,
 DI24, DI23, DI22, DI21, DI20, DI19, DI18, DI17, DI16, DI15,
 DI14, DI13, DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5,
 DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR4X611_
`else
module MPR4X611( A1, A0, SYNC_IN, DO610, DO609, DO608, DO607,
 DO606, DO605, DO604, DO603, DO602, DO601, DO600, DO599,
 DO598, DO597, DO596, DO595, DO594, DO593, DO592, DO591,
 DO590, DO589, DO588, DO587, DO586, DO585, DO584, DO583,
 DO582, DO581, DO580, DO579, DO578, DO577, DO576, DO575,
 DO574, DO573, DO572, DO571, DO570, DO569, DO568, DO567,
 DO566, DO565, DO564, DO563, DO562, DO561, DO560, DO559,
 DO558, DO557, DO556, DO555, DO554, DO553, DO552, DO551,
 DO550, DO549, DO548, DO547, DO546, DO545, DO544, DO543,
 DO542, DO541, DO540, DO539, DO538, DO537, DO536, DO535,
 DO534, DO533, DO532, DO531, DO530, DO529, DO528, DO527,
 DO526, DO525, DO524, DO523, DO522, DO521, DO520, DO519,
 DO518, DO517, DO516, DO515, DO514, DO513, DO512, DO511,
 DO510, DO509, DO508, DO507, DO506, DO505, DO504, DO503,
 DO502, DO501, DO500, DO499, DO498, DO497, DO496, DO495,
 DO494, DO493, DO492, DO491, DO490, DO489, DO488, DO487,
 DO486, DO485, DO484, DO483, DO482, DO481, DO480, DO479,
 DO478, DO477, DO476, DO475, DO474, DO473, DO472, DO471,
 DO470, DO469, DO468, DO467, DO466, DO465, DO464, DO463,
 DO462, DO461, DO460, DO459, DO458, DO457, DO456, DO455,
 DO454, DO453, DO452, DO451, DO450, DO449, DO448, DO447,
 DO446, DO445, DO444, DO443, DO442, DO441, DO440, DO439,
 DO438, DO437, DO436, DO435, DO434, DO433, DO432, DO431,
 DO430, DO429, DO428, DO427, DO426, DO425, DO424, DO423,
 DO422, DO421, DO420, DO419, DO418, DO417, DO416, DO415,
 DO414, DO413, DO412, DO411, DO410, DO409, DO408, DO407,
 DO406, DO405, DO404, DO403, DO402, DO401, DO400, DO399,
 DO398, DO397, DO396, DO395, DO394, DO393, DO392, DO391,
 DO390, DO389, DO388, DO387, DO386, DO385, DO384, DO383,
 DO382, DO381, DO380, DO379, DO378, DO377, DO376, DO375,
 DO374, DO373, DO372, DO371, DO370, DO369, DO368, DO367,
 DO366, DO365, DO364, DO363, DO362, DO361, DO360, DO359,
 DO358, DO357, DO356, DO355, DO354, DO353, DO352, DO351,
 DO350, DO349, DO348, DO347, DO346, DO345, DO344, DO343,
 DO342, DO341, DO340, DO339, DO338, DO337, DO336, DO335,
 DO334, DO333, DO332, DO331, DO330, DO329, DO328, DO327,
 DO326, DO325, DO324, DO323, DO322, DO321, DO320, DO319,
 DO318, DO317, DO316, DO315, DO314, DO313, DO312, DO311,
 DO310, DO309, DO308, DO307, DO306, DO305, DO304, DO303,
 DO302, DO301, DO300, DO299, DO298, DO297, DO296, DO295,
 DO294, DO293, DO292, DO291, DO290, DO289, DO288, DO287,
 DO286, DO285, DO284, DO283, DO282, DO281, DO280, DO279,
 DO278, DO277, DO276, DO275, DO274, DO273, DO272, DO271,
 DO270, DO269, DO268, DO267, DO266, DO265, DO264, DO263,
 DO262, DO261, DO260, DO259, DO258, DO257, DO256, DO255,
 DO254, DO253, DO252, DO251, DO250, DO249, DO248, DO247,
 DO246, DO245, DO244, DO243, DO242, DO241, DO240, DO239,
 DO238, DO237, DO236, DO235, DO234, DO233, DO232, DO231,
 DO230, DO229, DO228, DO227, DO226, DO225, DO224, DO223,
 DO222, DO221, DO220, DO219, DO218, DO217, DO216, DO215,
 DO214, DO213, DO212, DO211, DO210, DO209, DO208, DO207,
 DO206, DO205, DO204, DO203, DO202, DO201, DO200, DO199,
 DO198, DO197, DO196, DO195, DO194, DO193, DO192, DO191,
 DO190, DO189, DO188, DO187, DO186, DO185, DO184, DO183,
 DO182, DO181, DO180, DO179, DO178, DO177, DO176, DO175,
 DO174, DO173, DO172, DO171, DO170, DO169, DO168, DO167,
 DO166, DO165, DO164, DO163, DO162, DO161, DO160, DO159,
 DO158, DO157, DO156, DO155, DO154, DO153, DO152, DO151,
 DO150, DO149, DO148, DO147, DO146, DO145, DO144, DO143,
 DO142, DO141, DO140, DO139, DO138, DO137, DO136, DO135,
 DO134, DO133, DO132, DO131, DO130, DO129, DO128, DO127,
 DO126, DO125, DO124, DO123, DO122, DO121, DO120, DO119,
 DO118, DO117, DO116, DO115, DO114, DO113, DO112, DO111,
 DO110, DO109, DO108, DO107, DO106, DO105, DO104, DO103,
 DO102, DO101, DO100, DO99, DO98, DO97, DO96, DO95,
 DO94, DO93, DO92, DO91, DO90, DO89, DO88, DO87,
 DO86, DO85, DO84, DO83, DO82, DO81, DO80, DO79,
 DO78, DO77, DO76, DO75, DO74, DO73, DO72, DO71,
 DO70, DO69, DO68, DO67, DO66, DO65, DO64, DO63,
 DO62, DO61, DO60, DO59, DO58, DO57, DO56, DO55,
 DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47,
 DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39,
 DO38, DO37, DO36, DO35, DO34, DO33, DO32, DO31,
 DO30, DO29, DO28, DO27, DO26, DO25, DO24, DO23,
 DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15,
 DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7,
 DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT);
input  A1, A0, SYNC_IN;
output  DO610, DO609, DO608, DO607, DO606, DO605, DO604, DO603,
 DO602, DO601, DO600, DO599, DO598, DO597, DO596, DO595, DO594, DO593,
 DO592, DO591, DO590, DO589, DO588, DO587, DO586, DO585, DO584, DO583,
 DO582, DO581, DO580, DO579, DO578, DO577, DO576, DO575, DO574, DO573,
 DO572, DO571, DO570, DO569, DO568, DO567, DO566, DO565, DO564, DO563,
 DO562, DO561, DO560, DO559, DO558, DO557, DO556, DO555, DO554, DO553,
 DO552, DO551, DO550, DO549, DO548, DO547, DO546, DO545, DO544, DO543,
 DO542, DO541, DO540, DO539, DO538, DO537, DO536, DO535, DO534, DO533,
 DO532, DO531, DO530, DO529, DO528, DO527, DO526, DO525, DO524, DO523,
 DO522, DO521, DO520, DO519, DO518, DO517, DO516, DO515, DO514, DO513,
 DO512, DO511, DO510, DO509, DO508, DO507, DO506, DO505, DO504, DO503,
 DO502, DO501, DO500, DO499, DO498, DO497, DO496, DO495, DO494, DO493,
 DO492, DO491, DO490, DO489, DO488, DO487, DO486, DO485, DO484, DO483,
 DO482, DO481, DO480, DO479, DO478, DO477, DO476, DO475, DO474, DO473,
 DO472, DO471, DO470, DO469, DO468, DO467, DO466, DO465, DO464, DO463,
 DO462, DO461, DO460, DO459, DO458, DO457, DO456, DO455, DO454, DO453,
 DO452, DO451, DO450, DO449, DO448, DO447, DO446, DO445, DO444, DO443,
 DO442, DO441, DO440, DO439, DO438, DO437, DO436, DO435, DO434, DO433,
 DO432, DO431, DO430, DO429, DO428, DO427, DO426, DO425, DO424, DO423,
 DO422, DO421, DO420, DO419, DO418, DO417, DO416, DO415, DO414, DO413,
 DO412, DO411, DO410, DO409, DO408, DO407, DO406, DO405, DO404, DO403,
 DO402, DO401, DO400, DO399, DO398, DO397, DO396, DO395, DO394, DO393,
 DO392, DO391, DO390, DO389, DO388, DO387, DO386, DO385, DO384, DO383,
 DO382, DO381, DO380, DO379, DO378, DO377, DO376, DO375, DO374, DO373,
 DO372, DO371, DO370, DO369, DO368, DO367, DO366, DO365, DO364, DO363,
 DO362, DO361, DO360, DO359, DO358, DO357, DO356, DO355, DO354, DO353,
 DO352, DO351, DO350, DO349, DO348, DO347, DO346, DO345, DO344, DO343,
 DO342, DO341, DO340, DO339, DO338, DO337, DO336, DO335, DO334, DO333,
 DO332, DO331, DO330, DO329, DO328, DO327, DO326, DO325, DO324, DO323,
 DO322, DO321, DO320, DO319, DO318, DO317, DO316, DO315, DO314, DO313,
 DO312, DO311, DO310, DO309, DO308, DO307, DO306, DO305, DO304, DO303,
 DO302, DO301, DO300, DO299, DO298, DO297, DO296, DO295, DO294, DO293,
 DO292, DO291, DO290, DO289, DO288, DO287, DO286, DO285, DO284, DO283,
 DO282, DO281, DO280, DO279, DO278, DO277, DO276, DO275, DO274, DO273,
 DO272, DO271, DO270, DO269, DO268, DO267, DO266, DO265, DO264, DO263,
 DO262, DO261, DO260, DO259, DO258, DO257, DO256, DO255, DO254, DO253,
 DO252, DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244, DO243,
 DO242, DO241, DO240, DO239, DO238, DO237, DO236, DO235, DO234, DO233,
 DO232, DO231, DO230, DO229, DO228, DO227, DO226, DO225, DO224, DO223,
 DO222, DO221, DO220, DO219, DO218, DO217, DO216, DO215, DO214, DO213,
 DO212, DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204, DO203,
 DO202, DO201, DO200, DO199, DO198, DO197, DO196, DO195, DO194, DO193,
 DO192, DO191, DO190, DO189, DO188, DO187, DO186, DO185, DO184, DO183,
 DO182, DO181, DO180, DO179, DO178, DO177, DO176, DO175, DO174, DO173,
 DO172, DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164, DO163,
 DO162, DO161, DO160, DO159, DO158, DO157, DO156, DO155, DO154, DO153,
 DO152, DO151, DO150, DO149, DO148, DO147, DO146, DO145, DO144, DO143,
 DO142, DO141, DO140, DO139, DO138, DO137, DO136, DO135, DO134, DO133,
 DO132, DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124, DO123,
 DO122, DO121, DO120, DO119, DO118, DO117, DO116, DO115, DO114, DO113,
 DO112, DO111, DO110, DO109, DO108, DO107, DO106, DO105, DO104, DO103,
 DO102, DO101, DO100, DO99, DO98, DO97, DO96, DO95, DO94, DO93,
 DO92, DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84, DO83,
 DO82, DO81, DO80, DO79, DO78, DO77, DO76, DO75, DO74, DO73,
 DO72, DO71, DO70, DO69, DO68, DO67, DO66, DO65, DO64, DO63,
 DO62, DO61, DO60, DO59, DO58, DO57, DO56, DO55, DO54, DO53,
 DO52, DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44, DO43,
 DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35, DO34, DO33,
 DO32, DO31, DO30, DO29, DO28, DO27, DO26, DO25, DO24, DO23,
 DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14, DO13,
 DO12, DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4, DO3,
 DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR4X611_
`endif
`define MPW4X611_MPR4X611
`endif
`endif
