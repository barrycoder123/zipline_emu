
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_gfifo_port_1_2 ( tkout, tkin, ireq, cbid, len, idata, CGFtsReq, 
	CGFcbid, CGFlen, CGFidata, CGFfull, CLBreq, CLBrd, CLBwr, CLBfull, 
	Rtkin);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output tkout;
input tkin;
input ireq;
input [19:0] cbid;
input [11:0] len;
input [0:0] idata;
output CGFtsReq;
output [19:0] CGFcbid;
output [11:0] CGFlen;
output [511:0] CGFidata;
input CGFfull;
output CLBreq;
input [3:0] CLBrd;
input [3:0] CLBwr;
input CLBfull;
input Rtkin;
wire fclk;
wire enq;
wire CLBreqWhileFull;
`_2_ wire en;
`_2_ wire ack;
`_2_ wire [0:0] odata;
`_2_ wire oreq;
`_2_ wire [19:0] ocbid;
`_2_ wire [19:0] xcbid;
`_2_ wire [11:0] olen;
`_2_ wire [11:0] xlen;
`_2_ wire [0:0] sel;
`_2_ wire [0:0] xdata;
wire [31:0] i;
`_2_ wire ireqR;
supply1 n5;
Q_ASSIGN U0 ( .B(len[0]), .A(xlen[0]));
Q_ASSIGN U1 ( .B(len[0]), .A(olen[0]));
Q_ASSIGN U2 ( .B(len[1]), .A(xlen[1]));
Q_ASSIGN U3 ( .B(len[1]), .A(olen[1]));
Q_ASSIGN U4 ( .B(len[2]), .A(xlen[2]));
Q_ASSIGN U5 ( .B(len[2]), .A(olen[2]));
Q_ASSIGN U6 ( .B(len[3]), .A(xlen[3]));
Q_ASSIGN U7 ( .B(len[3]), .A(olen[3]));
Q_ASSIGN U8 ( .B(len[4]), .A(xlen[4]));
Q_ASSIGN U9 ( .B(len[4]), .A(olen[4]));
Q_ASSIGN U10 ( .B(len[5]), .A(xlen[5]));
Q_ASSIGN U11 ( .B(len[5]), .A(olen[5]));
Q_ASSIGN U12 ( .B(len[6]), .A(xlen[6]));
Q_ASSIGN U13 ( .B(len[6]), .A(olen[6]));
Q_ASSIGN U14 ( .B(len[7]), .A(xlen[7]));
Q_ASSIGN U15 ( .B(len[7]), .A(olen[7]));
Q_ASSIGN U16 ( .B(len[8]), .A(xlen[8]));
Q_ASSIGN U17 ( .B(len[8]), .A(olen[8]));
Q_ASSIGN U18 ( .B(len[9]), .A(xlen[9]));
Q_ASSIGN U19 ( .B(len[9]), .A(olen[9]));
Q_ASSIGN U20 ( .B(len[10]), .A(xlen[10]));
Q_ASSIGN U21 ( .B(len[10]), .A(olen[10]));
Q_ASSIGN U22 ( .B(len[11]), .A(xlen[11]));
Q_ASSIGN U23 ( .B(len[11]), .A(olen[11]));
Q_BUF U24 ( .A(ocbid[0]), .Z(xcbid[0]));
Q_BUF U25 ( .A(ocbid[1]), .Z(xcbid[1]));
Q_BUF U26 ( .A(ocbid[2]), .Z(xcbid[2]));
Q_BUF U27 ( .A(ocbid[3]), .Z(xcbid[3]));
Q_BUF U28 ( .A(ocbid[4]), .Z(xcbid[4]));
Q_BUF U29 ( .A(ocbid[5]), .Z(xcbid[5]));
Q_BUF U30 ( .A(ocbid[6]), .Z(xcbid[6]));
Q_BUF U31 ( .A(ocbid[7]), .Z(xcbid[7]));
Q_BUF U32 ( .A(ocbid[8]), .Z(xcbid[8]));
Q_BUF U33 ( .A(ocbid[9]), .Z(xcbid[9]));
Q_BUF U34 ( .A(ocbid[10]), .Z(xcbid[10]));
Q_BUF U35 ( .A(ocbid[11]), .Z(xcbid[11]));
Q_BUF U36 ( .A(ocbid[12]), .Z(xcbid[12]));
Q_BUF U37 ( .A(ocbid[13]), .Z(xcbid[13]));
Q_BUF U38 ( .A(ocbid[14]), .Z(xcbid[14]));
Q_BUF U39 ( .A(ocbid[15]), .Z(xcbid[15]));
Q_BUF U40 ( .A(ocbid[16]), .Z(xcbid[16]));
Q_BUF U41 ( .A(ocbid[17]), .Z(xcbid[17]));
Q_BUF U42 ( .A(ocbid[18]), .Z(xcbid[18]));
Q_BUF U43 ( .A(ocbid[19]), .Z(xcbid[19]));
Q_BUF U44 ( .A(odata[0]), .Z(xdata[0]));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_EV_WOR_START qi ( .A(CLBreqWhileFull));
Q_INV U47 ( .A(n4), .Z(tkout));
Q_XNR2 U48 ( .A0(oreq), .A1(ack), .Z(n4));
Q_CCLKCHK cchk ( .sig(ireq));
Q_AN02 U50 ( .A0(enq), .A1(CLBfull), .Z(CLBreqWhileFull));
Q_AN02 U51 ( .A0(n2), .A1(n3), .Z(enq));
Q_INV U52 ( .A(xc_top.GFLock2), .Z(n3));
Q_XOR2 U53 ( .A0(ireq), .A1(ireqR), .Z(n2));
Q_BUFZP U54 ( .OE(CLBreqWhileFull), .A(n5), .Z(xc_top.GFLBfull));
Q_BUFZP U55 ( .OE(en), .A(xcbid[0]), .Z(CGFcbid[0]));
Q_BUFZP U56 ( .OE(en), .A(xcbid[1]), .Z(CGFcbid[1]));
Q_BUFZP U57 ( .OE(en), .A(xcbid[2]), .Z(CGFcbid[2]));
Q_BUFZP U58 ( .OE(en), .A(xcbid[3]), .Z(CGFcbid[3]));
Q_BUFZP U59 ( .OE(en), .A(xcbid[4]), .Z(CGFcbid[4]));
Q_BUFZP U60 ( .OE(en), .A(xcbid[5]), .Z(CGFcbid[5]));
Q_BUFZP U61 ( .OE(en), .A(xcbid[6]), .Z(CGFcbid[6]));
Q_BUFZP U62 ( .OE(en), .A(xcbid[7]), .Z(CGFcbid[7]));
Q_BUFZP U63 ( .OE(en), .A(xcbid[8]), .Z(CGFcbid[8]));
Q_BUFZP U64 ( .OE(en), .A(xcbid[9]), .Z(CGFcbid[9]));
Q_BUFZP U65 ( .OE(en), .A(xcbid[10]), .Z(CGFcbid[10]));
Q_BUFZP U66 ( .OE(en), .A(xcbid[11]), .Z(CGFcbid[11]));
Q_BUFZP U67 ( .OE(en), .A(xcbid[12]), .Z(CGFcbid[12]));
Q_BUFZP U68 ( .OE(en), .A(xcbid[13]), .Z(CGFcbid[13]));
Q_BUFZP U69 ( .OE(en), .A(xcbid[14]), .Z(CGFcbid[14]));
Q_BUFZP U70 ( .OE(en), .A(xcbid[15]), .Z(CGFcbid[15]));
Q_BUFZP U71 ( .OE(en), .A(xcbid[16]), .Z(CGFcbid[16]));
Q_BUFZP U72 ( .OE(en), .A(xcbid[17]), .Z(CGFcbid[17]));
Q_BUFZP U73 ( .OE(en), .A(xcbid[18]), .Z(CGFcbid[18]));
Q_BUFZP U74 ( .OE(en), .A(xcbid[19]), .Z(CGFcbid[19]));
Q_BUFZP U75 ( .OE(en), .A(len[0]), .Z(CGFlen[0]));
Q_BUFZP U76 ( .OE(en), .A(len[1]), .Z(CGFlen[1]));
Q_BUFZP U77 ( .OE(en), .A(len[2]), .Z(CGFlen[2]));
Q_BUFZP U78 ( .OE(en), .A(len[3]), .Z(CGFlen[3]));
Q_BUFZP U79 ( .OE(en), .A(len[4]), .Z(CGFlen[4]));
Q_BUFZP U80 ( .OE(en), .A(len[5]), .Z(CGFlen[5]));
Q_BUFZP U81 ( .OE(en), .A(len[6]), .Z(CGFlen[6]));
Q_BUFZP U82 ( .OE(en), .A(len[7]), .Z(CGFlen[7]));
Q_BUFZP U83 ( .OE(en), .A(len[8]), .Z(CGFlen[8]));
Q_BUFZP U84 ( .OE(en), .A(len[9]), .Z(CGFlen[9]));
Q_BUFZP U85 ( .OE(en), .A(len[10]), .Z(CGFlen[10]));
Q_BUFZP U86 ( .OE(en), .A(len[11]), .Z(CGFlen[11]));
Q_BUFZP U87 ( .OE(en), .A(xdata[0]), .Z(CGFidata[0]));
Q_BUFZP U88 ( .OE(enq), .A(n5), .Z(CLBreq));
Q_BUFZP U89 ( .OE(enq), .A(n5), .Z(CGFtsReq));
Q_INV U90 ( .A(CLBwr[2]), .Z(n6));
ixc_bind \genblk3.b5 ( CLBfull, IXC_GFIFO.O.O.LBfull);
ixc_bind_4 \genblk3.b4 ( CLBwr[3:0], IXC_GFIFO.O.O.LBwr[3:0]);
ixc_bind_4 \genblk3.b3 ( CLBrd[3:0], IXC_GFIFO.O.O.LBrd[3:0]);
ixc_bind \genblk3.b2 ( CLBreq, IXC_GFIFO.O.O.LBreq);
ixc_bind \genblk3.b1 ( CGFfull, IXC_GFIFO.O.O.GFfull);
ixc_bind \genblk3.b0 ( CGFtsReq, IXC_GFIFO.O.O.GFtsReq);
Q_MX02 U97 ( .S(xc_top.GFLock2), .A0(oreq), .A1(ireq), .Z(n8));
Q_FDP0UA U98 ( .D(n9), .QTFCLK( ), .Q(ack));
Q_MX02 U99 ( .S(n14), .A0(ack), .A1(n8), .Z(n9));
Q_FDP0UA U100 ( .D(n10), .QTFCLK( ), .Q(en));
Q_NR02 U101 ( .A0(xc_top.GFLock2), .A1(n11), .Z(n10));
Q_OR02 U102 ( .A0(xc_top.GFLock2), .A1(n12), .Z(n14));
Q_INV U103 ( .A(n11), .Z(n12));
Q_OR03 U104 ( .A0(n4), .A1(tkin), .A2(n13), .Z(n11));
Q_OR02 U105 ( .A0(Rtkin), .A1(CGFfull), .Z(n13));
Q_MX02 U106 ( .S(CLBfull), .A0(ireq), .A1(ireqR), .Z(n15));
Q_FDP0UA U107 ( .D(n15), .QTFCLK( ), .Q(ireqR));
Q_AN02 U108 ( .A0(CLBwr[0]), .A1(n6), .Z(n16));
Q_AN02 U109 ( .A0(CLBwr[1]), .A1(n6), .Z(n17));
Q_INV U110 ( .A(n16), .Z(n18));
Q_INV U111 ( .A(n17), .Z(n19));
Q_NR02 U112 ( .A0(n17), .A1(n16), .Z(n20));
Q_AN02 U113 ( .A0(n19), .A1(n16), .Z(n21));
Q_AN02 U114 ( .A0(n17), .A1(n18), .Z(n22));
Q_AN02 U115 ( .A0(n17), .A1(n16), .Z(n23));
Q_AN02 U116 ( .A0(n20), .A1(n6), .Z(n24));
Q_LDP0 \_zzLB_REG[0][0] ( .G(n24), .D(cbid[0]), .Q(\_zzLB[0][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][1] ( .G(n24), .D(cbid[1]), .Q(\_zzLB[0][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][2] ( .G(n24), .D(cbid[2]), .Q(\_zzLB[0][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][3] ( .G(n24), .D(cbid[3]), .Q(\_zzLB[0][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][4] ( .G(n24), .D(cbid[4]), .Q(\_zzLB[0][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][5] ( .G(n24), .D(cbid[5]), .Q(\_zzLB[0][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][6] ( .G(n24), .D(cbid[6]), .Q(\_zzLB[0][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][7] ( .G(n24), .D(cbid[7]), .Q(\_zzLB[0][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][8] ( .G(n24), .D(cbid[8]), .Q(\_zzLB[0][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][9] ( .G(n24), .D(cbid[9]), .Q(\_zzLB[0][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][10] ( .G(n24), .D(cbid[10]), .Q(\_zzLB[0][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][11] ( .G(n24), .D(cbid[11]), .Q(\_zzLB[0][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][12] ( .G(n24), .D(cbid[12]), .Q(\_zzLB[0][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][13] ( .G(n24), .D(cbid[13]), .Q(\_zzLB[0][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][14] ( .G(n24), .D(cbid[14]), .Q(\_zzLB[0][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][15] ( .G(n24), .D(cbid[15]), .Q(\_zzLB[0][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][16] ( .G(n24), .D(cbid[16]), .Q(\_zzLB[0][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][17] ( .G(n24), .D(cbid[17]), .Q(\_zzLB[0][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][18] ( .G(n24), .D(cbid[18]), .Q(\_zzLB[0][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][19] ( .G(n24), .D(cbid[19]), .Q(\_zzLB[0][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][20] ( .G(n24), .D(idata[0]), .Q(\_zzLB[0][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][21] ( .G(n24), .D(ireq), .Q(\_zzLB[0][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][0] ( .G(n21), .D(cbid[0]), .Q(\_zzLB[1][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][1] ( .G(n21), .D(cbid[1]), .Q(\_zzLB[1][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][2] ( .G(n21), .D(cbid[2]), .Q(\_zzLB[1][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][3] ( .G(n21), .D(cbid[3]), .Q(\_zzLB[1][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][4] ( .G(n21), .D(cbid[4]), .Q(\_zzLB[1][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][5] ( .G(n21), .D(cbid[5]), .Q(\_zzLB[1][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][6] ( .G(n21), .D(cbid[6]), .Q(\_zzLB[1][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][7] ( .G(n21), .D(cbid[7]), .Q(\_zzLB[1][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][8] ( .G(n21), .D(cbid[8]), .Q(\_zzLB[1][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][9] ( .G(n21), .D(cbid[9]), .Q(\_zzLB[1][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][10] ( .G(n21), .D(cbid[10]), .Q(\_zzLB[1][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][11] ( .G(n21), .D(cbid[11]), .Q(\_zzLB[1][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][12] ( .G(n21), .D(cbid[12]), .Q(\_zzLB[1][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][13] ( .G(n21), .D(cbid[13]), .Q(\_zzLB[1][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][14] ( .G(n21), .D(cbid[14]), .Q(\_zzLB[1][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][15] ( .G(n21), .D(cbid[15]), .Q(\_zzLB[1][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][16] ( .G(n21), .D(cbid[16]), .Q(\_zzLB[1][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][17] ( .G(n21), .D(cbid[17]), .Q(\_zzLB[1][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][18] ( .G(n21), .D(cbid[18]), .Q(\_zzLB[1][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][19] ( .G(n21), .D(cbid[19]), .Q(\_zzLB[1][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][20] ( .G(n21), .D(idata[0]), .Q(\_zzLB[1][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][21] ( .G(n21), .D(ireq), .Q(\_zzLB[1][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][0] ( .G(n22), .D(cbid[0]), .Q(\_zzLB[2][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][1] ( .G(n22), .D(cbid[1]), .Q(\_zzLB[2][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][2] ( .G(n22), .D(cbid[2]), .Q(\_zzLB[2][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][3] ( .G(n22), .D(cbid[3]), .Q(\_zzLB[2][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][4] ( .G(n22), .D(cbid[4]), .Q(\_zzLB[2][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][5] ( .G(n22), .D(cbid[5]), .Q(\_zzLB[2][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][6] ( .G(n22), .D(cbid[6]), .Q(\_zzLB[2][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][7] ( .G(n22), .D(cbid[7]), .Q(\_zzLB[2][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][8] ( .G(n22), .D(cbid[8]), .Q(\_zzLB[2][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][9] ( .G(n22), .D(cbid[9]), .Q(\_zzLB[2][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][10] ( .G(n22), .D(cbid[10]), .Q(\_zzLB[2][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][11] ( .G(n22), .D(cbid[11]), .Q(\_zzLB[2][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][12] ( .G(n22), .D(cbid[12]), .Q(\_zzLB[2][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][13] ( .G(n22), .D(cbid[13]), .Q(\_zzLB[2][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][14] ( .G(n22), .D(cbid[14]), .Q(\_zzLB[2][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][15] ( .G(n22), .D(cbid[15]), .Q(\_zzLB[2][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][16] ( .G(n22), .D(cbid[16]), .Q(\_zzLB[2][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][17] ( .G(n22), .D(cbid[17]), .Q(\_zzLB[2][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][18] ( .G(n22), .D(cbid[18]), .Q(\_zzLB[2][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][19] ( .G(n22), .D(cbid[19]), .Q(\_zzLB[2][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][20] ( .G(n22), .D(idata[0]), .Q(\_zzLB[2][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][21] ( .G(n22), .D(ireq), .Q(\_zzLB[2][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][0] ( .G(n23), .D(cbid[0]), .Q(\_zzLB[3][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][1] ( .G(n23), .D(cbid[1]), .Q(\_zzLB[3][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][2] ( .G(n23), .D(cbid[2]), .Q(\_zzLB[3][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][3] ( .G(n23), .D(cbid[3]), .Q(\_zzLB[3][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][4] ( .G(n23), .D(cbid[4]), .Q(\_zzLB[3][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][5] ( .G(n23), .D(cbid[5]), .Q(\_zzLB[3][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][6] ( .G(n23), .D(cbid[6]), .Q(\_zzLB[3][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][7] ( .G(n23), .D(cbid[7]), .Q(\_zzLB[3][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][8] ( .G(n23), .D(cbid[8]), .Q(\_zzLB[3][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][9] ( .G(n23), .D(cbid[9]), .Q(\_zzLB[3][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][10] ( .G(n23), .D(cbid[10]), .Q(\_zzLB[3][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][11] ( .G(n23), .D(cbid[11]), .Q(\_zzLB[3][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][12] ( .G(n23), .D(cbid[12]), .Q(\_zzLB[3][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][13] ( .G(n23), .D(cbid[13]), .Q(\_zzLB[3][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][14] ( .G(n23), .D(cbid[14]), .Q(\_zzLB[3][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][15] ( .G(n23), .D(cbid[15]), .Q(\_zzLB[3][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][16] ( .G(n23), .D(cbid[16]), .Q(\_zzLB[3][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][17] ( .G(n23), .D(cbid[17]), .Q(\_zzLB[3][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][18] ( .G(n23), .D(cbid[18]), .Q(\_zzLB[3][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][19] ( .G(n23), .D(cbid[19]), .Q(\_zzLB[3][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][20] ( .G(n23), .D(idata[0]), .Q(\_zzLB[3][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][21] ( .G(n23), .D(ireq), .Q(\_zzLB[3][21] ), .QN( ));
Q_MX04 U205 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][0] ), .A1(\_zzLB[1][0] ), .A2(\_zzLB[2][0] ), .A3(\_zzLB[3][0] ), .Z(ocbid[0]));
Q_MX04 U206 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][1] ), .A1(\_zzLB[1][1] ), .A2(\_zzLB[2][1] ), .A3(\_zzLB[3][1] ), .Z(ocbid[1]));
Q_MX04 U207 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][2] ), .A1(\_zzLB[1][2] ), .A2(\_zzLB[2][2] ), .A3(\_zzLB[3][2] ), .Z(ocbid[2]));
Q_MX04 U208 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][3] ), .A1(\_zzLB[1][3] ), .A2(\_zzLB[2][3] ), .A3(\_zzLB[3][3] ), .Z(ocbid[3]));
Q_MX04 U209 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][4] ), .A1(\_zzLB[1][4] ), .A2(\_zzLB[2][4] ), .A3(\_zzLB[3][4] ), .Z(ocbid[4]));
Q_MX04 U210 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][5] ), .A1(\_zzLB[1][5] ), .A2(\_zzLB[2][5] ), .A3(\_zzLB[3][5] ), .Z(ocbid[5]));
Q_MX04 U211 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][6] ), .A1(\_zzLB[1][6] ), .A2(\_zzLB[2][6] ), .A3(\_zzLB[3][6] ), .Z(ocbid[6]));
Q_MX04 U212 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][7] ), .A1(\_zzLB[1][7] ), .A2(\_zzLB[2][7] ), .A3(\_zzLB[3][7] ), .Z(ocbid[7]));
Q_MX04 U213 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][8] ), .A1(\_zzLB[1][8] ), .A2(\_zzLB[2][8] ), .A3(\_zzLB[3][8] ), .Z(ocbid[8]));
Q_MX04 U214 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][9] ), .A1(\_zzLB[1][9] ), .A2(\_zzLB[2][9] ), .A3(\_zzLB[3][9] ), .Z(ocbid[9]));
Q_MX04 U215 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][10] ), .A1(\_zzLB[1][10] ), .A2(\_zzLB[2][10] ), .A3(\_zzLB[3][10] ), .Z(ocbid[10]));
Q_MX04 U216 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][11] ), .A1(\_zzLB[1][11] ), .A2(\_zzLB[2][11] ), .A3(\_zzLB[3][11] ), .Z(ocbid[11]));
Q_MX04 U217 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][12] ), .A1(\_zzLB[1][12] ), .A2(\_zzLB[2][12] ), .A3(\_zzLB[3][12] ), .Z(ocbid[12]));
Q_MX04 U218 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][13] ), .A1(\_zzLB[1][13] ), .A2(\_zzLB[2][13] ), .A3(\_zzLB[3][13] ), .Z(ocbid[13]));
Q_MX04 U219 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][14] ), .A1(\_zzLB[1][14] ), .A2(\_zzLB[2][14] ), .A3(\_zzLB[3][14] ), .Z(ocbid[14]));
Q_MX04 U220 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][15] ), .A1(\_zzLB[1][15] ), .A2(\_zzLB[2][15] ), .A3(\_zzLB[3][15] ), .Z(ocbid[15]));
Q_MX04 U221 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][16] ), .A1(\_zzLB[1][16] ), .A2(\_zzLB[2][16] ), .A3(\_zzLB[3][16] ), .Z(ocbid[16]));
Q_MX04 U222 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][17] ), .A1(\_zzLB[1][17] ), .A2(\_zzLB[2][17] ), .A3(\_zzLB[3][17] ), .Z(ocbid[17]));
Q_MX04 U223 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][18] ), .A1(\_zzLB[1][18] ), .A2(\_zzLB[2][18] ), .A3(\_zzLB[3][18] ), .Z(ocbid[18]));
Q_MX04 U224 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][19] ), .A1(\_zzLB[1][19] ), .A2(\_zzLB[2][19] ), .A3(\_zzLB[3][19] ), .Z(ocbid[19]));
Q_MX04 U225 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][20] ), .A1(\_zzLB[1][20] ), .A2(\_zzLB[2][20] ), .A3(\_zzLB[3][20] ), .Z(odata[0]));
Q_MX04 U226 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][21] ), .A1(\_zzLB[1][21] ), .A2(\_zzLB[2][21] ), .A3(\_zzLB[3][21] ), .Z(oreq));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "_zzLB 1 21 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_gfifo_port"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
