
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_drbg_reggen ( set_drbg_expired_int, kdf_drbg_ctrl, seed0_valid, 
	seed0_internal_state_key, seed0_internal_state_value, 
	seed0_reseed_interval, seed1_valid, seed1_internal_state_key, 
	seed1_internal_state_value, seed1_reseed_interval, clk, rst_n, 
	wr_stb, wr_data, reg_addr, o_kdf_drbg_ctrl, 
	o_kdf_drbg_seed_0_reseed_interval_0, 
	o_kdf_drbg_seed_0_reseed_interval_1, 
	o_kdf_drbg_seed_0_state_key_127_96, 
	o_kdf_drbg_seed_0_state_key_159_128, 
	o_kdf_drbg_seed_0_state_key_191_160, 
	o_kdf_drbg_seed_0_state_key_223_192, 
	o_kdf_drbg_seed_0_state_key_255_224, 
	o_kdf_drbg_seed_0_state_key_31_0, o_kdf_drbg_seed_0_state_key_63_32, 
	o_kdf_drbg_seed_0_state_key_95_64, 
	o_kdf_drbg_seed_0_state_value_127_96, 
	o_kdf_drbg_seed_0_state_value_31_0, 
	o_kdf_drbg_seed_0_state_value_63_32, 
	o_kdf_drbg_seed_0_state_value_95_64, 
	o_kdf_drbg_seed_1_reseed_interval_0, 
	o_kdf_drbg_seed_1_reseed_interval_1, 
	o_kdf_drbg_seed_1_state_key_127_96, 
	o_kdf_drbg_seed_1_state_key_159_128, 
	o_kdf_drbg_seed_1_state_key_191_160, 
	o_kdf_drbg_seed_1_state_key_223_192, 
	o_kdf_drbg_seed_1_state_key_255_224, 
	o_kdf_drbg_seed_1_state_key_31_0, o_kdf_drbg_seed_1_state_key_63_32, 
	o_kdf_drbg_seed_1_state_key_95_64, 
	o_kdf_drbg_seed_1_state_value_127_96, 
	o_kdf_drbg_seed_1_state_value_31_0, 
	o_kdf_drbg_seed_1_state_value_63_32, 
	o_kdf_drbg_seed_1_state_value_95_64, seed0_invalidate, 
	seed1_invalidate);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output set_drbg_expired_int;
output [1:0] kdf_drbg_ctrl;
output seed0_valid;
output [255:0] seed0_internal_state_key;
output [127:0] seed0_internal_state_value;
output [47:0] seed0_reseed_interval;
output seed1_valid;
output [255:0] seed1_internal_state_key;
output [127:0] seed1_internal_state_value;
output [47:0] seed1_reseed_interval;
input clk;
input rst_n;
input wr_stb;
input [31:0] wr_data;
input [10:0] reg_addr;
input [1:0] o_kdf_drbg_ctrl;
input [31:0] o_kdf_drbg_seed_0_reseed_interval_0;
input [15:0] o_kdf_drbg_seed_0_reseed_interval_1;
input [31:0] o_kdf_drbg_seed_0_state_key_127_96;
input [31:0] o_kdf_drbg_seed_0_state_key_159_128;
input [31:0] o_kdf_drbg_seed_0_state_key_191_160;
input [31:0] o_kdf_drbg_seed_0_state_key_223_192;
input [31:0] o_kdf_drbg_seed_0_state_key_255_224;
input [31:0] o_kdf_drbg_seed_0_state_key_31_0;
input [31:0] o_kdf_drbg_seed_0_state_key_63_32;
input [31:0] o_kdf_drbg_seed_0_state_key_95_64;
input [31:0] o_kdf_drbg_seed_0_state_value_127_96;
input [31:0] o_kdf_drbg_seed_0_state_value_31_0;
input [31:0] o_kdf_drbg_seed_0_state_value_63_32;
input [31:0] o_kdf_drbg_seed_0_state_value_95_64;
input [31:0] o_kdf_drbg_seed_1_reseed_interval_0;
input [15:0] o_kdf_drbg_seed_1_reseed_interval_1;
input [31:0] o_kdf_drbg_seed_1_state_key_127_96;
input [31:0] o_kdf_drbg_seed_1_state_key_159_128;
input [31:0] o_kdf_drbg_seed_1_state_key_191_160;
input [31:0] o_kdf_drbg_seed_1_state_key_223_192;
input [31:0] o_kdf_drbg_seed_1_state_key_255_224;
input [31:0] o_kdf_drbg_seed_1_state_key_31_0;
input [31:0] o_kdf_drbg_seed_1_state_key_63_32;
input [31:0] o_kdf_drbg_seed_1_state_key_95_64;
input [31:0] o_kdf_drbg_seed_1_state_value_127_96;
input [31:0] o_kdf_drbg_seed_1_state_value_31_0;
input [31:0] o_kdf_drbg_seed_1_state_value_63_32;
input [31:0] o_kdf_drbg_seed_1_state_value_95_64;
input seed0_invalidate;
input seed1_invalidate;
wire _zy_simnet_seed0_valid_0_w$;
wire _zy_simnet_seed1_valid_1_w$;
ixc_assign _zz_strnp_8 ( _zy_simnet_seed1_valid_1_w$, seed1_valid);
ixc_assign _zz_strnp_7 ( _zy_simnet_seed0_valid_0_w$, seed0_valid);
ixc_assign_48 _zz_strnp_6 ( seed1_reseed_interval[47:0], { 
	o_kdf_drbg_seed_1_reseed_interval_1[15], 
	o_kdf_drbg_seed_1_reseed_interval_1[14], 
	o_kdf_drbg_seed_1_reseed_interval_1[13], 
	o_kdf_drbg_seed_1_reseed_interval_1[12], 
	o_kdf_drbg_seed_1_reseed_interval_1[11], 
	o_kdf_drbg_seed_1_reseed_interval_1[10], 
	o_kdf_drbg_seed_1_reseed_interval_1[9], 
	o_kdf_drbg_seed_1_reseed_interval_1[8], 
	o_kdf_drbg_seed_1_reseed_interval_1[7], 
	o_kdf_drbg_seed_1_reseed_interval_1[6], 
	o_kdf_drbg_seed_1_reseed_interval_1[5], 
	o_kdf_drbg_seed_1_reseed_interval_1[4], 
	o_kdf_drbg_seed_1_reseed_interval_1[3], 
	o_kdf_drbg_seed_1_reseed_interval_1[2], 
	o_kdf_drbg_seed_1_reseed_interval_1[1], 
	o_kdf_drbg_seed_1_reseed_interval_1[0], 
	o_kdf_drbg_seed_1_reseed_interval_0[31], 
	o_kdf_drbg_seed_1_reseed_interval_0[30], 
	o_kdf_drbg_seed_1_reseed_interval_0[29], 
	o_kdf_drbg_seed_1_reseed_interval_0[28], 
	o_kdf_drbg_seed_1_reseed_interval_0[27], 
	o_kdf_drbg_seed_1_reseed_interval_0[26], 
	o_kdf_drbg_seed_1_reseed_interval_0[25], 
	o_kdf_drbg_seed_1_reseed_interval_0[24], 
	o_kdf_drbg_seed_1_reseed_interval_0[23], 
	o_kdf_drbg_seed_1_reseed_interval_0[22], 
	o_kdf_drbg_seed_1_reseed_interval_0[21], 
	o_kdf_drbg_seed_1_reseed_interval_0[20], 
	o_kdf_drbg_seed_1_reseed_interval_0[19], 
	o_kdf_drbg_seed_1_reseed_interval_0[18], 
	o_kdf_drbg_seed_1_reseed_interval_0[17], 
	o_kdf_drbg_seed_1_reseed_interval_0[16], 
	o_kdf_drbg_seed_1_reseed_interval_0[15], 
	o_kdf_drbg_seed_1_reseed_interval_0[14], 
	o_kdf_drbg_seed_1_reseed_interval_0[13], 
	o_kdf_drbg_seed_1_reseed_interval_0[12], 
	o_kdf_drbg_seed_1_reseed_interval_0[11], 
	o_kdf_drbg_seed_1_reseed_interval_0[10], 
	o_kdf_drbg_seed_1_reseed_interval_0[9], 
	o_kdf_drbg_seed_1_reseed_interval_0[8], 
	o_kdf_drbg_seed_1_reseed_interval_0[7], 
	o_kdf_drbg_seed_1_reseed_interval_0[6], 
	o_kdf_drbg_seed_1_reseed_interval_0[5], 
	o_kdf_drbg_seed_1_reseed_interval_0[4], 
	o_kdf_drbg_seed_1_reseed_interval_0[3], 
	o_kdf_drbg_seed_1_reseed_interval_0[2], 
	o_kdf_drbg_seed_1_reseed_interval_0[1], 
	o_kdf_drbg_seed_1_reseed_interval_0[0]});
ixc_assign_128 _zz_strnp_5 ( seed1_internal_state_value[127:0], { 
	o_kdf_drbg_seed_1_state_value_127_96[31], 
	o_kdf_drbg_seed_1_state_value_127_96[30], 
	o_kdf_drbg_seed_1_state_value_127_96[29], 
	o_kdf_drbg_seed_1_state_value_127_96[28], 
	o_kdf_drbg_seed_1_state_value_127_96[27], 
	o_kdf_drbg_seed_1_state_value_127_96[26], 
	o_kdf_drbg_seed_1_state_value_127_96[25], 
	o_kdf_drbg_seed_1_state_value_127_96[24], 
	o_kdf_drbg_seed_1_state_value_127_96[23], 
	o_kdf_drbg_seed_1_state_value_127_96[22], 
	o_kdf_drbg_seed_1_state_value_127_96[21], 
	o_kdf_drbg_seed_1_state_value_127_96[20], 
	o_kdf_drbg_seed_1_state_value_127_96[19], 
	o_kdf_drbg_seed_1_state_value_127_96[18], 
	o_kdf_drbg_seed_1_state_value_127_96[17], 
	o_kdf_drbg_seed_1_state_value_127_96[16], 
	o_kdf_drbg_seed_1_state_value_127_96[15], 
	o_kdf_drbg_seed_1_state_value_127_96[14], 
	o_kdf_drbg_seed_1_state_value_127_96[13], 
	o_kdf_drbg_seed_1_state_value_127_96[12], 
	o_kdf_drbg_seed_1_state_value_127_96[11], 
	o_kdf_drbg_seed_1_state_value_127_96[10], 
	o_kdf_drbg_seed_1_state_value_127_96[9], 
	o_kdf_drbg_seed_1_state_value_127_96[8], 
	o_kdf_drbg_seed_1_state_value_127_96[7], 
	o_kdf_drbg_seed_1_state_value_127_96[6], 
	o_kdf_drbg_seed_1_state_value_127_96[5], 
	o_kdf_drbg_seed_1_state_value_127_96[4], 
	o_kdf_drbg_seed_1_state_value_127_96[3], 
	o_kdf_drbg_seed_1_state_value_127_96[2], 
	o_kdf_drbg_seed_1_state_value_127_96[1], 
	o_kdf_drbg_seed_1_state_value_127_96[0], 
	o_kdf_drbg_seed_1_state_value_95_64[31], 
	o_kdf_drbg_seed_1_state_value_95_64[30], 
	o_kdf_drbg_seed_1_state_value_95_64[29], 
	o_kdf_drbg_seed_1_state_value_95_64[28], 
	o_kdf_drbg_seed_1_state_value_95_64[27], 
	o_kdf_drbg_seed_1_state_value_95_64[26], 
	o_kdf_drbg_seed_1_state_value_95_64[25], 
	o_kdf_drbg_seed_1_state_value_95_64[24], 
	o_kdf_drbg_seed_1_state_value_95_64[23], 
	o_kdf_drbg_seed_1_state_value_95_64[22], 
	o_kdf_drbg_seed_1_state_value_95_64[21], 
	o_kdf_drbg_seed_1_state_value_95_64[20], 
	o_kdf_drbg_seed_1_state_value_95_64[19], 
	o_kdf_drbg_seed_1_state_value_95_64[18], 
	o_kdf_drbg_seed_1_state_value_95_64[17], 
	o_kdf_drbg_seed_1_state_value_95_64[16], 
	o_kdf_drbg_seed_1_state_value_95_64[15], 
	o_kdf_drbg_seed_1_state_value_95_64[14], 
	o_kdf_drbg_seed_1_state_value_95_64[13], 
	o_kdf_drbg_seed_1_state_value_95_64[12], 
	o_kdf_drbg_seed_1_state_value_95_64[11], 
	o_kdf_drbg_seed_1_state_value_95_64[10], 
	o_kdf_drbg_seed_1_state_value_95_64[9], 
	o_kdf_drbg_seed_1_state_value_95_64[8], 
	o_kdf_drbg_seed_1_state_value_95_64[7], 
	o_kdf_drbg_seed_1_state_value_95_64[6], 
	o_kdf_drbg_seed_1_state_value_95_64[5], 
	o_kdf_drbg_seed_1_state_value_95_64[4], 
	o_kdf_drbg_seed_1_state_value_95_64[3], 
	o_kdf_drbg_seed_1_state_value_95_64[2], 
	o_kdf_drbg_seed_1_state_value_95_64[1], 
	o_kdf_drbg_seed_1_state_value_95_64[0], 
	o_kdf_drbg_seed_1_state_value_63_32[31], 
	o_kdf_drbg_seed_1_state_value_63_32[30], 
	o_kdf_drbg_seed_1_state_value_63_32[29], 
	o_kdf_drbg_seed_1_state_value_63_32[28], 
	o_kdf_drbg_seed_1_state_value_63_32[27], 
	o_kdf_drbg_seed_1_state_value_63_32[26], 
	o_kdf_drbg_seed_1_state_value_63_32[25], 
	o_kdf_drbg_seed_1_state_value_63_32[24], 
	o_kdf_drbg_seed_1_state_value_63_32[23], 
	o_kdf_drbg_seed_1_state_value_63_32[22], 
	o_kdf_drbg_seed_1_state_value_63_32[21], 
	o_kdf_drbg_seed_1_state_value_63_32[20], 
	o_kdf_drbg_seed_1_state_value_63_32[19], 
	o_kdf_drbg_seed_1_state_value_63_32[18], 
	o_kdf_drbg_seed_1_state_value_63_32[17], 
	o_kdf_drbg_seed_1_state_value_63_32[16], 
	o_kdf_drbg_seed_1_state_value_63_32[15], 
	o_kdf_drbg_seed_1_state_value_63_32[14], 
	o_kdf_drbg_seed_1_state_value_63_32[13], 
	o_kdf_drbg_seed_1_state_value_63_32[12], 
	o_kdf_drbg_seed_1_state_value_63_32[11], 
	o_kdf_drbg_seed_1_state_value_63_32[10], 
	o_kdf_drbg_seed_1_state_value_63_32[9], 
	o_kdf_drbg_seed_1_state_value_63_32[8], 
	o_kdf_drbg_seed_1_state_value_63_32[7], 
	o_kdf_drbg_seed_1_state_value_63_32[6], 
	o_kdf_drbg_seed_1_state_value_63_32[5], 
	o_kdf_drbg_seed_1_state_value_63_32[4], 
	o_kdf_drbg_seed_1_state_value_63_32[3], 
	o_kdf_drbg_seed_1_state_value_63_32[2], 
	o_kdf_drbg_seed_1_state_value_63_32[1], 
	o_kdf_drbg_seed_1_state_value_63_32[0], 
	o_kdf_drbg_seed_1_state_value_31_0[31], 
	o_kdf_drbg_seed_1_state_value_31_0[30], 
	o_kdf_drbg_seed_1_state_value_31_0[29], 
	o_kdf_drbg_seed_1_state_value_31_0[28], 
	o_kdf_drbg_seed_1_state_value_31_0[27], 
	o_kdf_drbg_seed_1_state_value_31_0[26], 
	o_kdf_drbg_seed_1_state_value_31_0[25], 
	o_kdf_drbg_seed_1_state_value_31_0[24], 
	o_kdf_drbg_seed_1_state_value_31_0[23], 
	o_kdf_drbg_seed_1_state_value_31_0[22], 
	o_kdf_drbg_seed_1_state_value_31_0[21], 
	o_kdf_drbg_seed_1_state_value_31_0[20], 
	o_kdf_drbg_seed_1_state_value_31_0[19], 
	o_kdf_drbg_seed_1_state_value_31_0[18], 
	o_kdf_drbg_seed_1_state_value_31_0[17], 
	o_kdf_drbg_seed_1_state_value_31_0[16], 
	o_kdf_drbg_seed_1_state_value_31_0[15], 
	o_kdf_drbg_seed_1_state_value_31_0[14], 
	o_kdf_drbg_seed_1_state_value_31_0[13], 
	o_kdf_drbg_seed_1_state_value_31_0[12], 
	o_kdf_drbg_seed_1_state_value_31_0[11], 
	o_kdf_drbg_seed_1_state_value_31_0[10], 
	o_kdf_drbg_seed_1_state_value_31_0[9], 
	o_kdf_drbg_seed_1_state_value_31_0[8], 
	o_kdf_drbg_seed_1_state_value_31_0[7], 
	o_kdf_drbg_seed_1_state_value_31_0[6], 
	o_kdf_drbg_seed_1_state_value_31_0[5], 
	o_kdf_drbg_seed_1_state_value_31_0[4], 
	o_kdf_drbg_seed_1_state_value_31_0[3], 
	o_kdf_drbg_seed_1_state_value_31_0[2], 
	o_kdf_drbg_seed_1_state_value_31_0[1], 
	o_kdf_drbg_seed_1_state_value_31_0[0]});
ixc_assign_256 _zz_strnp_4 ( seed1_internal_state_key[255:0], { 
	o_kdf_drbg_seed_1_state_key_255_224[31], 
	o_kdf_drbg_seed_1_state_key_255_224[30], 
	o_kdf_drbg_seed_1_state_key_255_224[29], 
	o_kdf_drbg_seed_1_state_key_255_224[28], 
	o_kdf_drbg_seed_1_state_key_255_224[27], 
	o_kdf_drbg_seed_1_state_key_255_224[26], 
	o_kdf_drbg_seed_1_state_key_255_224[25], 
	o_kdf_drbg_seed_1_state_key_255_224[24], 
	o_kdf_drbg_seed_1_state_key_255_224[23], 
	o_kdf_drbg_seed_1_state_key_255_224[22], 
	o_kdf_drbg_seed_1_state_key_255_224[21], 
	o_kdf_drbg_seed_1_state_key_255_224[20], 
	o_kdf_drbg_seed_1_state_key_255_224[19], 
	o_kdf_drbg_seed_1_state_key_255_224[18], 
	o_kdf_drbg_seed_1_state_key_255_224[17], 
	o_kdf_drbg_seed_1_state_key_255_224[16], 
	o_kdf_drbg_seed_1_state_key_255_224[15], 
	o_kdf_drbg_seed_1_state_key_255_224[14], 
	o_kdf_drbg_seed_1_state_key_255_224[13], 
	o_kdf_drbg_seed_1_state_key_255_224[12], 
	o_kdf_drbg_seed_1_state_key_255_224[11], 
	o_kdf_drbg_seed_1_state_key_255_224[10], 
	o_kdf_drbg_seed_1_state_key_255_224[9], 
	o_kdf_drbg_seed_1_state_key_255_224[8], 
	o_kdf_drbg_seed_1_state_key_255_224[7], 
	o_kdf_drbg_seed_1_state_key_255_224[6], 
	o_kdf_drbg_seed_1_state_key_255_224[5], 
	o_kdf_drbg_seed_1_state_key_255_224[4], 
	o_kdf_drbg_seed_1_state_key_255_224[3], 
	o_kdf_drbg_seed_1_state_key_255_224[2], 
	o_kdf_drbg_seed_1_state_key_255_224[1], 
	o_kdf_drbg_seed_1_state_key_255_224[0], 
	o_kdf_drbg_seed_1_state_key_223_192[31], 
	o_kdf_drbg_seed_1_state_key_223_192[30], 
	o_kdf_drbg_seed_1_state_key_223_192[29], 
	o_kdf_drbg_seed_1_state_key_223_192[28], 
	o_kdf_drbg_seed_1_state_key_223_192[27], 
	o_kdf_drbg_seed_1_state_key_223_192[26], 
	o_kdf_drbg_seed_1_state_key_223_192[25], 
	o_kdf_drbg_seed_1_state_key_223_192[24], 
	o_kdf_drbg_seed_1_state_key_223_192[23], 
	o_kdf_drbg_seed_1_state_key_223_192[22], 
	o_kdf_drbg_seed_1_state_key_223_192[21], 
	o_kdf_drbg_seed_1_state_key_223_192[20], 
	o_kdf_drbg_seed_1_state_key_223_192[19], 
	o_kdf_drbg_seed_1_state_key_223_192[18], 
	o_kdf_drbg_seed_1_state_key_223_192[17], 
	o_kdf_drbg_seed_1_state_key_223_192[16], 
	o_kdf_drbg_seed_1_state_key_223_192[15], 
	o_kdf_drbg_seed_1_state_key_223_192[14], 
	o_kdf_drbg_seed_1_state_key_223_192[13], 
	o_kdf_drbg_seed_1_state_key_223_192[12], 
	o_kdf_drbg_seed_1_state_key_223_192[11], 
	o_kdf_drbg_seed_1_state_key_223_192[10], 
	o_kdf_drbg_seed_1_state_key_223_192[9], 
	o_kdf_drbg_seed_1_state_key_223_192[8], 
	o_kdf_drbg_seed_1_state_key_223_192[7], 
	o_kdf_drbg_seed_1_state_key_223_192[6], 
	o_kdf_drbg_seed_1_state_key_223_192[5], 
	o_kdf_drbg_seed_1_state_key_223_192[4], 
	o_kdf_drbg_seed_1_state_key_223_192[3], 
	o_kdf_drbg_seed_1_state_key_223_192[2], 
	o_kdf_drbg_seed_1_state_key_223_192[1], 
	o_kdf_drbg_seed_1_state_key_223_192[0], 
	o_kdf_drbg_seed_1_state_key_191_160[31], 
	o_kdf_drbg_seed_1_state_key_191_160[30], 
	o_kdf_drbg_seed_1_state_key_191_160[29], 
	o_kdf_drbg_seed_1_state_key_191_160[28], 
	o_kdf_drbg_seed_1_state_key_191_160[27], 
	o_kdf_drbg_seed_1_state_key_191_160[26], 
	o_kdf_drbg_seed_1_state_key_191_160[25], 
	o_kdf_drbg_seed_1_state_key_191_160[24], 
	o_kdf_drbg_seed_1_state_key_191_160[23], 
	o_kdf_drbg_seed_1_state_key_191_160[22], 
	o_kdf_drbg_seed_1_state_key_191_160[21], 
	o_kdf_drbg_seed_1_state_key_191_160[20], 
	o_kdf_drbg_seed_1_state_key_191_160[19], 
	o_kdf_drbg_seed_1_state_key_191_160[18], 
	o_kdf_drbg_seed_1_state_key_191_160[17], 
	o_kdf_drbg_seed_1_state_key_191_160[16], 
	o_kdf_drbg_seed_1_state_key_191_160[15], 
	o_kdf_drbg_seed_1_state_key_191_160[14], 
	o_kdf_drbg_seed_1_state_key_191_160[13], 
	o_kdf_drbg_seed_1_state_key_191_160[12], 
	o_kdf_drbg_seed_1_state_key_191_160[11], 
	o_kdf_drbg_seed_1_state_key_191_160[10], 
	o_kdf_drbg_seed_1_state_key_191_160[9], 
	o_kdf_drbg_seed_1_state_key_191_160[8], 
	o_kdf_drbg_seed_1_state_key_191_160[7], 
	o_kdf_drbg_seed_1_state_key_191_160[6], 
	o_kdf_drbg_seed_1_state_key_191_160[5], 
	o_kdf_drbg_seed_1_state_key_191_160[4], 
	o_kdf_drbg_seed_1_state_key_191_160[3], 
	o_kdf_drbg_seed_1_state_key_191_160[2], 
	o_kdf_drbg_seed_1_state_key_191_160[1], 
	o_kdf_drbg_seed_1_state_key_191_160[0], 
	o_kdf_drbg_seed_1_state_key_159_128[31], 
	o_kdf_drbg_seed_1_state_key_159_128[30], 
	o_kdf_drbg_seed_1_state_key_159_128[29], 
	o_kdf_drbg_seed_1_state_key_159_128[28], 
	o_kdf_drbg_seed_1_state_key_159_128[27], 
	o_kdf_drbg_seed_1_state_key_159_128[26], 
	o_kdf_drbg_seed_1_state_key_159_128[25], 
	o_kdf_drbg_seed_1_state_key_159_128[24], 
	o_kdf_drbg_seed_1_state_key_159_128[23], 
	o_kdf_drbg_seed_1_state_key_159_128[22], 
	o_kdf_drbg_seed_1_state_key_159_128[21], 
	o_kdf_drbg_seed_1_state_key_159_128[20], 
	o_kdf_drbg_seed_1_state_key_159_128[19], 
	o_kdf_drbg_seed_1_state_key_159_128[18], 
	o_kdf_drbg_seed_1_state_key_159_128[17], 
	o_kdf_drbg_seed_1_state_key_159_128[16], 
	o_kdf_drbg_seed_1_state_key_159_128[15], 
	o_kdf_drbg_seed_1_state_key_159_128[14], 
	o_kdf_drbg_seed_1_state_key_159_128[13], 
	o_kdf_drbg_seed_1_state_key_159_128[12], 
	o_kdf_drbg_seed_1_state_key_159_128[11], 
	o_kdf_drbg_seed_1_state_key_159_128[10], 
	o_kdf_drbg_seed_1_state_key_159_128[9], 
	o_kdf_drbg_seed_1_state_key_159_128[8], 
	o_kdf_drbg_seed_1_state_key_159_128[7], 
	o_kdf_drbg_seed_1_state_key_159_128[6], 
	o_kdf_drbg_seed_1_state_key_159_128[5], 
	o_kdf_drbg_seed_1_state_key_159_128[4], 
	o_kdf_drbg_seed_1_state_key_159_128[3], 
	o_kdf_drbg_seed_1_state_key_159_128[2], 
	o_kdf_drbg_seed_1_state_key_159_128[1], 
	o_kdf_drbg_seed_1_state_key_159_128[0], 
	o_kdf_drbg_seed_1_state_key_127_96[31], 
	o_kdf_drbg_seed_1_state_key_127_96[30], 
	o_kdf_drbg_seed_1_state_key_127_96[29], 
	o_kdf_drbg_seed_1_state_key_127_96[28], 
	o_kdf_drbg_seed_1_state_key_127_96[27], 
	o_kdf_drbg_seed_1_state_key_127_96[26], 
	o_kdf_drbg_seed_1_state_key_127_96[25], 
	o_kdf_drbg_seed_1_state_key_127_96[24], 
	o_kdf_drbg_seed_1_state_key_127_96[23], 
	o_kdf_drbg_seed_1_state_key_127_96[22], 
	o_kdf_drbg_seed_1_state_key_127_96[21], 
	o_kdf_drbg_seed_1_state_key_127_96[20], 
	o_kdf_drbg_seed_1_state_key_127_96[19], 
	o_kdf_drbg_seed_1_state_key_127_96[18], 
	o_kdf_drbg_seed_1_state_key_127_96[17], 
	o_kdf_drbg_seed_1_state_key_127_96[16], 
	o_kdf_drbg_seed_1_state_key_127_96[15], 
	o_kdf_drbg_seed_1_state_key_127_96[14], 
	o_kdf_drbg_seed_1_state_key_127_96[13], 
	o_kdf_drbg_seed_1_state_key_127_96[12], 
	o_kdf_drbg_seed_1_state_key_127_96[11], 
	o_kdf_drbg_seed_1_state_key_127_96[10], 
	o_kdf_drbg_seed_1_state_key_127_96[9], 
	o_kdf_drbg_seed_1_state_key_127_96[8], 
	o_kdf_drbg_seed_1_state_key_127_96[7], 
	o_kdf_drbg_seed_1_state_key_127_96[6], 
	o_kdf_drbg_seed_1_state_key_127_96[5], 
	o_kdf_drbg_seed_1_state_key_127_96[4], 
	o_kdf_drbg_seed_1_state_key_127_96[3], 
	o_kdf_drbg_seed_1_state_key_127_96[2], 
	o_kdf_drbg_seed_1_state_key_127_96[1], 
	o_kdf_drbg_seed_1_state_key_127_96[0], 
	o_kdf_drbg_seed_1_state_key_95_64[31], 
	o_kdf_drbg_seed_1_state_key_95_64[30], 
	o_kdf_drbg_seed_1_state_key_95_64[29], 
	o_kdf_drbg_seed_1_state_key_95_64[28], 
	o_kdf_drbg_seed_1_state_key_95_64[27], 
	o_kdf_drbg_seed_1_state_key_95_64[26], 
	o_kdf_drbg_seed_1_state_key_95_64[25], 
	o_kdf_drbg_seed_1_state_key_95_64[24], 
	o_kdf_drbg_seed_1_state_key_95_64[23], 
	o_kdf_drbg_seed_1_state_key_95_64[22], 
	o_kdf_drbg_seed_1_state_key_95_64[21], 
	o_kdf_drbg_seed_1_state_key_95_64[20], 
	o_kdf_drbg_seed_1_state_key_95_64[19], 
	o_kdf_drbg_seed_1_state_key_95_64[18], 
	o_kdf_drbg_seed_1_state_key_95_64[17], 
	o_kdf_drbg_seed_1_state_key_95_64[16], 
	o_kdf_drbg_seed_1_state_key_95_64[15], 
	o_kdf_drbg_seed_1_state_key_95_64[14], 
	o_kdf_drbg_seed_1_state_key_95_64[13], 
	o_kdf_drbg_seed_1_state_key_95_64[12], 
	o_kdf_drbg_seed_1_state_key_95_64[11], 
	o_kdf_drbg_seed_1_state_key_95_64[10], 
	o_kdf_drbg_seed_1_state_key_95_64[9], 
	o_kdf_drbg_seed_1_state_key_95_64[8], 
	o_kdf_drbg_seed_1_state_key_95_64[7], 
	o_kdf_drbg_seed_1_state_key_95_64[6], 
	o_kdf_drbg_seed_1_state_key_95_64[5], 
	o_kdf_drbg_seed_1_state_key_95_64[4], 
	o_kdf_drbg_seed_1_state_key_95_64[3], 
	o_kdf_drbg_seed_1_state_key_95_64[2], 
	o_kdf_drbg_seed_1_state_key_95_64[1], 
	o_kdf_drbg_seed_1_state_key_95_64[0], 
	o_kdf_drbg_seed_1_state_key_63_32[31], 
	o_kdf_drbg_seed_1_state_key_63_32[30], 
	o_kdf_drbg_seed_1_state_key_63_32[29], 
	o_kdf_drbg_seed_1_state_key_63_32[28], 
	o_kdf_drbg_seed_1_state_key_63_32[27], 
	o_kdf_drbg_seed_1_state_key_63_32[26], 
	o_kdf_drbg_seed_1_state_key_63_32[25], 
	o_kdf_drbg_seed_1_state_key_63_32[24], 
	o_kdf_drbg_seed_1_state_key_63_32[23], 
	o_kdf_drbg_seed_1_state_key_63_32[22], 
	o_kdf_drbg_seed_1_state_key_63_32[21], 
	o_kdf_drbg_seed_1_state_key_63_32[20], 
	o_kdf_drbg_seed_1_state_key_63_32[19], 
	o_kdf_drbg_seed_1_state_key_63_32[18], 
	o_kdf_drbg_seed_1_state_key_63_32[17], 
	o_kdf_drbg_seed_1_state_key_63_32[16], 
	o_kdf_drbg_seed_1_state_key_63_32[15], 
	o_kdf_drbg_seed_1_state_key_63_32[14], 
	o_kdf_drbg_seed_1_state_key_63_32[13], 
	o_kdf_drbg_seed_1_state_key_63_32[12], 
	o_kdf_drbg_seed_1_state_key_63_32[11], 
	o_kdf_drbg_seed_1_state_key_63_32[10], 
	o_kdf_drbg_seed_1_state_key_63_32[9], 
	o_kdf_drbg_seed_1_state_key_63_32[8], 
	o_kdf_drbg_seed_1_state_key_63_32[7], 
	o_kdf_drbg_seed_1_state_key_63_32[6], 
	o_kdf_drbg_seed_1_state_key_63_32[5], 
	o_kdf_drbg_seed_1_state_key_63_32[4], 
	o_kdf_drbg_seed_1_state_key_63_32[3], 
	o_kdf_drbg_seed_1_state_key_63_32[2], 
	o_kdf_drbg_seed_1_state_key_63_32[1], 
	o_kdf_drbg_seed_1_state_key_63_32[0], 
	o_kdf_drbg_seed_1_state_key_31_0[31], 
	o_kdf_drbg_seed_1_state_key_31_0[30], 
	o_kdf_drbg_seed_1_state_key_31_0[29], 
	o_kdf_drbg_seed_1_state_key_31_0[28], 
	o_kdf_drbg_seed_1_state_key_31_0[27], 
	o_kdf_drbg_seed_1_state_key_31_0[26], 
	o_kdf_drbg_seed_1_state_key_31_0[25], 
	o_kdf_drbg_seed_1_state_key_31_0[24], 
	o_kdf_drbg_seed_1_state_key_31_0[23], 
	o_kdf_drbg_seed_1_state_key_31_0[22], 
	o_kdf_drbg_seed_1_state_key_31_0[21], 
	o_kdf_drbg_seed_1_state_key_31_0[20], 
	o_kdf_drbg_seed_1_state_key_31_0[19], 
	o_kdf_drbg_seed_1_state_key_31_0[18], 
	o_kdf_drbg_seed_1_state_key_31_0[17], 
	o_kdf_drbg_seed_1_state_key_31_0[16], 
	o_kdf_drbg_seed_1_state_key_31_0[15], 
	o_kdf_drbg_seed_1_state_key_31_0[14], 
	o_kdf_drbg_seed_1_state_key_31_0[13], 
	o_kdf_drbg_seed_1_state_key_31_0[12], 
	o_kdf_drbg_seed_1_state_key_31_0[11], 
	o_kdf_drbg_seed_1_state_key_31_0[10], 
	o_kdf_drbg_seed_1_state_key_31_0[9], 
	o_kdf_drbg_seed_1_state_key_31_0[8], 
	o_kdf_drbg_seed_1_state_key_31_0[7], 
	o_kdf_drbg_seed_1_state_key_31_0[6], 
	o_kdf_drbg_seed_1_state_key_31_0[5], 
	o_kdf_drbg_seed_1_state_key_31_0[4], 
	o_kdf_drbg_seed_1_state_key_31_0[3], 
	o_kdf_drbg_seed_1_state_key_31_0[2], 
	o_kdf_drbg_seed_1_state_key_31_0[1], 
	o_kdf_drbg_seed_1_state_key_31_0[0]});
ixc_assign_48 _zz_strnp_3 ( seed0_reseed_interval[47:0], { 
	o_kdf_drbg_seed_0_reseed_interval_1[15], 
	o_kdf_drbg_seed_0_reseed_interval_1[14], 
	o_kdf_drbg_seed_0_reseed_interval_1[13], 
	o_kdf_drbg_seed_0_reseed_interval_1[12], 
	o_kdf_drbg_seed_0_reseed_interval_1[11], 
	o_kdf_drbg_seed_0_reseed_interval_1[10], 
	o_kdf_drbg_seed_0_reseed_interval_1[9], 
	o_kdf_drbg_seed_0_reseed_interval_1[8], 
	o_kdf_drbg_seed_0_reseed_interval_1[7], 
	o_kdf_drbg_seed_0_reseed_interval_1[6], 
	o_kdf_drbg_seed_0_reseed_interval_1[5], 
	o_kdf_drbg_seed_0_reseed_interval_1[4], 
	o_kdf_drbg_seed_0_reseed_interval_1[3], 
	o_kdf_drbg_seed_0_reseed_interval_1[2], 
	o_kdf_drbg_seed_0_reseed_interval_1[1], 
	o_kdf_drbg_seed_0_reseed_interval_1[0], 
	o_kdf_drbg_seed_0_reseed_interval_0[31], 
	o_kdf_drbg_seed_0_reseed_interval_0[30], 
	o_kdf_drbg_seed_0_reseed_interval_0[29], 
	o_kdf_drbg_seed_0_reseed_interval_0[28], 
	o_kdf_drbg_seed_0_reseed_interval_0[27], 
	o_kdf_drbg_seed_0_reseed_interval_0[26], 
	o_kdf_drbg_seed_0_reseed_interval_0[25], 
	o_kdf_drbg_seed_0_reseed_interval_0[24], 
	o_kdf_drbg_seed_0_reseed_interval_0[23], 
	o_kdf_drbg_seed_0_reseed_interval_0[22], 
	o_kdf_drbg_seed_0_reseed_interval_0[21], 
	o_kdf_drbg_seed_0_reseed_interval_0[20], 
	o_kdf_drbg_seed_0_reseed_interval_0[19], 
	o_kdf_drbg_seed_0_reseed_interval_0[18], 
	o_kdf_drbg_seed_0_reseed_interval_0[17], 
	o_kdf_drbg_seed_0_reseed_interval_0[16], 
	o_kdf_drbg_seed_0_reseed_interval_0[15], 
	o_kdf_drbg_seed_0_reseed_interval_0[14], 
	o_kdf_drbg_seed_0_reseed_interval_0[13], 
	o_kdf_drbg_seed_0_reseed_interval_0[12], 
	o_kdf_drbg_seed_0_reseed_interval_0[11], 
	o_kdf_drbg_seed_0_reseed_interval_0[10], 
	o_kdf_drbg_seed_0_reseed_interval_0[9], 
	o_kdf_drbg_seed_0_reseed_interval_0[8], 
	o_kdf_drbg_seed_0_reseed_interval_0[7], 
	o_kdf_drbg_seed_0_reseed_interval_0[6], 
	o_kdf_drbg_seed_0_reseed_interval_0[5], 
	o_kdf_drbg_seed_0_reseed_interval_0[4], 
	o_kdf_drbg_seed_0_reseed_interval_0[3], 
	o_kdf_drbg_seed_0_reseed_interval_0[2], 
	o_kdf_drbg_seed_0_reseed_interval_0[1], 
	o_kdf_drbg_seed_0_reseed_interval_0[0]});
ixc_assign_128 _zz_strnp_2 ( seed0_internal_state_value[127:0], { 
	o_kdf_drbg_seed_0_state_value_127_96[31], 
	o_kdf_drbg_seed_0_state_value_127_96[30], 
	o_kdf_drbg_seed_0_state_value_127_96[29], 
	o_kdf_drbg_seed_0_state_value_127_96[28], 
	o_kdf_drbg_seed_0_state_value_127_96[27], 
	o_kdf_drbg_seed_0_state_value_127_96[26], 
	o_kdf_drbg_seed_0_state_value_127_96[25], 
	o_kdf_drbg_seed_0_state_value_127_96[24], 
	o_kdf_drbg_seed_0_state_value_127_96[23], 
	o_kdf_drbg_seed_0_state_value_127_96[22], 
	o_kdf_drbg_seed_0_state_value_127_96[21], 
	o_kdf_drbg_seed_0_state_value_127_96[20], 
	o_kdf_drbg_seed_0_state_value_127_96[19], 
	o_kdf_drbg_seed_0_state_value_127_96[18], 
	o_kdf_drbg_seed_0_state_value_127_96[17], 
	o_kdf_drbg_seed_0_state_value_127_96[16], 
	o_kdf_drbg_seed_0_state_value_127_96[15], 
	o_kdf_drbg_seed_0_state_value_127_96[14], 
	o_kdf_drbg_seed_0_state_value_127_96[13], 
	o_kdf_drbg_seed_0_state_value_127_96[12], 
	o_kdf_drbg_seed_0_state_value_127_96[11], 
	o_kdf_drbg_seed_0_state_value_127_96[10], 
	o_kdf_drbg_seed_0_state_value_127_96[9], 
	o_kdf_drbg_seed_0_state_value_127_96[8], 
	o_kdf_drbg_seed_0_state_value_127_96[7], 
	o_kdf_drbg_seed_0_state_value_127_96[6], 
	o_kdf_drbg_seed_0_state_value_127_96[5], 
	o_kdf_drbg_seed_0_state_value_127_96[4], 
	o_kdf_drbg_seed_0_state_value_127_96[3], 
	o_kdf_drbg_seed_0_state_value_127_96[2], 
	o_kdf_drbg_seed_0_state_value_127_96[1], 
	o_kdf_drbg_seed_0_state_value_127_96[0], 
	o_kdf_drbg_seed_0_state_value_95_64[31], 
	o_kdf_drbg_seed_0_state_value_95_64[30], 
	o_kdf_drbg_seed_0_state_value_95_64[29], 
	o_kdf_drbg_seed_0_state_value_95_64[28], 
	o_kdf_drbg_seed_0_state_value_95_64[27], 
	o_kdf_drbg_seed_0_state_value_95_64[26], 
	o_kdf_drbg_seed_0_state_value_95_64[25], 
	o_kdf_drbg_seed_0_state_value_95_64[24], 
	o_kdf_drbg_seed_0_state_value_95_64[23], 
	o_kdf_drbg_seed_0_state_value_95_64[22], 
	o_kdf_drbg_seed_0_state_value_95_64[21], 
	o_kdf_drbg_seed_0_state_value_95_64[20], 
	o_kdf_drbg_seed_0_state_value_95_64[19], 
	o_kdf_drbg_seed_0_state_value_95_64[18], 
	o_kdf_drbg_seed_0_state_value_95_64[17], 
	o_kdf_drbg_seed_0_state_value_95_64[16], 
	o_kdf_drbg_seed_0_state_value_95_64[15], 
	o_kdf_drbg_seed_0_state_value_95_64[14], 
	o_kdf_drbg_seed_0_state_value_95_64[13], 
	o_kdf_drbg_seed_0_state_value_95_64[12], 
	o_kdf_drbg_seed_0_state_value_95_64[11], 
	o_kdf_drbg_seed_0_state_value_95_64[10], 
	o_kdf_drbg_seed_0_state_value_95_64[9], 
	o_kdf_drbg_seed_0_state_value_95_64[8], 
	o_kdf_drbg_seed_0_state_value_95_64[7], 
	o_kdf_drbg_seed_0_state_value_95_64[6], 
	o_kdf_drbg_seed_0_state_value_95_64[5], 
	o_kdf_drbg_seed_0_state_value_95_64[4], 
	o_kdf_drbg_seed_0_state_value_95_64[3], 
	o_kdf_drbg_seed_0_state_value_95_64[2], 
	o_kdf_drbg_seed_0_state_value_95_64[1], 
	o_kdf_drbg_seed_0_state_value_95_64[0], 
	o_kdf_drbg_seed_0_state_value_63_32[31], 
	o_kdf_drbg_seed_0_state_value_63_32[30], 
	o_kdf_drbg_seed_0_state_value_63_32[29], 
	o_kdf_drbg_seed_0_state_value_63_32[28], 
	o_kdf_drbg_seed_0_state_value_63_32[27], 
	o_kdf_drbg_seed_0_state_value_63_32[26], 
	o_kdf_drbg_seed_0_state_value_63_32[25], 
	o_kdf_drbg_seed_0_state_value_63_32[24], 
	o_kdf_drbg_seed_0_state_value_63_32[23], 
	o_kdf_drbg_seed_0_state_value_63_32[22], 
	o_kdf_drbg_seed_0_state_value_63_32[21], 
	o_kdf_drbg_seed_0_state_value_63_32[20], 
	o_kdf_drbg_seed_0_state_value_63_32[19], 
	o_kdf_drbg_seed_0_state_value_63_32[18], 
	o_kdf_drbg_seed_0_state_value_63_32[17], 
	o_kdf_drbg_seed_0_state_value_63_32[16], 
	o_kdf_drbg_seed_0_state_value_63_32[15], 
	o_kdf_drbg_seed_0_state_value_63_32[14], 
	o_kdf_drbg_seed_0_state_value_63_32[13], 
	o_kdf_drbg_seed_0_state_value_63_32[12], 
	o_kdf_drbg_seed_0_state_value_63_32[11], 
	o_kdf_drbg_seed_0_state_value_63_32[10], 
	o_kdf_drbg_seed_0_state_value_63_32[9], 
	o_kdf_drbg_seed_0_state_value_63_32[8], 
	o_kdf_drbg_seed_0_state_value_63_32[7], 
	o_kdf_drbg_seed_0_state_value_63_32[6], 
	o_kdf_drbg_seed_0_state_value_63_32[5], 
	o_kdf_drbg_seed_0_state_value_63_32[4], 
	o_kdf_drbg_seed_0_state_value_63_32[3], 
	o_kdf_drbg_seed_0_state_value_63_32[2], 
	o_kdf_drbg_seed_0_state_value_63_32[1], 
	o_kdf_drbg_seed_0_state_value_63_32[0], 
	o_kdf_drbg_seed_0_state_value_31_0[31], 
	o_kdf_drbg_seed_0_state_value_31_0[30], 
	o_kdf_drbg_seed_0_state_value_31_0[29], 
	o_kdf_drbg_seed_0_state_value_31_0[28], 
	o_kdf_drbg_seed_0_state_value_31_0[27], 
	o_kdf_drbg_seed_0_state_value_31_0[26], 
	o_kdf_drbg_seed_0_state_value_31_0[25], 
	o_kdf_drbg_seed_0_state_value_31_0[24], 
	o_kdf_drbg_seed_0_state_value_31_0[23], 
	o_kdf_drbg_seed_0_state_value_31_0[22], 
	o_kdf_drbg_seed_0_state_value_31_0[21], 
	o_kdf_drbg_seed_0_state_value_31_0[20], 
	o_kdf_drbg_seed_0_state_value_31_0[19], 
	o_kdf_drbg_seed_0_state_value_31_0[18], 
	o_kdf_drbg_seed_0_state_value_31_0[17], 
	o_kdf_drbg_seed_0_state_value_31_0[16], 
	o_kdf_drbg_seed_0_state_value_31_0[15], 
	o_kdf_drbg_seed_0_state_value_31_0[14], 
	o_kdf_drbg_seed_0_state_value_31_0[13], 
	o_kdf_drbg_seed_0_state_value_31_0[12], 
	o_kdf_drbg_seed_0_state_value_31_0[11], 
	o_kdf_drbg_seed_0_state_value_31_0[10], 
	o_kdf_drbg_seed_0_state_value_31_0[9], 
	o_kdf_drbg_seed_0_state_value_31_0[8], 
	o_kdf_drbg_seed_0_state_value_31_0[7], 
	o_kdf_drbg_seed_0_state_value_31_0[6], 
	o_kdf_drbg_seed_0_state_value_31_0[5], 
	o_kdf_drbg_seed_0_state_value_31_0[4], 
	o_kdf_drbg_seed_0_state_value_31_0[3], 
	o_kdf_drbg_seed_0_state_value_31_0[2], 
	o_kdf_drbg_seed_0_state_value_31_0[1], 
	o_kdf_drbg_seed_0_state_value_31_0[0]});
ixc_assign_256 _zz_strnp_1 ( seed0_internal_state_key[255:0], { 
	o_kdf_drbg_seed_0_state_key_255_224[31], 
	o_kdf_drbg_seed_0_state_key_255_224[30], 
	o_kdf_drbg_seed_0_state_key_255_224[29], 
	o_kdf_drbg_seed_0_state_key_255_224[28], 
	o_kdf_drbg_seed_0_state_key_255_224[27], 
	o_kdf_drbg_seed_0_state_key_255_224[26], 
	o_kdf_drbg_seed_0_state_key_255_224[25], 
	o_kdf_drbg_seed_0_state_key_255_224[24], 
	o_kdf_drbg_seed_0_state_key_255_224[23], 
	o_kdf_drbg_seed_0_state_key_255_224[22], 
	o_kdf_drbg_seed_0_state_key_255_224[21], 
	o_kdf_drbg_seed_0_state_key_255_224[20], 
	o_kdf_drbg_seed_0_state_key_255_224[19], 
	o_kdf_drbg_seed_0_state_key_255_224[18], 
	o_kdf_drbg_seed_0_state_key_255_224[17], 
	o_kdf_drbg_seed_0_state_key_255_224[16], 
	o_kdf_drbg_seed_0_state_key_255_224[15], 
	o_kdf_drbg_seed_0_state_key_255_224[14], 
	o_kdf_drbg_seed_0_state_key_255_224[13], 
	o_kdf_drbg_seed_0_state_key_255_224[12], 
	o_kdf_drbg_seed_0_state_key_255_224[11], 
	o_kdf_drbg_seed_0_state_key_255_224[10], 
	o_kdf_drbg_seed_0_state_key_255_224[9], 
	o_kdf_drbg_seed_0_state_key_255_224[8], 
	o_kdf_drbg_seed_0_state_key_255_224[7], 
	o_kdf_drbg_seed_0_state_key_255_224[6], 
	o_kdf_drbg_seed_0_state_key_255_224[5], 
	o_kdf_drbg_seed_0_state_key_255_224[4], 
	o_kdf_drbg_seed_0_state_key_255_224[3], 
	o_kdf_drbg_seed_0_state_key_255_224[2], 
	o_kdf_drbg_seed_0_state_key_255_224[1], 
	o_kdf_drbg_seed_0_state_key_255_224[0], 
	o_kdf_drbg_seed_0_state_key_223_192[31], 
	o_kdf_drbg_seed_0_state_key_223_192[30], 
	o_kdf_drbg_seed_0_state_key_223_192[29], 
	o_kdf_drbg_seed_0_state_key_223_192[28], 
	o_kdf_drbg_seed_0_state_key_223_192[27], 
	o_kdf_drbg_seed_0_state_key_223_192[26], 
	o_kdf_drbg_seed_0_state_key_223_192[25], 
	o_kdf_drbg_seed_0_state_key_223_192[24], 
	o_kdf_drbg_seed_0_state_key_223_192[23], 
	o_kdf_drbg_seed_0_state_key_223_192[22], 
	o_kdf_drbg_seed_0_state_key_223_192[21], 
	o_kdf_drbg_seed_0_state_key_223_192[20], 
	o_kdf_drbg_seed_0_state_key_223_192[19], 
	o_kdf_drbg_seed_0_state_key_223_192[18], 
	o_kdf_drbg_seed_0_state_key_223_192[17], 
	o_kdf_drbg_seed_0_state_key_223_192[16], 
	o_kdf_drbg_seed_0_state_key_223_192[15], 
	o_kdf_drbg_seed_0_state_key_223_192[14], 
	o_kdf_drbg_seed_0_state_key_223_192[13], 
	o_kdf_drbg_seed_0_state_key_223_192[12], 
	o_kdf_drbg_seed_0_state_key_223_192[11], 
	o_kdf_drbg_seed_0_state_key_223_192[10], 
	o_kdf_drbg_seed_0_state_key_223_192[9], 
	o_kdf_drbg_seed_0_state_key_223_192[8], 
	o_kdf_drbg_seed_0_state_key_223_192[7], 
	o_kdf_drbg_seed_0_state_key_223_192[6], 
	o_kdf_drbg_seed_0_state_key_223_192[5], 
	o_kdf_drbg_seed_0_state_key_223_192[4], 
	o_kdf_drbg_seed_0_state_key_223_192[3], 
	o_kdf_drbg_seed_0_state_key_223_192[2], 
	o_kdf_drbg_seed_0_state_key_223_192[1], 
	o_kdf_drbg_seed_0_state_key_223_192[0], 
	o_kdf_drbg_seed_0_state_key_191_160[31], 
	o_kdf_drbg_seed_0_state_key_191_160[30], 
	o_kdf_drbg_seed_0_state_key_191_160[29], 
	o_kdf_drbg_seed_0_state_key_191_160[28], 
	o_kdf_drbg_seed_0_state_key_191_160[27], 
	o_kdf_drbg_seed_0_state_key_191_160[26], 
	o_kdf_drbg_seed_0_state_key_191_160[25], 
	o_kdf_drbg_seed_0_state_key_191_160[24], 
	o_kdf_drbg_seed_0_state_key_191_160[23], 
	o_kdf_drbg_seed_0_state_key_191_160[22], 
	o_kdf_drbg_seed_0_state_key_191_160[21], 
	o_kdf_drbg_seed_0_state_key_191_160[20], 
	o_kdf_drbg_seed_0_state_key_191_160[19], 
	o_kdf_drbg_seed_0_state_key_191_160[18], 
	o_kdf_drbg_seed_0_state_key_191_160[17], 
	o_kdf_drbg_seed_0_state_key_191_160[16], 
	o_kdf_drbg_seed_0_state_key_191_160[15], 
	o_kdf_drbg_seed_0_state_key_191_160[14], 
	o_kdf_drbg_seed_0_state_key_191_160[13], 
	o_kdf_drbg_seed_0_state_key_191_160[12], 
	o_kdf_drbg_seed_0_state_key_191_160[11], 
	o_kdf_drbg_seed_0_state_key_191_160[10], 
	o_kdf_drbg_seed_0_state_key_191_160[9], 
	o_kdf_drbg_seed_0_state_key_191_160[8], 
	o_kdf_drbg_seed_0_state_key_191_160[7], 
	o_kdf_drbg_seed_0_state_key_191_160[6], 
	o_kdf_drbg_seed_0_state_key_191_160[5], 
	o_kdf_drbg_seed_0_state_key_191_160[4], 
	o_kdf_drbg_seed_0_state_key_191_160[3], 
	o_kdf_drbg_seed_0_state_key_191_160[2], 
	o_kdf_drbg_seed_0_state_key_191_160[1], 
	o_kdf_drbg_seed_0_state_key_191_160[0], 
	o_kdf_drbg_seed_0_state_key_159_128[31], 
	o_kdf_drbg_seed_0_state_key_159_128[30], 
	o_kdf_drbg_seed_0_state_key_159_128[29], 
	o_kdf_drbg_seed_0_state_key_159_128[28], 
	o_kdf_drbg_seed_0_state_key_159_128[27], 
	o_kdf_drbg_seed_0_state_key_159_128[26], 
	o_kdf_drbg_seed_0_state_key_159_128[25], 
	o_kdf_drbg_seed_0_state_key_159_128[24], 
	o_kdf_drbg_seed_0_state_key_159_128[23], 
	o_kdf_drbg_seed_0_state_key_159_128[22], 
	o_kdf_drbg_seed_0_state_key_159_128[21], 
	o_kdf_drbg_seed_0_state_key_159_128[20], 
	o_kdf_drbg_seed_0_state_key_159_128[19], 
	o_kdf_drbg_seed_0_state_key_159_128[18], 
	o_kdf_drbg_seed_0_state_key_159_128[17], 
	o_kdf_drbg_seed_0_state_key_159_128[16], 
	o_kdf_drbg_seed_0_state_key_159_128[15], 
	o_kdf_drbg_seed_0_state_key_159_128[14], 
	o_kdf_drbg_seed_0_state_key_159_128[13], 
	o_kdf_drbg_seed_0_state_key_159_128[12], 
	o_kdf_drbg_seed_0_state_key_159_128[11], 
	o_kdf_drbg_seed_0_state_key_159_128[10], 
	o_kdf_drbg_seed_0_state_key_159_128[9], 
	o_kdf_drbg_seed_0_state_key_159_128[8], 
	o_kdf_drbg_seed_0_state_key_159_128[7], 
	o_kdf_drbg_seed_0_state_key_159_128[6], 
	o_kdf_drbg_seed_0_state_key_159_128[5], 
	o_kdf_drbg_seed_0_state_key_159_128[4], 
	o_kdf_drbg_seed_0_state_key_159_128[3], 
	o_kdf_drbg_seed_0_state_key_159_128[2], 
	o_kdf_drbg_seed_0_state_key_159_128[1], 
	o_kdf_drbg_seed_0_state_key_159_128[0], 
	o_kdf_drbg_seed_0_state_key_127_96[31], 
	o_kdf_drbg_seed_0_state_key_127_96[30], 
	o_kdf_drbg_seed_0_state_key_127_96[29], 
	o_kdf_drbg_seed_0_state_key_127_96[28], 
	o_kdf_drbg_seed_0_state_key_127_96[27], 
	o_kdf_drbg_seed_0_state_key_127_96[26], 
	o_kdf_drbg_seed_0_state_key_127_96[25], 
	o_kdf_drbg_seed_0_state_key_127_96[24], 
	o_kdf_drbg_seed_0_state_key_127_96[23], 
	o_kdf_drbg_seed_0_state_key_127_96[22], 
	o_kdf_drbg_seed_0_state_key_127_96[21], 
	o_kdf_drbg_seed_0_state_key_127_96[20], 
	o_kdf_drbg_seed_0_state_key_127_96[19], 
	o_kdf_drbg_seed_0_state_key_127_96[18], 
	o_kdf_drbg_seed_0_state_key_127_96[17], 
	o_kdf_drbg_seed_0_state_key_127_96[16], 
	o_kdf_drbg_seed_0_state_key_127_96[15], 
	o_kdf_drbg_seed_0_state_key_127_96[14], 
	o_kdf_drbg_seed_0_state_key_127_96[13], 
	o_kdf_drbg_seed_0_state_key_127_96[12], 
	o_kdf_drbg_seed_0_state_key_127_96[11], 
	o_kdf_drbg_seed_0_state_key_127_96[10], 
	o_kdf_drbg_seed_0_state_key_127_96[9], 
	o_kdf_drbg_seed_0_state_key_127_96[8], 
	o_kdf_drbg_seed_0_state_key_127_96[7], 
	o_kdf_drbg_seed_0_state_key_127_96[6], 
	o_kdf_drbg_seed_0_state_key_127_96[5], 
	o_kdf_drbg_seed_0_state_key_127_96[4], 
	o_kdf_drbg_seed_0_state_key_127_96[3], 
	o_kdf_drbg_seed_0_state_key_127_96[2], 
	o_kdf_drbg_seed_0_state_key_127_96[1], 
	o_kdf_drbg_seed_0_state_key_127_96[0], 
	o_kdf_drbg_seed_0_state_key_95_64[31], 
	o_kdf_drbg_seed_0_state_key_95_64[30], 
	o_kdf_drbg_seed_0_state_key_95_64[29], 
	o_kdf_drbg_seed_0_state_key_95_64[28], 
	o_kdf_drbg_seed_0_state_key_95_64[27], 
	o_kdf_drbg_seed_0_state_key_95_64[26], 
	o_kdf_drbg_seed_0_state_key_95_64[25], 
	o_kdf_drbg_seed_0_state_key_95_64[24], 
	o_kdf_drbg_seed_0_state_key_95_64[23], 
	o_kdf_drbg_seed_0_state_key_95_64[22], 
	o_kdf_drbg_seed_0_state_key_95_64[21], 
	o_kdf_drbg_seed_0_state_key_95_64[20], 
	o_kdf_drbg_seed_0_state_key_95_64[19], 
	o_kdf_drbg_seed_0_state_key_95_64[18], 
	o_kdf_drbg_seed_0_state_key_95_64[17], 
	o_kdf_drbg_seed_0_state_key_95_64[16], 
	o_kdf_drbg_seed_0_state_key_95_64[15], 
	o_kdf_drbg_seed_0_state_key_95_64[14], 
	o_kdf_drbg_seed_0_state_key_95_64[13], 
	o_kdf_drbg_seed_0_state_key_95_64[12], 
	o_kdf_drbg_seed_0_state_key_95_64[11], 
	o_kdf_drbg_seed_0_state_key_95_64[10], 
	o_kdf_drbg_seed_0_state_key_95_64[9], 
	o_kdf_drbg_seed_0_state_key_95_64[8], 
	o_kdf_drbg_seed_0_state_key_95_64[7], 
	o_kdf_drbg_seed_0_state_key_95_64[6], 
	o_kdf_drbg_seed_0_state_key_95_64[5], 
	o_kdf_drbg_seed_0_state_key_95_64[4], 
	o_kdf_drbg_seed_0_state_key_95_64[3], 
	o_kdf_drbg_seed_0_state_key_95_64[2], 
	o_kdf_drbg_seed_0_state_key_95_64[1], 
	o_kdf_drbg_seed_0_state_key_95_64[0], 
	o_kdf_drbg_seed_0_state_key_63_32[31], 
	o_kdf_drbg_seed_0_state_key_63_32[30], 
	o_kdf_drbg_seed_0_state_key_63_32[29], 
	o_kdf_drbg_seed_0_state_key_63_32[28], 
	o_kdf_drbg_seed_0_state_key_63_32[27], 
	o_kdf_drbg_seed_0_state_key_63_32[26], 
	o_kdf_drbg_seed_0_state_key_63_32[25], 
	o_kdf_drbg_seed_0_state_key_63_32[24], 
	o_kdf_drbg_seed_0_state_key_63_32[23], 
	o_kdf_drbg_seed_0_state_key_63_32[22], 
	o_kdf_drbg_seed_0_state_key_63_32[21], 
	o_kdf_drbg_seed_0_state_key_63_32[20], 
	o_kdf_drbg_seed_0_state_key_63_32[19], 
	o_kdf_drbg_seed_0_state_key_63_32[18], 
	o_kdf_drbg_seed_0_state_key_63_32[17], 
	o_kdf_drbg_seed_0_state_key_63_32[16], 
	o_kdf_drbg_seed_0_state_key_63_32[15], 
	o_kdf_drbg_seed_0_state_key_63_32[14], 
	o_kdf_drbg_seed_0_state_key_63_32[13], 
	o_kdf_drbg_seed_0_state_key_63_32[12], 
	o_kdf_drbg_seed_0_state_key_63_32[11], 
	o_kdf_drbg_seed_0_state_key_63_32[10], 
	o_kdf_drbg_seed_0_state_key_63_32[9], 
	o_kdf_drbg_seed_0_state_key_63_32[8], 
	o_kdf_drbg_seed_0_state_key_63_32[7], 
	o_kdf_drbg_seed_0_state_key_63_32[6], 
	o_kdf_drbg_seed_0_state_key_63_32[5], 
	o_kdf_drbg_seed_0_state_key_63_32[4], 
	o_kdf_drbg_seed_0_state_key_63_32[3], 
	o_kdf_drbg_seed_0_state_key_63_32[2], 
	o_kdf_drbg_seed_0_state_key_63_32[1], 
	o_kdf_drbg_seed_0_state_key_63_32[0], 
	o_kdf_drbg_seed_0_state_key_31_0[31], 
	o_kdf_drbg_seed_0_state_key_31_0[30], 
	o_kdf_drbg_seed_0_state_key_31_0[29], 
	o_kdf_drbg_seed_0_state_key_31_0[28], 
	o_kdf_drbg_seed_0_state_key_31_0[27], 
	o_kdf_drbg_seed_0_state_key_31_0[26], 
	o_kdf_drbg_seed_0_state_key_31_0[25], 
	o_kdf_drbg_seed_0_state_key_31_0[24], 
	o_kdf_drbg_seed_0_state_key_31_0[23], 
	o_kdf_drbg_seed_0_state_key_31_0[22], 
	o_kdf_drbg_seed_0_state_key_31_0[21], 
	o_kdf_drbg_seed_0_state_key_31_0[20], 
	o_kdf_drbg_seed_0_state_key_31_0[19], 
	o_kdf_drbg_seed_0_state_key_31_0[18], 
	o_kdf_drbg_seed_0_state_key_31_0[17], 
	o_kdf_drbg_seed_0_state_key_31_0[16], 
	o_kdf_drbg_seed_0_state_key_31_0[15], 
	o_kdf_drbg_seed_0_state_key_31_0[14], 
	o_kdf_drbg_seed_0_state_key_31_0[13], 
	o_kdf_drbg_seed_0_state_key_31_0[12], 
	o_kdf_drbg_seed_0_state_key_31_0[11], 
	o_kdf_drbg_seed_0_state_key_31_0[10], 
	o_kdf_drbg_seed_0_state_key_31_0[9], 
	o_kdf_drbg_seed_0_state_key_31_0[8], 
	o_kdf_drbg_seed_0_state_key_31_0[7], 
	o_kdf_drbg_seed_0_state_key_31_0[6], 
	o_kdf_drbg_seed_0_state_key_31_0[5], 
	o_kdf_drbg_seed_0_state_key_31_0[4], 
	o_kdf_drbg_seed_0_state_key_31_0[3], 
	o_kdf_drbg_seed_0_state_key_31_0[2], 
	o_kdf_drbg_seed_0_state_key_31_0[1], 
	o_kdf_drbg_seed_0_state_key_31_0[0]});
ixc_assign_2 _zz_strnp_0 ( kdf_drbg_ctrl[1:0], { seed1_valid, seed0_valid});
Q_AN02 U9 ( .A0(seed1_valid), .A1(seed1_invalidate), .Z(n1));
Q_AO21 U10 ( .A0(seed0_valid), .A1(seed0_invalidate), .B0(n1), .Z(set_drbg_expired_int));
Q_INV U11 ( .A(reg_addr[3]), .Z(n2));
Q_INV U12 ( .A(reg_addr[8]), .Z(n3));
Q_INV U13 ( .A(reg_addr[9]), .Z(n4));
Q_OR03 U14 ( .A0(reg_addr[10]), .A1(n4), .A2(n3), .Z(n5));
Q_OR03 U15 ( .A0(reg_addr[7]), .A1(reg_addr[6]), .A2(reg_addr[5]), .Z(n6));
Q_OR03 U16 ( .A0(reg_addr[4]), .A1(n2), .A2(reg_addr[2]), .Z(n7));
Q_OR03 U17 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n5), .Z(n8));
Q_NR03 U18 ( .A0(n6), .A1(n7), .A2(n8), .Z(n9));
Q_AN02 U19 ( .A0(wr_stb), .A1(n9), .Z(n13));
Q_AN02 U20 ( .A0(n12), .A1(wr_data[0]), .Z(n10));
Q_OR02 U21 ( .A0(seed0_invalidate), .A1(n13), .Z(n11));
Q_INV U22 ( .A(seed0_invalidate), .Z(n12));
Q_AN02 U23 ( .A0(n16), .A1(wr_data[1]), .Z(n14));
Q_OR02 U24 ( .A0(seed1_invalidate), .A1(n13), .Z(n15));
Q_INV U25 ( .A(seed1_invalidate), .Z(n16));
Q_FDP4EP seed1_valid_REG  ( .CK(clk), .CE(n15), .R(n17), .D(n14), .Q(seed1_valid));
Q_INV U27 ( .A(rst_n), .Z(n17));
Q_FDP4EP seed0_valid_REG  ( .CK(clk), .CE(n11), .R(n17), .D(n10), .Q(seed0_valid));
endmodule
