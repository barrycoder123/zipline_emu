architecture module of sfifo_conns is
  component sfifo_conns_0
  end component ;


begin
  sc0 : sfifo_conns_0
     ;
end module;
